// This is the unpowered netlist.
module posit_unit (clk,
    rst,
    io_in,
    io_out);
 input clk;
 input rst;
 input [2:0] io_in;
 output [3:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire \cmd[0] ;
 wire \cmd[6] ;
 wire \cmd[7] ;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \in_reg[0] ;
 wire \in_reg[10] ;
 wire \in_reg[11] ;
 wire \in_reg[12] ;
 wire \in_reg[13] ;
 wire \in_reg[14] ;
 wire \in_reg[15] ;
 wire \in_reg[1] ;
 wire \in_reg[2] ;
 wire \in_reg[3] ;
 wire \in_reg[4] ;
 wire \in_reg[5] ;
 wire \in_reg[6] ;
 wire \in_reg[7] ;
 wire \in_reg[8] ;
 wire \in_reg[9] ;
 wire net6;
 wire net7;
 wire clknet_0_clk;
 wire last_SCLK;
 wire mode;
 wire \out_reg[0] ;
 wire \out_reg[10] ;
 wire \out_reg[11] ;
 wire \out_reg[12] ;
 wire \out_reg[13] ;
 wire \out_reg[14] ;
 wire \out_reg[15] ;
 wire \out_reg[1] ;
 wire \out_reg[2] ;
 wire \out_reg[3] ;
 wire \out_reg[4] ;
 wire \out_reg[5] ;
 wire \out_reg[6] ;
 wire \out_reg[7] ;
 wire \out_reg[8] ;
 wire \out_reg[9] ;
 wire \posit_add.in1[0] ;
 wire \posit_add.in1[10] ;
 wire \posit_add.in1[11] ;
 wire \posit_add.in1[12] ;
 wire \posit_add.in1[13] ;
 wire \posit_add.in1[14] ;
 wire \posit_add.in1[15] ;
 wire \posit_add.in1[1] ;
 wire \posit_add.in1[2] ;
 wire \posit_add.in1[3] ;
 wire \posit_add.in1[4] ;
 wire \posit_add.in1[5] ;
 wire \posit_add.in1[6] ;
 wire \posit_add.in1[7] ;
 wire \posit_add.in1[8] ;
 wire \posit_add.in1[9] ;
 wire \posit_add.in2[0] ;
 wire \posit_add.in2[10] ;
 wire \posit_add.in2[11] ;
 wire \posit_add.in2[12] ;
 wire \posit_add.in2[13] ;
 wire \posit_add.in2[14] ;
 wire \posit_add.in2[15] ;
 wire \posit_add.in2[1] ;
 wire \posit_add.in2[2] ;
 wire \posit_add.in2[3] ;
 wire \posit_add.in2[4] ;
 wire \posit_add.in2[5] ;
 wire \posit_add.in2[6] ;
 wire \posit_add.in2[7] ;
 wire \posit_add.in2[8] ;
 wire \posit_add.in2[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sky130_fd_sc_hd__buf_2 _4257_ (.A(net4),
    .X(_0635_));
 sky130_fd_sc_hd__or4_1 _4258_ (.A(\in_reg[5] ),
    .B(\in_reg[4] ),
    .C(\in_reg[7] ),
    .D(\in_reg[6] ),
    .X(_0646_));
 sky130_fd_sc_hd__or4_1 _4259_ (.A(\in_reg[1] ),
    .B(\in_reg[0] ),
    .C(\in_reg[3] ),
    .D(\in_reg[2] ),
    .X(_0657_));
 sky130_fd_sc_hd__or3_1 _4260_ (.A(\counter[2] ),
    .B(\counter[1] ),
    .C(\counter[0] ),
    .X(_0668_));
 sky130_fd_sc_hd__nor4b_2 _4261_ (.A(\counter[4] ),
    .B(mode),
    .C(_0668_),
    .D_N(\counter[3] ),
    .Y(_0679_));
 sky130_fd_sc_hd__o21ai_1 _4262_ (.A1(_0646_),
    .A2(_0657_),
    .B1(_0679_),
    .Y(_0690_));
 sky130_fd_sc_hd__clkbuf_4 _4263_ (.A(net1),
    .X(_0701_));
 sky130_fd_sc_hd__or3b_2 _4264_ (.A(_0635_),
    .B(_0690_),
    .C_N(_0701_),
    .X(_0712_));
 sky130_fd_sc_hd__mux2_1 _4265_ (.A0(\in_reg[0] ),
    .A1(\cmd[0] ),
    .S(_0712_),
    .X(_0723_));
 sky130_fd_sc_hd__clkbuf_1 _4266_ (.A(_0723_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _4267_ (.A0(\in_reg[6] ),
    .A1(\cmd[6] ),
    .S(_0712_),
    .X(_0744_));
 sky130_fd_sc_hd__clkbuf_1 _4268_ (.A(_0744_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _4269_ (.A0(\in_reg[7] ),
    .A1(\cmd[7] ),
    .S(_0712_),
    .X(_0765_));
 sky130_fd_sc_hd__clkbuf_1 _4270_ (.A(_0765_),
    .X(_0002_));
 sky130_fd_sc_hd__nor2b_1 _4271_ (.A(last_SCLK),
    .B_N(net2),
    .Y(_0786_));
 sky130_fd_sc_hd__nand2_1 _4272_ (.A(net1),
    .B(_0786_),
    .Y(_0797_));
 sky130_fd_sc_hd__or2_1 _4273_ (.A(net4),
    .B(_0797_),
    .X(_0808_));
 sky130_fd_sc_hd__clkbuf_4 _4274_ (.A(_0808_),
    .X(_0819_));
 sky130_fd_sc_hd__buf_4 _4275_ (.A(_0819_),
    .X(_0830_));
 sky130_fd_sc_hd__mux2_1 _4276_ (.A0(net3),
    .A1(\in_reg[0] ),
    .S(_0830_),
    .X(_0841_));
 sky130_fd_sc_hd__clkbuf_1 _4277_ (.A(_0841_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _4278_ (.A0(\in_reg[0] ),
    .A1(\in_reg[1] ),
    .S(_0830_),
    .X(_0862_));
 sky130_fd_sc_hd__clkbuf_1 _4279_ (.A(_0862_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _4280_ (.A0(\in_reg[1] ),
    .A1(\in_reg[2] ),
    .S(_0830_),
    .X(_0883_));
 sky130_fd_sc_hd__clkbuf_1 _4281_ (.A(_0883_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _4282_ (.A0(\in_reg[2] ),
    .A1(\in_reg[3] ),
    .S(_0830_),
    .X(_0904_));
 sky130_fd_sc_hd__clkbuf_1 _4283_ (.A(_0904_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _4284_ (.A0(\in_reg[3] ),
    .A1(\in_reg[4] ),
    .S(_0830_),
    .X(_0925_));
 sky130_fd_sc_hd__clkbuf_1 _4285_ (.A(_0925_),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _4286_ (.A0(\in_reg[4] ),
    .A1(\in_reg[5] ),
    .S(_0830_),
    .X(_0946_));
 sky130_fd_sc_hd__clkbuf_1 _4287_ (.A(_0946_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _4288_ (.A0(\in_reg[5] ),
    .A1(\in_reg[6] ),
    .S(_0830_),
    .X(_0967_));
 sky130_fd_sc_hd__clkbuf_1 _4289_ (.A(_0967_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _4290_ (.A0(\in_reg[6] ),
    .A1(\in_reg[7] ),
    .S(_0830_),
    .X(_0988_));
 sky130_fd_sc_hd__clkbuf_1 _4291_ (.A(_0988_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _4292_ (.A0(\in_reg[7] ),
    .A1(\in_reg[8] ),
    .S(_0830_),
    .X(_1009_));
 sky130_fd_sc_hd__clkbuf_1 _4293_ (.A(_1009_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _4294_ (.A0(\in_reg[8] ),
    .A1(\in_reg[9] ),
    .S(_0830_),
    .X(_1030_));
 sky130_fd_sc_hd__clkbuf_1 _4295_ (.A(_1030_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _4296_ (.A0(\in_reg[9] ),
    .A1(\in_reg[10] ),
    .S(_0819_),
    .X(_1051_));
 sky130_fd_sc_hd__clkbuf_1 _4297_ (.A(_1051_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _4298_ (.A0(\in_reg[10] ),
    .A1(\in_reg[11] ),
    .S(_0819_),
    .X(_1072_));
 sky130_fd_sc_hd__clkbuf_1 _4299_ (.A(_1072_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _4300_ (.A0(\in_reg[11] ),
    .A1(\in_reg[12] ),
    .S(_0819_),
    .X(_1093_));
 sky130_fd_sc_hd__clkbuf_1 _4301_ (.A(_1093_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _4302_ (.A0(\in_reg[12] ),
    .A1(\in_reg[13] ),
    .S(_0819_),
    .X(_1114_));
 sky130_fd_sc_hd__clkbuf_1 _4303_ (.A(_1114_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _4304_ (.A0(\in_reg[13] ),
    .A1(\in_reg[14] ),
    .S(_0819_),
    .X(_1135_));
 sky130_fd_sc_hd__clkbuf_1 _4305_ (.A(_1135_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _4306_ (.A0(\in_reg[14] ),
    .A1(\in_reg[15] ),
    .S(_0819_),
    .X(_1156_));
 sky130_fd_sc_hd__clkbuf_1 _4307_ (.A(_1156_),
    .X(_0018_));
 sky130_fd_sc_hd__buf_4 _4308_ (.A(_0701_),
    .X(_1177_));
 sky130_fd_sc_hd__mux2_1 _4309_ (.A0(last_SCLK),
    .A1(net2),
    .S(_1177_),
    .X(_1188_));
 sky130_fd_sc_hd__and2b_1 _4310_ (.A_N(_0635_),
    .B(_1188_),
    .X(_1199_));
 sky130_fd_sc_hd__clkbuf_1 _4311_ (.A(_1199_),
    .X(_0019_));
 sky130_fd_sc_hd__buf_2 _4312_ (.A(_0635_),
    .X(_1220_));
 sky130_fd_sc_hd__nor2b_2 _4313_ (.A(_0786_),
    .B_N(_0701_),
    .Y(_1231_));
 sky130_fd_sc_hd__clkbuf_4 _4314_ (.A(\posit_add.in1[15] ),
    .X(_1242_));
 sky130_fd_sc_hd__buf_4 _4315_ (.A(_1242_),
    .X(_1253_));
 sky130_fd_sc_hd__buf_2 _4316_ (.A(\posit_add.in2[15] ),
    .X(_1264_));
 sky130_fd_sc_hd__buf_4 _4317_ (.A(_1264_),
    .X(_1275_));
 sky130_fd_sc_hd__xor2_2 _4318_ (.A(_1253_),
    .B(_1275_),
    .X(_1286_));
 sky130_fd_sc_hd__clkbuf_4 _4319_ (.A(_1286_),
    .X(_1297_));
 sky130_fd_sc_hd__clkbuf_4 _4320_ (.A(_1297_),
    .X(_1308_));
 sky130_fd_sc_hd__clkbuf_2 _4321_ (.A(_1308_),
    .X(_1319_));
 sky130_fd_sc_hd__clkbuf_4 _4322_ (.A(_1319_),
    .X(_1330_));
 sky130_fd_sc_hd__or4_1 _4323_ (.A(\posit_add.in2[0] ),
    .B(\posit_add.in2[1] ),
    .C(\posit_add.in2[3] ),
    .D(\posit_add.in2[2] ),
    .X(_1341_));
 sky130_fd_sc_hd__buf_2 _4324_ (.A(_1341_),
    .X(_1352_));
 sky130_fd_sc_hd__or4_1 _4325_ (.A(\posit_add.in2[7] ),
    .B(\posit_add.in2[5] ),
    .C(\posit_add.in2[4] ),
    .D(\posit_add.in2[6] ),
    .X(_1363_));
 sky130_fd_sc_hd__clkbuf_2 _4326_ (.A(_1363_),
    .X(_1374_));
 sky130_fd_sc_hd__nor2_1 _4327_ (.A(_1352_),
    .B(_1374_),
    .Y(_1385_));
 sky130_fd_sc_hd__or4_1 _4328_ (.A(\posit_add.in2[11] ),
    .B(\posit_add.in2[9] ),
    .C(\posit_add.in2[8] ),
    .D(\posit_add.in2[10] ),
    .X(_1396_));
 sky130_fd_sc_hd__or2_1 _4329_ (.A(\posit_add.in2[13] ),
    .B(\posit_add.in2[12] ),
    .X(_1407_));
 sky130_fd_sc_hd__o41a_2 _4330_ (.A1(_1341_),
    .A2(_1374_),
    .A3(_1396_),
    .A4(_1407_),
    .B1(\posit_add.in2[15] ),
    .X(_1418_));
 sky130_fd_sc_hd__xnor2_4 _4331_ (.A(\posit_add.in2[14] ),
    .B(_1418_),
    .Y(_1429_));
 sky130_fd_sc_hd__o31a_1 _4332_ (.A1(_1341_),
    .A2(_1374_),
    .A3(_1396_),
    .B1(_1264_),
    .X(_1440_));
 sky130_fd_sc_hd__xnor2_4 _4333_ (.A(\posit_add.in2[12] ),
    .B(_1440_),
    .Y(_1451_));
 sky130_fd_sc_hd__or3_1 _4334_ (.A(\posit_add.in2[9] ),
    .B(\posit_add.in2[8] ),
    .C(\posit_add.in2[10] ),
    .X(_1462_));
 sky130_fd_sc_hd__o31a_1 _4335_ (.A1(_1341_),
    .A2(_1374_),
    .A3(_1462_),
    .B1(_1264_),
    .X(_1473_));
 sky130_fd_sc_hd__xnor2_4 _4336_ (.A(\posit_add.in2[11] ),
    .B(_1473_),
    .Y(_1484_));
 sky130_fd_sc_hd__or3_2 _4337_ (.A(_1429_),
    .B(_1451_),
    .C(_1484_),
    .X(_1495_));
 sky130_fd_sc_hd__buf_2 _4338_ (.A(_1429_),
    .X(_1506_));
 sky130_fd_sc_hd__nand3_2 _4339_ (.A(_1506_),
    .B(_1451_),
    .C(_1484_),
    .Y(_1517_));
 sky130_fd_sc_hd__o41a_2 _4340_ (.A1(\posit_add.in2[12] ),
    .A2(_1352_),
    .A3(_1374_),
    .A4(_1396_),
    .B1(_1264_),
    .X(_1528_));
 sky130_fd_sc_hd__xnor2_4 _4341_ (.A(\posit_add.in2[13] ),
    .B(_1528_),
    .Y(_1539_));
 sky130_fd_sc_hd__xor2_4 _4342_ (.A(_1429_),
    .B(_1539_),
    .X(_1550_));
 sky130_fd_sc_hd__a21oi_4 _4343_ (.A1(_1495_),
    .A2(_1517_),
    .B1(_1550_),
    .Y(_1561_));
 sky130_fd_sc_hd__o41a_2 _4344_ (.A1(\posit_add.in2[9] ),
    .A2(\posit_add.in2[8] ),
    .A3(_1352_),
    .A4(_1374_),
    .B1(_1264_),
    .X(_1572_));
 sky130_fd_sc_hd__xnor2_4 _4345_ (.A(\posit_add.in2[10] ),
    .B(_1572_),
    .Y(_1583_));
 sky130_fd_sc_hd__o31a_1 _4346_ (.A1(\posit_add.in2[8] ),
    .A2(_1352_),
    .A3(_1374_),
    .B1(_1264_),
    .X(_1594_));
 sky130_fd_sc_hd__xor2_2 _4347_ (.A(\posit_add.in2[9] ),
    .B(_1594_),
    .X(_1605_));
 sky130_fd_sc_hd__o21a_1 _4348_ (.A1(_1429_),
    .A2(_1583_),
    .B1(_1605_),
    .X(_1616_));
 sky130_fd_sc_hd__a21oi_1 _4349_ (.A1(_1506_),
    .A2(_1583_),
    .B1(_1605_),
    .Y(_1627_));
 sky130_fd_sc_hd__nor2_2 _4350_ (.A(_1616_),
    .B(_1627_),
    .Y(_1638_));
 sky130_fd_sc_hd__o21a_1 _4351_ (.A1(_1352_),
    .A2(_1374_),
    .B1(_1264_),
    .X(_1649_));
 sky130_fd_sc_hd__xnor2_2 _4352_ (.A(\posit_add.in2[8] ),
    .B(_1649_),
    .Y(_1660_));
 sky130_fd_sc_hd__o41a_2 _4353_ (.A1(\posit_add.in2[5] ),
    .A2(\posit_add.in2[4] ),
    .A3(\posit_add.in2[6] ),
    .A4(_1352_),
    .B1(_1264_),
    .X(_1671_));
 sky130_fd_sc_hd__xor2_4 _4354_ (.A(\posit_add.in2[7] ),
    .B(_1671_),
    .X(_1682_));
 sky130_fd_sc_hd__a21oi_1 _4355_ (.A1(_1506_),
    .A2(_1660_),
    .B1(_1682_),
    .Y(_1693_));
 sky130_fd_sc_hd__o21a_1 _4356_ (.A1(_1429_),
    .A2(_1660_),
    .B1(_1682_),
    .X(_1704_));
 sky130_fd_sc_hd__nor2_1 _4357_ (.A(_1693_),
    .B(_1704_),
    .Y(_1715_));
 sky130_fd_sc_hd__nand3_4 _4358_ (.A(_1561_),
    .B(_1638_),
    .C(_1715_),
    .Y(_1726_));
 sky130_fd_sc_hd__or2_2 _4359_ (.A(_1385_),
    .B(_1726_),
    .X(_1737_));
 sky130_fd_sc_hd__clkbuf_4 _4360_ (.A(_1737_),
    .X(_1748_));
 sky130_fd_sc_hd__nand2_1 _4361_ (.A(_1638_),
    .B(_1715_),
    .Y(_1759_));
 sky130_fd_sc_hd__or2_1 _4362_ (.A(\posit_add.in2[0] ),
    .B(\posit_add.in2[1] ),
    .X(_1770_));
 sky130_fd_sc_hd__clkbuf_4 _4363_ (.A(_1429_),
    .X(_1781_));
 sky130_fd_sc_hd__nand2_2 _4364_ (.A(_1275_),
    .B(_1770_),
    .Y(_1792_));
 sky130_fd_sc_hd__xor2_4 _4365_ (.A(\posit_add.in2[2] ),
    .B(_1792_),
    .X(_1803_));
 sky130_fd_sc_hd__nand2_1 _4366_ (.A(_1781_),
    .B(_1803_),
    .Y(_1814_));
 sky130_fd_sc_hd__o21a_2 _4367_ (.A1(\posit_add.in2[2] ),
    .A2(_1770_),
    .B1(_1275_),
    .X(_1825_));
 sky130_fd_sc_hd__xnor2_4 _4368_ (.A(\posit_add.in2[3] ),
    .B(_1825_),
    .Y(_1836_));
 sky130_fd_sc_hd__nand2_1 _4369_ (.A(_1275_),
    .B(_1352_),
    .Y(_1847_));
 sky130_fd_sc_hd__xor2_4 _4370_ (.A(\posit_add.in2[4] ),
    .B(_1847_),
    .X(_1858_));
 sky130_fd_sc_hd__nand2_1 _4371_ (.A(_1506_),
    .B(_1858_),
    .Y(_1869_));
 sky130_fd_sc_hd__xor2_1 _4372_ (.A(\posit_add.in2[3] ),
    .B(_1825_),
    .X(_1880_));
 sky130_fd_sc_hd__o21a_1 _4373_ (.A1(_1429_),
    .A2(_1858_),
    .B1(_1880_),
    .X(_1891_));
 sky130_fd_sc_hd__o21ai_2 _4374_ (.A1(\posit_add.in2[4] ),
    .A2(_1352_),
    .B1(_1264_),
    .Y(_1902_));
 sky130_fd_sc_hd__xnor2_4 _4375_ (.A(\posit_add.in2[5] ),
    .B(_1902_),
    .Y(_1913_));
 sky130_fd_sc_hd__xnor2_1 _4376_ (.A(_1429_),
    .B(_1913_),
    .Y(_1924_));
 sky130_fd_sc_hd__o31a_1 _4377_ (.A1(\posit_add.in2[5] ),
    .A2(\posit_add.in2[4] ),
    .A3(_1352_),
    .B1(_1264_),
    .X(_1935_));
 sky130_fd_sc_hd__xor2_4 _4378_ (.A(\posit_add.in2[6] ),
    .B(_1935_),
    .X(_1946_));
 sky130_fd_sc_hd__xnor2_1 _4379_ (.A(_1429_),
    .B(_1946_),
    .Y(_1957_));
 sky130_fd_sc_hd__a2111o_1 _4380_ (.A1(_1836_),
    .A2(_1869_),
    .B1(_1891_),
    .C1(_1924_),
    .D1(_1957_),
    .X(_1968_));
 sky130_fd_sc_hd__o21ba_1 _4381_ (.A1(_1770_),
    .A2(_1814_),
    .B1_N(_1968_),
    .X(_1979_));
 sky130_fd_sc_hd__o21ai_4 _4382_ (.A1(_1759_),
    .A2(_1979_),
    .B1(_1561_),
    .Y(_1990_));
 sky130_fd_sc_hd__and3_1 _4383_ (.A(_1561_),
    .B(_1638_),
    .C(_1715_),
    .X(_2001_));
 sky130_fd_sc_hd__clkbuf_2 _4384_ (.A(_2001_),
    .X(_2012_));
 sky130_fd_sc_hd__nand2_2 _4385_ (.A(\posit_add.in2[0] ),
    .B(_1275_),
    .Y(_2023_));
 sky130_fd_sc_hd__xor2_4 _4386_ (.A(\posit_add.in2[1] ),
    .B(_2023_),
    .X(_2034_));
 sky130_fd_sc_hd__or2_1 _4387_ (.A(_1506_),
    .B(_1803_),
    .X(_2045_));
 sky130_fd_sc_hd__nor2_1 _4388_ (.A(\posit_add.in2[0] ),
    .B(_2034_),
    .Y(_2056_));
 sky130_fd_sc_hd__o22a_1 _4389_ (.A1(_1814_),
    .A2(_2034_),
    .B1(_2045_),
    .B2(_2056_),
    .X(_2067_));
 sky130_fd_sc_hd__xor2_1 _4390_ (.A(_1506_),
    .B(_1913_),
    .X(_2078_));
 sky130_fd_sc_hd__or2_1 _4391_ (.A(_1506_),
    .B(_1858_),
    .X(_2089_));
 sky130_fd_sc_hd__a31o_1 _4392_ (.A1(_2078_),
    .A2(_2089_),
    .A3(_1869_),
    .B1(_1957_),
    .X(_2100_));
 sky130_fd_sc_hd__mux2_2 _4393_ (.A0(_2067_),
    .A1(_2100_),
    .S(_1968_),
    .X(_2111_));
 sky130_fd_sc_hd__a21o_1 _4394_ (.A1(_1495_),
    .A2(_1517_),
    .B1(_1550_),
    .X(_2122_));
 sky130_fd_sc_hd__xnor2_1 _4395_ (.A(_1506_),
    .B(_1660_),
    .Y(_2133_));
 sky130_fd_sc_hd__and2_1 _4396_ (.A(_1506_),
    .B(_1583_),
    .X(_2144_));
 sky130_fd_sc_hd__nor2_1 _4397_ (.A(_1781_),
    .B(_1583_),
    .Y(_2155_));
 sky130_fd_sc_hd__o32a_1 _4398_ (.A1(_1616_),
    .A2(_1627_),
    .A3(_2133_),
    .B1(_2144_),
    .B2(_2155_),
    .X(_2166_));
 sky130_fd_sc_hd__nor2_1 _4399_ (.A(_1781_),
    .B(_1451_),
    .Y(_2177_));
 sky130_fd_sc_hd__and2_1 _4400_ (.A(_1506_),
    .B(_1451_),
    .X(_2188_));
 sky130_fd_sc_hd__or3_1 _4401_ (.A(_2177_),
    .B(_2188_),
    .C(_1550_),
    .X(_2199_));
 sky130_fd_sc_hd__o21ai_2 _4402_ (.A1(_2122_),
    .A2(_2166_),
    .B1(_2199_),
    .Y(_2210_));
 sky130_fd_sc_hd__a21o_2 _4403_ (.A1(_2012_),
    .A2(_2111_),
    .B1(_2210_),
    .X(_2221_));
 sky130_fd_sc_hd__a211oi_1 _4404_ (.A1(_2012_),
    .A2(_2111_),
    .B1(_2210_),
    .C1(_1858_),
    .Y(_2232_));
 sky130_fd_sc_hd__nor2_1 _4405_ (.A(_2034_),
    .B(_2045_),
    .Y(_2243_));
 sky130_fd_sc_hd__and4_1 _4406_ (.A(\posit_add.in2[0] ),
    .B(_1781_),
    .C(_1803_),
    .D(_2034_),
    .X(_2254_));
 sky130_fd_sc_hd__nor2_1 _4407_ (.A(_1957_),
    .B(_1924_),
    .Y(_2265_));
 sky130_fd_sc_hd__o31ai_1 _4408_ (.A1(_1968_),
    .A2(_2243_),
    .A3(_2254_),
    .B1(_2265_),
    .Y(_2276_));
 sky130_fd_sc_hd__a21oi_1 _4409_ (.A1(_1495_),
    .A2(_1517_),
    .B1(_1638_),
    .Y(_2287_));
 sky130_fd_sc_hd__a211oi_2 _4410_ (.A1(_2012_),
    .A2(_2276_),
    .B1(_2287_),
    .C1(_1550_),
    .Y(_2298_));
 sky130_fd_sc_hd__buf_2 _4411_ (.A(_2298_),
    .X(_2309_));
 sky130_fd_sc_hd__a211o_1 _4412_ (.A1(_1913_),
    .A2(_2221_),
    .B1(_2232_),
    .C1(_2309_),
    .X(_2320_));
 sky130_fd_sc_hd__o22ai_1 _4413_ (.A1(_1814_),
    .A2(_2034_),
    .B1(_2045_),
    .B2(_2056_),
    .Y(_2331_));
 sky130_fd_sc_hd__a31oi_1 _4414_ (.A1(_2078_),
    .A2(_2089_),
    .A3(_1869_),
    .B1(_1957_),
    .Y(_2342_));
 sky130_fd_sc_hd__mux2_2 _4415_ (.A0(_2331_),
    .A1(_2342_),
    .S(_1968_),
    .X(_2353_));
 sky130_fd_sc_hd__o21a_2 _4416_ (.A1(_2122_),
    .A2(_2166_),
    .B1(_2199_),
    .X(_2364_));
 sky130_fd_sc_hd__xnor2_1 _4417_ (.A(\posit_add.in2[2] ),
    .B(_1792_),
    .Y(_2375_));
 sky130_fd_sc_hd__o211a_1 _4418_ (.A1(_1726_),
    .A2(_2353_),
    .B1(_2364_),
    .C1(_2375_),
    .X(_2386_));
 sky130_fd_sc_hd__a211o_1 _4419_ (.A1(_2012_),
    .A2(_2276_),
    .B1(_2287_),
    .C1(_1550_),
    .X(_2397_));
 sky130_fd_sc_hd__buf_2 _4420_ (.A(_2397_),
    .X(_2408_));
 sky130_fd_sc_hd__a211o_1 _4421_ (.A1(_1880_),
    .A2(_2221_),
    .B1(_2386_),
    .C1(_2408_),
    .X(_2419_));
 sky130_fd_sc_hd__xnor2_1 _4422_ (.A(\posit_add.in2[1] ),
    .B(_2023_),
    .Y(_2430_));
 sky130_fd_sc_hd__a21oi_1 _4423_ (.A1(_2012_),
    .A2(_2111_),
    .B1(_2210_),
    .Y(_2441_));
 sky130_fd_sc_hd__buf_4 _4424_ (.A(_2441_),
    .X(_2452_));
 sky130_fd_sc_hd__a211o_1 _4425_ (.A1(_2012_),
    .A2(_2111_),
    .B1(_2210_),
    .C1(\posit_add.in2[0] ),
    .X(_2463_));
 sky130_fd_sc_hd__o21a_1 _4426_ (.A1(_1759_),
    .A2(_1979_),
    .B1(_1561_),
    .X(_2474_));
 sky130_fd_sc_hd__buf_2 _4427_ (.A(_2474_),
    .X(_2485_));
 sky130_fd_sc_hd__o2111a_1 _4428_ (.A1(_2430_),
    .A2(_2452_),
    .B1(_2463_),
    .C1(_2408_),
    .D1(_2485_),
    .X(_2496_));
 sky130_fd_sc_hd__a31o_4 _4429_ (.A1(_1990_),
    .A2(_2320_),
    .A3(_2419_),
    .B1(_2496_),
    .X(_2507_));
 sky130_fd_sc_hd__nand2_1 _4430_ (.A(_1748_),
    .B(_2507_),
    .Y(_2518_));
 sky130_fd_sc_hd__buf_4 _4431_ (.A(_2518_),
    .X(_2529_));
 sky130_fd_sc_hd__buf_2 _4432_ (.A(_2529_),
    .X(_2540_));
 sky130_fd_sc_hd__or4_2 _4433_ (.A(\posit_add.in1[0] ),
    .B(\posit_add.in1[3] ),
    .C(\posit_add.in1[2] ),
    .D(\posit_add.in1[1] ),
    .X(_2551_));
 sky130_fd_sc_hd__or4_1 _4434_ (.A(\posit_add.in1[6] ),
    .B(\posit_add.in1[5] ),
    .C(\posit_add.in1[4] ),
    .D(_2551_),
    .X(_2562_));
 sky130_fd_sc_hd__or4_2 _4435_ (.A(\posit_add.in1[9] ),
    .B(\posit_add.in1[8] ),
    .C(\posit_add.in1[7] ),
    .D(_2562_),
    .X(_2573_));
 sky130_fd_sc_hd__or2_1 _4436_ (.A(\posit_add.in1[13] ),
    .B(\posit_add.in1[12] ),
    .X(_2584_));
 sky130_fd_sc_hd__o41a_2 _4437_ (.A1(\posit_add.in1[11] ),
    .A2(\posit_add.in1[10] ),
    .A3(_2573_),
    .A4(_2584_),
    .B1(_1242_),
    .X(_2595_));
 sky130_fd_sc_hd__xnor2_4 _4438_ (.A(\posit_add.in1[14] ),
    .B(_2595_),
    .Y(_2606_));
 sky130_fd_sc_hd__or2_1 _4439_ (.A(\posit_add.in1[7] ),
    .B(_2562_),
    .X(_2617_));
 sky130_fd_sc_hd__nand2_1 _4440_ (.A(_1242_),
    .B(_2617_),
    .Y(_2628_));
 sky130_fd_sc_hd__xor2_2 _4441_ (.A(\posit_add.in1[8] ),
    .B(_2628_),
    .X(_2639_));
 sky130_fd_sc_hd__and2_1 _4442_ (.A(_2606_),
    .B(_2639_),
    .X(_2650_));
 sky130_fd_sc_hd__buf_4 _4443_ (.A(_2606_),
    .X(_2661_));
 sky130_fd_sc_hd__nor2_1 _4444_ (.A(_2661_),
    .B(_2639_),
    .Y(_2672_));
 sky130_fd_sc_hd__and2_1 _4445_ (.A(_1242_),
    .B(_2562_),
    .X(_2683_));
 sky130_fd_sc_hd__xor2_2 _4446_ (.A(\posit_add.in1[7] ),
    .B(_2683_),
    .X(_2694_));
 sky130_fd_sc_hd__mux2_1 _4447_ (.A0(_2650_),
    .A1(_2672_),
    .S(_2694_),
    .X(_2705_));
 sky130_fd_sc_hd__nand2_2 _4448_ (.A(_1242_),
    .B(_2573_),
    .Y(_2716_));
 sky130_fd_sc_hd__xnor2_4 _4449_ (.A(\posit_add.in1[10] ),
    .B(_2716_),
    .Y(_2727_));
 sky130_fd_sc_hd__xnor2_2 _4450_ (.A(_2606_),
    .B(_2727_),
    .Y(_2738_));
 sky130_fd_sc_hd__o21a_1 _4451_ (.A1(\posit_add.in1[8] ),
    .A2(_2617_),
    .B1(_1242_),
    .X(_2749_));
 sky130_fd_sc_hd__xor2_4 _4452_ (.A(\posit_add.in1[9] ),
    .B(_2749_),
    .X(_2760_));
 sky130_fd_sc_hd__xnor2_1 _4453_ (.A(_2661_),
    .B(_2760_),
    .Y(_2771_));
 sky130_fd_sc_hd__nor2_1 _4454_ (.A(_2738_),
    .B(_2771_),
    .Y(_2782_));
 sky130_fd_sc_hd__nand2_1 _4455_ (.A(_2705_),
    .B(_2782_),
    .Y(_2793_));
 sky130_fd_sc_hd__inv_2 _4456_ (.A(_2793_),
    .Y(_2804_));
 sky130_fd_sc_hd__o31a_1 _4457_ (.A1(\posit_add.in1[5] ),
    .A2(\posit_add.in1[4] ),
    .A3(_2551_),
    .B1(_1253_),
    .X(_2815_));
 sky130_fd_sc_hd__xor2_4 _4458_ (.A(\posit_add.in1[6] ),
    .B(_2815_),
    .X(_2826_));
 sky130_fd_sc_hd__xor2_1 _4459_ (.A(_2661_),
    .B(_2826_),
    .X(_2837_));
 sky130_fd_sc_hd__o21ai_2 _4460_ (.A1(\posit_add.in1[4] ),
    .A2(_2551_),
    .B1(_1242_),
    .Y(_2848_));
 sky130_fd_sc_hd__xnor2_4 _4461_ (.A(\posit_add.in1[5] ),
    .B(_2848_),
    .Y(_2859_));
 sky130_fd_sc_hd__xor2_1 _4462_ (.A(_2661_),
    .B(_2859_),
    .X(_2870_));
 sky130_fd_sc_hd__nand2_1 _4463_ (.A(_2837_),
    .B(_2870_),
    .Y(_2881_));
 sky130_fd_sc_hd__nand2_1 _4464_ (.A(_1242_),
    .B(_2551_),
    .Y(_2892_));
 sky130_fd_sc_hd__xnor2_4 _4465_ (.A(\posit_add.in1[4] ),
    .B(_2892_),
    .Y(_2903_));
 sky130_fd_sc_hd__xnor2_1 _4466_ (.A(_2661_),
    .B(_2903_),
    .Y(_2914_));
 sky130_fd_sc_hd__o31a_1 _4467_ (.A1(\posit_add.in1[0] ),
    .A2(\posit_add.in1[2] ),
    .A3(\posit_add.in1[1] ),
    .B1(\posit_add.in1[15] ),
    .X(_2925_));
 sky130_fd_sc_hd__xor2_4 _4468_ (.A(\posit_add.in1[3] ),
    .B(_2925_),
    .X(_2936_));
 sky130_fd_sc_hd__xnor2_1 _4469_ (.A(_2661_),
    .B(_2936_),
    .Y(_2947_));
 sky130_fd_sc_hd__or2_1 _4470_ (.A(_2914_),
    .B(_2947_),
    .X(_2958_));
 sky130_fd_sc_hd__clkbuf_4 _4471_ (.A(\posit_add.in1[0] ),
    .X(_2969_));
 sky130_fd_sc_hd__inv_4 _4472_ (.A(_2661_),
    .Y(_2980_));
 sky130_fd_sc_hd__or4_1 _4473_ (.A(_2969_),
    .B(\posit_add.in1[2] ),
    .C(\posit_add.in1[1] ),
    .D(_2980_),
    .X(_2991_));
 sky130_fd_sc_hd__or3b_2 _4474_ (.A(_2881_),
    .B(_2958_),
    .C_N(_2991_),
    .X(_3002_));
 sky130_fd_sc_hd__or3_2 _4475_ (.A(\posit_add.in1[11] ),
    .B(\posit_add.in1[10] ),
    .C(_2573_),
    .X(_3013_));
 sky130_fd_sc_hd__o21a_1 _4476_ (.A1(\posit_add.in1[12] ),
    .A2(_3013_),
    .B1(_1253_),
    .X(_3024_));
 sky130_fd_sc_hd__xnor2_4 _4477_ (.A(\posit_add.in1[13] ),
    .B(_3024_),
    .Y(_3035_));
 sky130_fd_sc_hd__xnor2_4 _4478_ (.A(_2980_),
    .B(_3035_),
    .Y(_3046_));
 sky130_fd_sc_hd__nand2_1 _4479_ (.A(_1253_),
    .B(_3013_),
    .Y(_3057_));
 sky130_fd_sc_hd__xnor2_4 _4480_ (.A(\posit_add.in1[12] ),
    .B(_3057_),
    .Y(_3068_));
 sky130_fd_sc_hd__xnor2_4 _4481_ (.A(_2980_),
    .B(_3068_),
    .Y(_3079_));
 sky130_fd_sc_hd__o21ai_2 _4482_ (.A1(\posit_add.in1[10] ),
    .A2(_2573_),
    .B1(_1253_),
    .Y(_3090_));
 sky130_fd_sc_hd__xnor2_4 _4483_ (.A(\posit_add.in1[11] ),
    .B(_3090_),
    .Y(_3101_));
 sky130_fd_sc_hd__xor2_2 _4484_ (.A(_2661_),
    .B(_3101_),
    .X(_3112_));
 sky130_fd_sc_hd__nand2_1 _4485_ (.A(_3079_),
    .B(_3112_),
    .Y(_3123_));
 sky130_fd_sc_hd__or2_2 _4486_ (.A(_3046_),
    .B(_3123_),
    .X(_3134_));
 sky130_fd_sc_hd__a21o_1 _4487_ (.A1(_2804_),
    .A2(_3002_),
    .B1(_3134_),
    .X(_3145_));
 sky130_fd_sc_hd__buf_2 _4488_ (.A(_3145_),
    .X(_3156_));
 sky130_fd_sc_hd__buf_4 _4489_ (.A(_3156_),
    .X(_3167_));
 sky130_fd_sc_hd__o21ai_2 _4490_ (.A1(\posit_add.in1[0] ),
    .A2(\posit_add.in1[1] ),
    .B1(_1242_),
    .Y(_3178_));
 sky130_fd_sc_hd__xnor2_4 _4491_ (.A(\posit_add.in1[2] ),
    .B(_3178_),
    .Y(_3189_));
 sky130_fd_sc_hd__xor2_1 _4492_ (.A(_2606_),
    .B(_3189_),
    .X(_3199_));
 sky130_fd_sc_hd__or2b_1 _4493_ (.A(_2969_),
    .B_N(\posit_add.in1[1] ),
    .X(_3210_));
 sky130_fd_sc_hd__nand2_1 _4494_ (.A(\posit_add.in1[0] ),
    .B(_1242_),
    .Y(_3221_));
 sky130_fd_sc_hd__xnor2_4 _4495_ (.A(\posit_add.in1[1] ),
    .B(_3221_),
    .Y(_3232_));
 sky130_fd_sc_hd__mux2_1 _4496_ (.A0(_3210_),
    .A1(_3232_),
    .S(_2606_),
    .X(_3243_));
 sky130_fd_sc_hd__a21oi_1 _4497_ (.A1(_3199_),
    .A2(_3243_),
    .B1(_2947_),
    .Y(_3253_));
 sky130_fd_sc_hd__o21ai_1 _4498_ (.A1(_2914_),
    .A2(_3253_),
    .B1(_2870_),
    .Y(_3264_));
 sky130_fd_sc_hd__a21oi_2 _4499_ (.A1(_2837_),
    .A2(_3264_),
    .B1(_2793_),
    .Y(_3275_));
 sky130_fd_sc_hd__nor3_2 _4500_ (.A(_2650_),
    .B(_2672_),
    .C(_2771_),
    .Y(_3285_));
 sky130_fd_sc_hd__o31ai_4 _4501_ (.A1(_2738_),
    .A2(_3275_),
    .A3(_3285_),
    .B1(_3112_),
    .Y(_3296_));
 sky130_fd_sc_hd__a21o_2 _4502_ (.A1(_3079_),
    .A2(_3296_),
    .B1(_3046_),
    .X(_3307_));
 sky130_fd_sc_hd__buf_2 _4503_ (.A(_3307_),
    .X(_3318_));
 sky130_fd_sc_hd__clkbuf_8 _4504_ (.A(_2661_),
    .X(_3328_));
 sky130_fd_sc_hd__xnor2_4 _4505_ (.A(_3328_),
    .B(_3068_),
    .Y(_3339_));
 sky130_fd_sc_hd__o31a_4 _4506_ (.A1(_2738_),
    .A2(_3275_),
    .A3(_3285_),
    .B1(_3112_),
    .X(_3349_));
 sky130_fd_sc_hd__xnor2_4 _4507_ (.A(_3328_),
    .B(_3035_),
    .Y(_3360_));
 sky130_fd_sc_hd__o211a_1 _4508_ (.A1(_3339_),
    .A2(_3349_),
    .B1(_2826_),
    .C1(_3360_),
    .X(_3371_));
 sky130_fd_sc_hd__xor2_1 _4509_ (.A(_2661_),
    .B(_3232_),
    .X(_3381_));
 sky130_fd_sc_hd__o211a_1 _4510_ (.A1(_2969_),
    .A2(_2980_),
    .B1(_3199_),
    .C1(_3381_),
    .X(_3392_));
 sky130_fd_sc_hd__nor2_1 _4511_ (.A(_2958_),
    .B(_3392_),
    .Y(_3403_));
 sky130_fd_sc_hd__o21ai_1 _4512_ (.A1(_2881_),
    .A2(_3403_),
    .B1(_2705_),
    .Y(_3414_));
 sky130_fd_sc_hd__a21oi_2 _4513_ (.A1(_2782_),
    .A2(_3414_),
    .B1(_3123_),
    .Y(_3424_));
 sky130_fd_sc_hd__nor2_1 _4514_ (.A(_3046_),
    .B(_3424_),
    .Y(_3435_));
 sky130_fd_sc_hd__clkbuf_4 _4515_ (.A(_3435_),
    .X(_3446_));
 sky130_fd_sc_hd__a211o_1 _4516_ (.A1(_2859_),
    .A2(_3318_),
    .B1(_3371_),
    .C1(_3446_),
    .X(_3456_));
 sky130_fd_sc_hd__o211a_1 _4517_ (.A1(_3339_),
    .A2(_3349_),
    .B1(_2903_),
    .C1(_3360_),
    .X(_3467_));
 sky130_fd_sc_hd__or2_2 _4518_ (.A(_3046_),
    .B(_3424_),
    .X(_3477_));
 sky130_fd_sc_hd__clkbuf_4 _4519_ (.A(_3477_),
    .X(_3488_));
 sky130_fd_sc_hd__a211o_1 _4520_ (.A1(_2936_),
    .A2(_3318_),
    .B1(_3467_),
    .C1(_3488_),
    .X(_3498_));
 sky130_fd_sc_hd__nand2_2 _4521_ (.A(_3456_),
    .B(_3498_),
    .Y(_3509_));
 sky130_fd_sc_hd__a21oi_4 _4522_ (.A1(_2804_),
    .A2(_3002_),
    .B1(_3134_),
    .Y(_3520_));
 sky130_fd_sc_hd__a21oi_4 _4523_ (.A1(_3079_),
    .A2(_3296_),
    .B1(_3046_),
    .Y(_3530_));
 sky130_fd_sc_hd__nand3_1 _4524_ (.A(_2969_),
    .B(_3446_),
    .C(_3530_),
    .Y(_3541_));
 sky130_fd_sc_hd__a211o_1 _4525_ (.A1(_3079_),
    .A2(_3296_),
    .B1(_3189_),
    .C1(_3046_),
    .X(_3552_));
 sky130_fd_sc_hd__o211ai_2 _4526_ (.A1(_3232_),
    .A2(_3530_),
    .B1(_3552_),
    .C1(_3488_),
    .Y(_3562_));
 sky130_fd_sc_hd__and3_1 _4527_ (.A(_3520_),
    .B(_3541_),
    .C(_3562_),
    .X(_3573_));
 sky130_fd_sc_hd__and3b_1 _4528_ (.A_N(_3134_),
    .B(_2617_),
    .C(_2804_),
    .X(_3583_));
 sky130_fd_sc_hd__clkbuf_4 _4529_ (.A(_3583_),
    .X(_3594_));
 sky130_fd_sc_hd__a211o_1 _4530_ (.A1(_3167_),
    .A2(_3509_),
    .B1(_3573_),
    .C1(_3594_),
    .X(_3604_));
 sky130_fd_sc_hd__clkbuf_4 _4531_ (.A(_3604_),
    .X(_3615_));
 sky130_fd_sc_hd__and3_1 _4532_ (.A(_2485_),
    .B(_2320_),
    .C(_2419_),
    .X(_3625_));
 sky130_fd_sc_hd__clkbuf_4 _4533_ (.A(_2221_),
    .X(_3635_));
 sky130_fd_sc_hd__inv_2 _4534_ (.A(_1660_),
    .Y(_3643_));
 sky130_fd_sc_hd__o211a_1 _4535_ (.A1(_1726_),
    .A2(_2353_),
    .B1(_2364_),
    .C1(_3643_),
    .X(_3651_));
 sky130_fd_sc_hd__a211o_1 _4536_ (.A1(_1605_),
    .A2(_3635_),
    .B1(_3651_),
    .C1(_2309_),
    .X(_3659_));
 sky130_fd_sc_hd__o211a_1 _4537_ (.A1(_1726_),
    .A2(_2353_),
    .B1(_2364_),
    .C1(_1946_),
    .X(_3665_));
 sky130_fd_sc_hd__a211o_1 _4538_ (.A1(_1682_),
    .A2(_3635_),
    .B1(_3665_),
    .C1(_2408_),
    .X(_3671_));
 sky130_fd_sc_hd__nor2_4 _4539_ (.A(_1385_),
    .B(_1726_),
    .Y(_3678_));
 sky130_fd_sc_hd__a31o_1 _4540_ (.A1(_1990_),
    .A2(_3659_),
    .A3(_3671_),
    .B1(_3678_),
    .X(_3684_));
 sky130_fd_sc_hd__clkbuf_4 _4541_ (.A(_1990_),
    .X(_3690_));
 sky130_fd_sc_hd__o21a_1 _4542_ (.A1(_2430_),
    .A2(_2452_),
    .B1(_2463_),
    .X(_3696_));
 sky130_fd_sc_hd__a31o_1 _4543_ (.A1(_3690_),
    .A2(_2408_),
    .A3(_3696_),
    .B1(_1737_),
    .X(_3698_));
 sky130_fd_sc_hd__o21ai_4 _4544_ (.A1(_3625_),
    .A2(_3684_),
    .B1(_3698_),
    .Y(_3699_));
 sky130_fd_sc_hd__clkbuf_4 _4545_ (.A(_3699_),
    .X(_3700_));
 sky130_fd_sc_hd__clkbuf_4 _4546_ (.A(_3700_),
    .X(_3701_));
 sky130_fd_sc_hd__a211o_4 _4547_ (.A1(_3541_),
    .A2(_3562_),
    .B1(_3594_),
    .C1(_3520_),
    .X(_3702_));
 sky130_fd_sc_hd__clkbuf_4 _4548_ (.A(_3702_),
    .X(_3703_));
 sky130_fd_sc_hd__nor2_1 _4549_ (.A(_3701_),
    .B(_3703_),
    .Y(_3704_));
 sky130_fd_sc_hd__o211a_1 _4550_ (.A1(_1726_),
    .A2(_2353_),
    .B1(_2364_),
    .C1(_1682_),
    .X(_3705_));
 sky130_fd_sc_hd__a211o_1 _4551_ (.A1(_3643_),
    .A2(_2221_),
    .B1(_3705_),
    .C1(_2309_),
    .X(_3706_));
 sky130_fd_sc_hd__o211a_1 _4552_ (.A1(_1726_),
    .A2(_2353_),
    .B1(_2364_),
    .C1(_1913_),
    .X(_3707_));
 sky130_fd_sc_hd__a211o_1 _4553_ (.A1(_1946_),
    .A2(_2221_),
    .B1(_3707_),
    .C1(_2408_),
    .X(_3708_));
 sky130_fd_sc_hd__and3_1 _4554_ (.A(\posit_add.in2[0] ),
    .B(_2408_),
    .C(_2221_),
    .X(_3709_));
 sky130_fd_sc_hd__a31o_1 _4555_ (.A1(_1737_),
    .A2(_3706_),
    .A3(_3708_),
    .B1(_3709_),
    .X(_3710_));
 sky130_fd_sc_hd__nand2_1 _4556_ (.A(_2485_),
    .B(_1737_),
    .Y(_3711_));
 sky130_fd_sc_hd__o211a_1 _4557_ (.A1(_1726_),
    .A2(_2353_),
    .B1(_2364_),
    .C1(_2034_),
    .X(_3712_));
 sky130_fd_sc_hd__a211o_1 _4558_ (.A1(_1803_),
    .A2(_2221_),
    .B1(_3712_),
    .C1(_2408_),
    .X(_3713_));
 sky130_fd_sc_hd__o211a_1 _4559_ (.A1(_1726_),
    .A2(_2353_),
    .B1(_2364_),
    .C1(_1836_),
    .X(_3714_));
 sky130_fd_sc_hd__a211o_1 _4560_ (.A1(_1858_),
    .A2(_2221_),
    .B1(_3714_),
    .C1(_2298_),
    .X(_3715_));
 sky130_fd_sc_hd__and2_1 _4561_ (.A(_3713_),
    .B(_3715_),
    .X(_3716_));
 sky130_fd_sc_hd__o2bb2a_2 _4562_ (.A1_N(_3690_),
    .A2_N(_3710_),
    .B1(_3711_),
    .B2(_3716_),
    .X(_3717_));
 sky130_fd_sc_hd__buf_2 _4563_ (.A(_3717_),
    .X(_3718_));
 sky130_fd_sc_hd__clkbuf_4 _4564_ (.A(_3718_),
    .X(_3719_));
 sky130_fd_sc_hd__or3b_1 _4565_ (.A(_2793_),
    .B(_3134_),
    .C_N(_2617_),
    .X(_3720_));
 sky130_fd_sc_hd__clkbuf_4 _4566_ (.A(_3720_),
    .X(_3721_));
 sky130_fd_sc_hd__clkbuf_4 _4567_ (.A(_3721_),
    .X(_3722_));
 sky130_fd_sc_hd__a211o_1 _4568_ (.A1(_3079_),
    .A2(_3296_),
    .B1(_3232_),
    .C1(_3046_),
    .X(_3723_));
 sky130_fd_sc_hd__o2111a_1 _4569_ (.A1(_2969_),
    .A2(_3530_),
    .B1(_3723_),
    .C1(_3167_),
    .D1(_3488_),
    .X(_3724_));
 sky130_fd_sc_hd__nand2_2 _4570_ (.A(_3722_),
    .B(_3724_),
    .Y(_3725_));
 sky130_fd_sc_hd__buf_2 _4571_ (.A(_3725_),
    .X(_3726_));
 sky130_fd_sc_hd__nor2_1 _4572_ (.A(_3719_),
    .B(_3726_),
    .Y(_3727_));
 sky130_fd_sc_hd__nand2_2 _4573_ (.A(_3704_),
    .B(_3727_),
    .Y(_3728_));
 sky130_fd_sc_hd__buf_4 _4574_ (.A(_3678_),
    .X(_3729_));
 sky130_fd_sc_hd__o211a_1 _4575_ (.A1(_2430_),
    .A2(_2441_),
    .B1(_2463_),
    .C1(_2298_),
    .X(_3730_));
 sky130_fd_sc_hd__a211o_1 _4576_ (.A1(_2012_),
    .A2(_2111_),
    .B1(_2210_),
    .C1(_2375_),
    .X(_3731_));
 sky130_fd_sc_hd__o211a_1 _4577_ (.A1(_1880_),
    .A2(_2452_),
    .B1(_3731_),
    .C1(_2397_),
    .X(_3732_));
 sky130_fd_sc_hd__o21ai_2 _4578_ (.A1(_3730_),
    .A2(_3732_),
    .B1(_3690_),
    .Y(_3733_));
 sky130_fd_sc_hd__or2_1 _4579_ (.A(_3729_),
    .B(_3733_),
    .X(_3734_));
 sky130_fd_sc_hd__clkbuf_4 _4580_ (.A(_3734_),
    .X(_3735_));
 sky130_fd_sc_hd__clkbuf_4 _4581_ (.A(_2485_),
    .X(_3736_));
 sky130_fd_sc_hd__or4b_1 _4582_ (.A(_3736_),
    .B(_2309_),
    .C(_3729_),
    .D_N(_3696_),
    .X(_3737_));
 sky130_fd_sc_hd__clkbuf_2 _4583_ (.A(_3737_),
    .X(_3738_));
 sky130_fd_sc_hd__clkbuf_4 _4584_ (.A(_3738_),
    .X(_3739_));
 sky130_fd_sc_hd__o211a_1 _4585_ (.A1(_3339_),
    .A2(_3349_),
    .B1(_2694_),
    .C1(_3360_),
    .X(_3740_));
 sky130_fd_sc_hd__a211o_1 _4586_ (.A1(_2826_),
    .A2(_3318_),
    .B1(_3740_),
    .C1(_3446_),
    .X(_3741_));
 sky130_fd_sc_hd__o211a_1 _4587_ (.A1(_3339_),
    .A2(_3349_),
    .B1(_2859_),
    .C1(_3360_),
    .X(_3742_));
 sky130_fd_sc_hd__a211o_1 _4588_ (.A1(_2903_),
    .A2(_3307_),
    .B1(_3742_),
    .C1(_3477_),
    .X(_3743_));
 sky130_fd_sc_hd__nand2_1 _4589_ (.A(_3741_),
    .B(_3743_),
    .Y(_3744_));
 sky130_fd_sc_hd__o211a_1 _4590_ (.A1(_3339_),
    .A2(_3349_),
    .B1(_2936_),
    .C1(_3360_),
    .X(_3745_));
 sky130_fd_sc_hd__a211o_2 _4591_ (.A1(_3189_),
    .A2(_3318_),
    .B1(_3745_),
    .C1(_3446_),
    .X(_3746_));
 sky130_fd_sc_hd__o211a_1 _4592_ (.A1(_3339_),
    .A2(_3349_),
    .B1(_3232_),
    .C1(_3360_),
    .X(_3747_));
 sky130_fd_sc_hd__a211o_2 _4593_ (.A1(_2969_),
    .A2(_3318_),
    .B1(_3747_),
    .C1(_3488_),
    .X(_3748_));
 sky130_fd_sc_hd__a21oi_1 _4594_ (.A1(_3746_),
    .A2(_3748_),
    .B1(_3167_),
    .Y(_3749_));
 sky130_fd_sc_hd__a211o_4 _4595_ (.A1(_3167_),
    .A2(_3744_),
    .B1(_3749_),
    .C1(_3594_),
    .X(_3750_));
 sky130_fd_sc_hd__a211o_1 _4596_ (.A1(_2903_),
    .A2(_3318_),
    .B1(_3742_),
    .C1(_3446_),
    .X(_3751_));
 sky130_fd_sc_hd__a211o_1 _4597_ (.A1(_3189_),
    .A2(_3318_),
    .B1(_3745_),
    .C1(_3488_),
    .X(_3752_));
 sky130_fd_sc_hd__o2111a_1 _4598_ (.A1(_2969_),
    .A2(_3530_),
    .B1(_3723_),
    .C1(_3520_),
    .D1(_3488_),
    .X(_3753_));
 sky130_fd_sc_hd__a31o_1 _4599_ (.A1(_3156_),
    .A2(_3751_),
    .A3(_3752_),
    .B1(_3753_),
    .X(_3754_));
 sky130_fd_sc_hd__nand2_2 _4600_ (.A(_3722_),
    .B(_3754_),
    .Y(_3755_));
 sky130_fd_sc_hd__nor4_2 _4601_ (.A(_3735_),
    .B(_3739_),
    .C(_3750_),
    .D(_3755_),
    .Y(_3756_));
 sky130_fd_sc_hd__a211o_1 _4602_ (.A1(_1682_),
    .A2(_2221_),
    .B1(_3665_),
    .C1(_2298_),
    .X(_3757_));
 sky130_fd_sc_hd__a211o_1 _4603_ (.A1(_1913_),
    .A2(_2221_),
    .B1(_2232_),
    .C1(_2408_),
    .X(_3758_));
 sky130_fd_sc_hd__a21o_1 _4604_ (.A1(_3757_),
    .A2(_3758_),
    .B1(_2485_),
    .X(_3759_));
 sky130_fd_sc_hd__o31a_1 _4605_ (.A1(_1990_),
    .A2(_3730_),
    .A3(_3732_),
    .B1(_1737_),
    .X(_3760_));
 sky130_fd_sc_hd__nand2_2 _4606_ (.A(_3759_),
    .B(_3760_),
    .Y(_3761_));
 sky130_fd_sc_hd__clkbuf_4 _4607_ (.A(_3761_),
    .X(_3762_));
 sky130_fd_sc_hd__clkbuf_4 _4608_ (.A(_3762_),
    .X(_3763_));
 sky130_fd_sc_hd__or2_1 _4609_ (.A(_3763_),
    .B(_3702_),
    .X(_3764_));
 sky130_fd_sc_hd__inv_2 _4610_ (.A(\posit_add.in2[0] ),
    .Y(_3765_));
 sky130_fd_sc_hd__or3_1 _4611_ (.A(_3765_),
    .B(_2408_),
    .C(_2452_),
    .X(_3766_));
 sky130_fd_sc_hd__a211o_1 _4612_ (.A1(_1803_),
    .A2(_3635_),
    .B1(_3712_),
    .C1(_2309_),
    .X(_3767_));
 sky130_fd_sc_hd__and2_1 _4613_ (.A(_3766_),
    .B(_3767_),
    .X(_3768_));
 sky130_fd_sc_hd__nor2_1 _4614_ (.A(_3736_),
    .B(_3768_),
    .Y(_3769_));
 sky130_fd_sc_hd__nand2_4 _4615_ (.A(_1748_),
    .B(_3769_),
    .Y(_3770_));
 sky130_fd_sc_hd__clkbuf_4 _4616_ (.A(_3770_),
    .X(_3771_));
 sky130_fd_sc_hd__buf_4 _4617_ (.A(_3594_),
    .X(_3772_));
 sky130_fd_sc_hd__a2111oi_2 _4618_ (.A1(_3167_),
    .A2(_3744_),
    .B1(_3749_),
    .C1(_3771_),
    .D1(_3772_),
    .Y(_3773_));
 sky130_fd_sc_hd__o31a_2 _4619_ (.A1(_3765_),
    .A2(_2309_),
    .A3(_2452_),
    .B1(_2474_),
    .X(_3774_));
 sky130_fd_sc_hd__a311oi_4 _4620_ (.A1(_1990_),
    .A2(_3713_),
    .A3(_3715_),
    .B1(_3774_),
    .C1(_3678_),
    .Y(_3775_));
 sky130_fd_sc_hd__clkbuf_4 _4621_ (.A(_3775_),
    .X(_3776_));
 sky130_fd_sc_hd__and3_1 _4622_ (.A(_3722_),
    .B(_3754_),
    .C(_3776_),
    .X(_3777_));
 sky130_fd_sc_hd__xor2_1 _4623_ (.A(_3773_),
    .B(_3777_),
    .X(_3778_));
 sky130_fd_sc_hd__xnor2_1 _4624_ (.A(_3764_),
    .B(_3778_),
    .Y(_3779_));
 sky130_fd_sc_hd__xnor2_1 _4625_ (.A(_3756_),
    .B(_3779_),
    .Y(_3780_));
 sky130_fd_sc_hd__nor2_1 _4626_ (.A(_3763_),
    .B(_3725_),
    .Y(_3781_));
 sky130_fd_sc_hd__a2111o_2 _4627_ (.A1(_3167_),
    .A2(_3509_),
    .B1(_3771_),
    .C1(_3573_),
    .D1(_3594_),
    .X(_3782_));
 sky130_fd_sc_hd__a211o_1 _4628_ (.A1(_2936_),
    .A2(_3307_),
    .B1(_3467_),
    .C1(_3435_),
    .X(_3783_));
 sky130_fd_sc_hd__o211a_1 _4629_ (.A1(_3339_),
    .A2(_3349_),
    .B1(_3189_),
    .C1(_3360_),
    .X(_3784_));
 sky130_fd_sc_hd__a211o_1 _4630_ (.A1(_3232_),
    .A2(_3307_),
    .B1(_3784_),
    .C1(_3477_),
    .X(_3785_));
 sky130_fd_sc_hd__o2111a_1 _4631_ (.A1(_3339_),
    .A2(_3349_),
    .B1(_3424_),
    .C1(_2969_),
    .D1(_3360_),
    .X(_3786_));
 sky130_fd_sc_hd__and2_1 _4632_ (.A(_3520_),
    .B(_3786_),
    .X(_3787_));
 sky130_fd_sc_hd__a31o_1 _4633_ (.A1(_3156_),
    .A2(_3783_),
    .A3(_3785_),
    .B1(_3787_),
    .X(_3788_));
 sky130_fd_sc_hd__and3_1 _4634_ (.A(_3721_),
    .B(_3776_),
    .C(_3788_),
    .X(_3789_));
 sky130_fd_sc_hd__xnor2_1 _4635_ (.A(_3782_),
    .B(_3789_),
    .Y(_3790_));
 sky130_fd_sc_hd__a311o_2 _4636_ (.A1(_3690_),
    .A2(_3713_),
    .A3(_3715_),
    .B1(_3774_),
    .C1(_3678_),
    .X(_3791_));
 sky130_fd_sc_hd__buf_4 _4637_ (.A(_3791_),
    .X(_3792_));
 sky130_fd_sc_hd__buf_2 _4638_ (.A(_3792_),
    .X(_3793_));
 sky130_fd_sc_hd__nand2_1 _4639_ (.A(_3721_),
    .B(_3788_),
    .Y(_3794_));
 sky130_fd_sc_hd__clkbuf_4 _4640_ (.A(_3794_),
    .X(_3795_));
 sky130_fd_sc_hd__or3_1 _4641_ (.A(_3793_),
    .B(_3795_),
    .C(_3782_),
    .X(_3796_));
 sky130_fd_sc_hd__a21bo_1 _4642_ (.A1(_3781_),
    .A2(_3790_),
    .B1_N(_3796_),
    .X(_3797_));
 sky130_fd_sc_hd__and2b_1 _4643_ (.A_N(_3780_),
    .B(_3797_),
    .X(_3798_));
 sky130_fd_sc_hd__a21o_1 _4644_ (.A1(_3756_),
    .A2(_3779_),
    .B1(_3798_),
    .X(_3799_));
 sky130_fd_sc_hd__clkbuf_4 _4645_ (.A(_3719_),
    .X(_3800_));
 sky130_fd_sc_hd__o21a_2 _4646_ (.A1(_3625_),
    .A2(_3684_),
    .B1(_3698_),
    .X(_3801_));
 sky130_fd_sc_hd__buf_4 _4647_ (.A(_3801_),
    .X(_3802_));
 sky130_fd_sc_hd__and2_1 _4648_ (.A(_3722_),
    .B(_3724_),
    .X(_3803_));
 sky130_fd_sc_hd__buf_4 _4649_ (.A(_3803_),
    .X(_3804_));
 sky130_fd_sc_hd__nand2_1 _4650_ (.A(_3802_),
    .B(_3804_),
    .Y(_3805_));
 sky130_fd_sc_hd__o21ai_1 _4651_ (.A1(_3800_),
    .A2(_3703_),
    .B1(_3805_),
    .Y(_3806_));
 sky130_fd_sc_hd__and3_1 _4652_ (.A(_3728_),
    .B(_3799_),
    .C(_3806_),
    .X(_3807_));
 sky130_fd_sc_hd__a211o_1 _4653_ (.A1(_1946_),
    .A2(_3635_),
    .B1(_3707_),
    .C1(_2309_),
    .X(_3808_));
 sky130_fd_sc_hd__a211o_1 _4654_ (.A1(_2012_),
    .A2(_2111_),
    .B1(_2210_),
    .C1(_1836_),
    .X(_3809_));
 sky130_fd_sc_hd__o211ai_2 _4655_ (.A1(_1858_),
    .A2(_2452_),
    .B1(_3809_),
    .C1(_2309_),
    .Y(_3810_));
 sky130_fd_sc_hd__a21o_1 _4656_ (.A1(_3808_),
    .A2(_3810_),
    .B1(_2485_),
    .X(_3811_));
 sky130_fd_sc_hd__a31oi_2 _4657_ (.A1(_2485_),
    .A2(_3766_),
    .A3(_3767_),
    .B1(_3678_),
    .Y(_3812_));
 sky130_fd_sc_hd__nand2_2 _4658_ (.A(_3811_),
    .B(_3812_),
    .Y(_3813_));
 sky130_fd_sc_hd__buf_2 _4659_ (.A(_3813_),
    .X(_3814_));
 sky130_fd_sc_hd__clkbuf_4 _4660_ (.A(_3814_),
    .X(_3815_));
 sky130_fd_sc_hd__clkbuf_4 _4661_ (.A(_3815_),
    .X(_3816_));
 sky130_fd_sc_hd__buf_4 _4662_ (.A(_3755_),
    .X(_3817_));
 sky130_fd_sc_hd__nor2_1 _4663_ (.A(_3816_),
    .B(_3817_),
    .Y(_3818_));
 sky130_fd_sc_hd__xnor2_1 _4664_ (.A(\posit_add.in1[8] ),
    .B(_2628_),
    .Y(_3819_));
 sky130_fd_sc_hd__o211a_1 _4665_ (.A1(_3339_),
    .A2(_3349_),
    .B1(_3819_),
    .C1(_3360_),
    .X(_3820_));
 sky130_fd_sc_hd__a211o_1 _4666_ (.A1(_2694_),
    .A2(_3318_),
    .B1(_3820_),
    .C1(_3488_),
    .X(_3821_));
 sky130_fd_sc_hd__o211a_1 _4667_ (.A1(_3339_),
    .A2(_3349_),
    .B1(_2727_),
    .C1(_3360_),
    .X(_3822_));
 sky130_fd_sc_hd__a211o_1 _4668_ (.A1(_2760_),
    .A2(_3318_),
    .B1(_3822_),
    .C1(_3446_),
    .X(_3823_));
 sky130_fd_sc_hd__nand2_1 _4669_ (.A(_3821_),
    .B(_3823_),
    .Y(_3824_));
 sky130_fd_sc_hd__mux2_1 _4670_ (.A0(_3509_),
    .A1(_3824_),
    .S(_3156_),
    .X(_3825_));
 sky130_fd_sc_hd__a21o_1 _4671_ (.A1(_3541_),
    .A2(_3562_),
    .B1(_3520_),
    .X(_3826_));
 sky130_fd_sc_hd__mux2_4 _4672_ (.A0(_3825_),
    .A1(_3826_),
    .S(_3594_),
    .X(_3827_));
 sky130_fd_sc_hd__clkbuf_4 _4673_ (.A(_3735_),
    .X(_3828_));
 sky130_fd_sc_hd__or2_1 _4674_ (.A(_3827_),
    .B(_3828_),
    .X(_3829_));
 sky130_fd_sc_hd__clkbuf_4 _4675_ (.A(_2408_),
    .X(_3830_));
 sky130_fd_sc_hd__and4_1 _4676_ (.A(_3690_),
    .B(_3830_),
    .C(_1748_),
    .D(_3696_),
    .X(_3831_));
 sky130_fd_sc_hd__clkbuf_4 _4677_ (.A(_3831_),
    .X(_3832_));
 sky130_fd_sc_hd__a211o_1 _4678_ (.A1(_2694_),
    .A2(_3307_),
    .B1(_3820_),
    .C1(_3435_),
    .X(_3833_));
 sky130_fd_sc_hd__a211o_1 _4679_ (.A1(_2859_),
    .A2(_3307_),
    .B1(_3371_),
    .C1(_3477_),
    .X(_3834_));
 sky130_fd_sc_hd__a21o_1 _4680_ (.A1(_3833_),
    .A2(_3834_),
    .B1(_3520_),
    .X(_3835_));
 sky130_fd_sc_hd__a21o_1 _4681_ (.A1(_3783_),
    .A2(_3785_),
    .B1(_3156_),
    .X(_3836_));
 sky130_fd_sc_hd__and3_1 _4682_ (.A(_3594_),
    .B(_3156_),
    .C(_3786_),
    .X(_3837_));
 sky130_fd_sc_hd__a31o_4 _4683_ (.A1(_3721_),
    .A2(_3835_),
    .A3(_3836_),
    .B1(_3837_),
    .X(_3838_));
 sky130_fd_sc_hd__nand2_1 _4684_ (.A(_3832_),
    .B(_3838_),
    .Y(_3839_));
 sky130_fd_sc_hd__a31oi_4 _4685_ (.A1(_3722_),
    .A2(_3835_),
    .A3(_3836_),
    .B1(_3837_),
    .Y(_3840_));
 sky130_fd_sc_hd__o22a_1 _4686_ (.A1(_3827_),
    .A2(_3739_),
    .B1(_3840_),
    .B2(_3828_),
    .X(_3841_));
 sky130_fd_sc_hd__o21ba_1 _4687_ (.A1(_3829_),
    .A2(_3839_),
    .B1_N(_3841_),
    .X(_3842_));
 sky130_fd_sc_hd__xnor2_1 _4688_ (.A(_3818_),
    .B(_3842_),
    .Y(_3843_));
 sky130_fd_sc_hd__nor2_1 _4689_ (.A(_3828_),
    .B(_3750_),
    .Y(_3844_));
 sky130_fd_sc_hd__buf_2 _4690_ (.A(_3739_),
    .X(_3845_));
 sky130_fd_sc_hd__a21oi_2 _4691_ (.A1(_3751_),
    .A2(_3752_),
    .B1(_3167_),
    .Y(_3846_));
 sky130_fd_sc_hd__a21o_1 _4692_ (.A1(_2826_),
    .A2(_3307_),
    .B1(_3740_),
    .X(_3847_));
 sky130_fd_sc_hd__a211o_1 _4693_ (.A1(_3079_),
    .A2(_3296_),
    .B1(_2760_),
    .C1(_3046_),
    .X(_3848_));
 sky130_fd_sc_hd__o211a_1 _4694_ (.A1(_3819_),
    .A2(_3530_),
    .B1(_3848_),
    .C1(_3477_),
    .X(_3849_));
 sky130_fd_sc_hd__a21o_1 _4695_ (.A1(_3446_),
    .A2(_3847_),
    .B1(_3849_),
    .X(_3850_));
 sky130_fd_sc_hd__nor2_1 _4696_ (.A(_3520_),
    .B(_3850_),
    .Y(_3851_));
 sky130_fd_sc_hd__nand2_1 _4697_ (.A(_3772_),
    .B(_3724_),
    .Y(_3852_));
 sky130_fd_sc_hd__o31a_1 _4698_ (.A1(_3772_),
    .A2(_3846_),
    .A3(_3851_),
    .B1(_3852_),
    .X(_3853_));
 sky130_fd_sc_hd__nor2_1 _4699_ (.A(_3845_),
    .B(_3853_),
    .Y(_3854_));
 sky130_fd_sc_hd__o31ai_4 _4700_ (.A1(_3772_),
    .A2(_3846_),
    .A3(_3851_),
    .B1(_3852_),
    .Y(_3855_));
 sky130_fd_sc_hd__and3_1 _4701_ (.A(_3832_),
    .B(_3855_),
    .C(_3844_),
    .X(_3856_));
 sky130_fd_sc_hd__o21ba_1 _4702_ (.A1(_3844_),
    .A2(_3854_),
    .B1_N(_3856_),
    .X(_3857_));
 sky130_fd_sc_hd__nor2_1 _4703_ (.A(_3816_),
    .B(_3795_),
    .Y(_3858_));
 sky130_fd_sc_hd__nand2_1 _4704_ (.A(_3857_),
    .B(_3858_),
    .Y(_3859_));
 sky130_fd_sc_hd__or2_1 _4705_ (.A(_3843_),
    .B(_3859_),
    .X(_3860_));
 sky130_fd_sc_hd__nand2_1 _4706_ (.A(_3843_),
    .B(_3859_),
    .Y(_3861_));
 sky130_fd_sc_hd__and2_1 _4707_ (.A(_3860_),
    .B(_3861_),
    .X(_3862_));
 sky130_fd_sc_hd__and2_1 _4708_ (.A(_3759_),
    .B(_3760_),
    .X(_3863_));
 sky130_fd_sc_hd__buf_2 _4709_ (.A(_3863_),
    .X(_3864_));
 sky130_fd_sc_hd__buf_2 _4710_ (.A(_3864_),
    .X(_3865_));
 sky130_fd_sc_hd__clkbuf_4 _4711_ (.A(_3865_),
    .X(_3866_));
 sky130_fd_sc_hd__and4_1 _4712_ (.A(_3721_),
    .B(_3156_),
    .C(_3746_),
    .D(_3748_),
    .X(_3867_));
 sky130_fd_sc_hd__clkbuf_4 _4713_ (.A(_3867_),
    .X(_3868_));
 sky130_fd_sc_hd__nand2_1 _4714_ (.A(_3866_),
    .B(_3868_),
    .Y(_3869_));
 sky130_fd_sc_hd__o22a_1 _4715_ (.A1(_3771_),
    .A2(_3840_),
    .B1(_3615_),
    .B2(_3793_),
    .X(_3870_));
 sky130_fd_sc_hd__nand2_1 _4716_ (.A(_3776_),
    .B(_3838_),
    .Y(_3871_));
 sky130_fd_sc_hd__or2_1 _4717_ (.A(_3871_),
    .B(_3782_),
    .X(_3872_));
 sky130_fd_sc_hd__o21ai_1 _4718_ (.A1(_3869_),
    .A2(_3870_),
    .B1(_3872_),
    .Y(_3873_));
 sky130_fd_sc_hd__or2_1 _4719_ (.A(_3793_),
    .B(_3750_),
    .X(_3874_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4720_ (.A(_3874_),
    .X(_3875_));
 sky130_fd_sc_hd__or2_1 _4721_ (.A(_2485_),
    .B(_3768_),
    .X(_3876_));
 sky130_fd_sc_hd__nor2_1 _4722_ (.A(_3729_),
    .B(_3876_),
    .Y(_3877_));
 sky130_fd_sc_hd__clkbuf_4 _4723_ (.A(_3877_),
    .X(_3878_));
 sky130_fd_sc_hd__nand2_1 _4724_ (.A(_3878_),
    .B(_3855_),
    .Y(_3879_));
 sky130_fd_sc_hd__xor2_1 _4725_ (.A(_3875_),
    .B(_3879_),
    .X(_3880_));
 sky130_fd_sc_hd__clkbuf_4 _4726_ (.A(_3866_),
    .X(_3881_));
 sky130_fd_sc_hd__a31oi_4 _4727_ (.A1(_3145_),
    .A2(_3783_),
    .A3(_3785_),
    .B1(_3787_),
    .Y(_3882_));
 sky130_fd_sc_hd__nor2_4 _4728_ (.A(_3772_),
    .B(_3882_),
    .Y(_3883_));
 sky130_fd_sc_hd__nand2_1 _4729_ (.A(_3881_),
    .B(_3883_),
    .Y(_3884_));
 sky130_fd_sc_hd__xnor2_1 _4730_ (.A(_3880_),
    .B(_3884_),
    .Y(_3885_));
 sky130_fd_sc_hd__xnor2_1 _4731_ (.A(_3856_),
    .B(_3885_),
    .Y(_3886_));
 sky130_fd_sc_hd__xnor2_1 _4732_ (.A(_3873_),
    .B(_3886_),
    .Y(_3887_));
 sky130_fd_sc_hd__nand2_1 _4733_ (.A(_3862_),
    .B(_3887_),
    .Y(_3888_));
 sky130_fd_sc_hd__or2_1 _4734_ (.A(_3862_),
    .B(_3887_),
    .X(_3889_));
 sky130_fd_sc_hd__nand2_1 _4735_ (.A(_3888_),
    .B(_3889_),
    .Y(_3890_));
 sky130_fd_sc_hd__xnor2_1 _4736_ (.A(_3857_),
    .B(_3858_),
    .Y(_3891_));
 sky130_fd_sc_hd__nor2_4 _4737_ (.A(_3729_),
    .B(_3733_),
    .Y(_3892_));
 sky130_fd_sc_hd__clkbuf_4 _4738_ (.A(_3892_),
    .X(_3893_));
 sky130_fd_sc_hd__a211oi_4 _4739_ (.A1(_3167_),
    .A2(_3509_),
    .B1(_3573_),
    .C1(_3772_),
    .Y(_3894_));
 sky130_fd_sc_hd__nand2_1 _4740_ (.A(_3893_),
    .B(_3894_),
    .Y(_3895_));
 sky130_fd_sc_hd__and4_1 _4741_ (.A(_3893_),
    .B(_3832_),
    .C(_3838_),
    .D(_3894_),
    .X(_3896_));
 sky130_fd_sc_hd__a21o_1 _4742_ (.A1(_3839_),
    .A2(_3895_),
    .B1(_3896_),
    .X(_3897_));
 sky130_fd_sc_hd__a21oi_2 _4743_ (.A1(_3808_),
    .A2(_3810_),
    .B1(_2485_),
    .Y(_3898_));
 sky130_fd_sc_hd__a31o_1 _4744_ (.A1(_2485_),
    .A2(_3766_),
    .A3(_3767_),
    .B1(_3678_),
    .X(_3899_));
 sky130_fd_sc_hd__nor2_4 _4745_ (.A(_3898_),
    .B(_3899_),
    .Y(_3900_));
 sky130_fd_sc_hd__buf_4 _4746_ (.A(_3900_),
    .X(_3901_));
 sky130_fd_sc_hd__nand2_1 _4747_ (.A(_3901_),
    .B(_3868_),
    .Y(_3902_));
 sky130_fd_sc_hd__or2_1 _4748_ (.A(_3897_),
    .B(_3902_),
    .X(_3903_));
 sky130_fd_sc_hd__o21ba_1 _4749_ (.A1(_3871_),
    .A2(_3782_),
    .B1_N(_3870_),
    .X(_3904_));
 sky130_fd_sc_hd__xnor2_1 _4750_ (.A(_3869_),
    .B(_3904_),
    .Y(_3905_));
 sky130_fd_sc_hd__xnor2_1 _4751_ (.A(_3896_),
    .B(_3905_),
    .Y(_3906_));
 sky130_fd_sc_hd__nor2_2 _4752_ (.A(_3772_),
    .B(_3826_),
    .Y(_3907_));
 sky130_fd_sc_hd__and2_1 _4753_ (.A(_3773_),
    .B(_3777_),
    .X(_3908_));
 sky130_fd_sc_hd__a31o_1 _4754_ (.A1(_3881_),
    .A2(_3907_),
    .A3(_3778_),
    .B1(_3908_),
    .X(_3909_));
 sky130_fd_sc_hd__xor2_1 _4755_ (.A(_3906_),
    .B(_3909_),
    .X(_3910_));
 sky130_fd_sc_hd__xor2_1 _4756_ (.A(_3891_),
    .B(_3903_),
    .X(_3911_));
 sky130_fd_sc_hd__or2b_1 _4757_ (.A(_3910_),
    .B_N(_3911_),
    .X(_3912_));
 sky130_fd_sc_hd__o21ai_2 _4758_ (.A1(_3891_),
    .A2(_3903_),
    .B1(_3912_),
    .Y(_3913_));
 sky130_fd_sc_hd__xor2_2 _4759_ (.A(_3890_),
    .B(_3913_),
    .X(_3914_));
 sky130_fd_sc_hd__nand2_1 _4760_ (.A(_3896_),
    .B(_3905_),
    .Y(_3915_));
 sky130_fd_sc_hd__or2b_1 _4761_ (.A(_3906_),
    .B_N(_3909_),
    .X(_3916_));
 sky130_fd_sc_hd__and3_1 _4762_ (.A(_3736_),
    .B(_3808_),
    .C(_3810_),
    .X(_3917_));
 sky130_fd_sc_hd__a21oi_1 _4763_ (.A1(_3643_),
    .A2(_3635_),
    .B1(_3705_),
    .Y(_3918_));
 sky130_fd_sc_hd__xnor2_1 _4764_ (.A(\posit_add.in2[9] ),
    .B(_1594_),
    .Y(_3919_));
 sky130_fd_sc_hd__mux2_1 _4765_ (.A0(_1583_),
    .A1(_3919_),
    .S(_2452_),
    .X(_3920_));
 sky130_fd_sc_hd__mux2_1 _4766_ (.A0(_3918_),
    .A1(_3920_),
    .S(_3830_),
    .X(_3921_));
 sky130_fd_sc_hd__o21ai_1 _4767_ (.A1(_3736_),
    .A2(_3921_),
    .B1(_1748_),
    .Y(_3922_));
 sky130_fd_sc_hd__a2bb2o_2 _4768_ (.A1_N(_3917_),
    .A2_N(_3922_),
    .B1(_3876_),
    .B2(_3729_),
    .X(_3923_));
 sky130_fd_sc_hd__clkbuf_4 _4769_ (.A(_3923_),
    .X(_3924_));
 sky130_fd_sc_hd__clkbuf_4 _4770_ (.A(_3924_),
    .X(_3925_));
 sky130_fd_sc_hd__nor2_1 _4771_ (.A(_3925_),
    .B(_3726_),
    .Y(_3926_));
 sky130_fd_sc_hd__or2_1 _4772_ (.A(_3924_),
    .B(_3702_),
    .X(_3927_));
 sky130_fd_sc_hd__or2_1 _4773_ (.A(_3927_),
    .B(_3805_),
    .X(_3928_));
 sky130_fd_sc_hd__o21a_1 _4774_ (.A1(_3926_),
    .A2(_3704_),
    .B1(_3928_),
    .X(_3929_));
 sky130_fd_sc_hd__nand4_4 _4775_ (.A(_3722_),
    .B(_3167_),
    .C(_3746_),
    .D(_3748_),
    .Y(_3930_));
 sky130_fd_sc_hd__nor2_1 _4776_ (.A(_3719_),
    .B(_3930_),
    .Y(_3931_));
 sky130_fd_sc_hd__xnor2_1 _4777_ (.A(_3929_),
    .B(_3931_),
    .Y(_3932_));
 sky130_fd_sc_hd__a21oi_1 _4778_ (.A1(_3915_),
    .A2(_3916_),
    .B1(_3932_),
    .Y(_3933_));
 sky130_fd_sc_hd__and3_1 _4779_ (.A(_3915_),
    .B(_3916_),
    .C(_3932_),
    .X(_3934_));
 sky130_fd_sc_hd__or2_1 _4780_ (.A(_3933_),
    .B(_3934_),
    .X(_3935_));
 sky130_fd_sc_hd__xnor2_2 _4781_ (.A(_3935_),
    .B(_3728_),
    .Y(_3936_));
 sky130_fd_sc_hd__xnor2_2 _4782_ (.A(_3914_),
    .B(_3936_),
    .Y(_3937_));
 sky130_fd_sc_hd__nand2_1 _4783_ (.A(_3728_),
    .B(_3806_),
    .Y(_3938_));
 sky130_fd_sc_hd__xnor2_1 _4784_ (.A(_3799_),
    .B(_3938_),
    .Y(_3939_));
 sky130_fd_sc_hd__xnor2_1 _4785_ (.A(_3910_),
    .B(_3911_),
    .Y(_3940_));
 sky130_fd_sc_hd__xnor2_1 _4786_ (.A(_3897_),
    .B(_3902_),
    .Y(_3941_));
 sky130_fd_sc_hd__or2_1 _4787_ (.A(_3739_),
    .B(_3750_),
    .X(_3942_));
 sky130_fd_sc_hd__and2_1 _4788_ (.A(_3722_),
    .B(_3754_),
    .X(_3943_));
 sky130_fd_sc_hd__nand2_1 _4789_ (.A(_3893_),
    .B(_3943_),
    .Y(_3944_));
 sky130_fd_sc_hd__a21o_1 _4790_ (.A1(_3942_),
    .A2(_3944_),
    .B1(_3756_),
    .X(_3945_));
 sky130_fd_sc_hd__or3_1 _4791_ (.A(_3816_),
    .B(_3702_),
    .C(_3945_),
    .X(_3946_));
 sky130_fd_sc_hd__xor2_1 _4792_ (.A(_3780_),
    .B(_3797_),
    .X(_3947_));
 sky130_fd_sc_hd__xnor2_1 _4793_ (.A(_3941_),
    .B(_3946_),
    .Y(_3948_));
 sky130_fd_sc_hd__nor2_1 _4794_ (.A(_3947_),
    .B(_3948_),
    .Y(_3949_));
 sky130_fd_sc_hd__o21ba_1 _4795_ (.A1(_3941_),
    .A2(_3946_),
    .B1_N(_3949_),
    .X(_3950_));
 sky130_fd_sc_hd__xnor2_1 _4796_ (.A(_3940_),
    .B(_3950_),
    .Y(_3951_));
 sky130_fd_sc_hd__or2b_1 _4797_ (.A(_3950_),
    .B_N(_3940_),
    .X(_3952_));
 sky130_fd_sc_hd__a21bo_1 _4798_ (.A1(_3939_),
    .A2(_3951_),
    .B1_N(_3952_),
    .X(_3953_));
 sky130_fd_sc_hd__xnor2_1 _4799_ (.A(_3937_),
    .B(_3953_),
    .Y(_3954_));
 sky130_fd_sc_hd__xnor2_1 _4800_ (.A(_3807_),
    .B(_3954_),
    .Y(_3955_));
 sky130_fd_sc_hd__or4_1 _4801_ (.A(_3735_),
    .B(_3739_),
    .C(_3604_),
    .D(_3794_),
    .X(_3956_));
 sky130_fd_sc_hd__xnor2_1 _4802_ (.A(_3781_),
    .B(_3790_),
    .Y(_3957_));
 sky130_fd_sc_hd__xnor2_1 _4803_ (.A(_3956_),
    .B(_3957_),
    .Y(_3958_));
 sky130_fd_sc_hd__nand2_1 _4804_ (.A(_3878_),
    .B(_3868_),
    .Y(_3959_));
 sky130_fd_sc_hd__or3_1 _4805_ (.A(_3793_),
    .B(_3817_),
    .C(_3959_),
    .X(_3960_));
 sky130_fd_sc_hd__or2_1 _4806_ (.A(_3958_),
    .B(_3960_),
    .X(_3961_));
 sky130_fd_sc_hd__o21a_1 _4807_ (.A1(_3956_),
    .A2(_3957_),
    .B1(_3961_),
    .X(_3962_));
 sky130_fd_sc_hd__or3_1 _4808_ (.A(_3800_),
    .B(_3726_),
    .C(_3962_),
    .X(_3963_));
 sky130_fd_sc_hd__xnor2_1 _4809_ (.A(_3939_),
    .B(_3951_),
    .Y(_3964_));
 sky130_fd_sc_hd__xnor2_1 _4810_ (.A(_3727_),
    .B(_3962_),
    .Y(_3965_));
 sky130_fd_sc_hd__and2_1 _4811_ (.A(_3947_),
    .B(_3948_),
    .X(_3966_));
 sky130_fd_sc_hd__or2_1 _4812_ (.A(_3949_),
    .B(_3966_),
    .X(_3967_));
 sky130_fd_sc_hd__xnor2_1 _4813_ (.A(_3958_),
    .B(_3960_),
    .Y(_3968_));
 sky130_fd_sc_hd__nor2_1 _4814_ (.A(_3815_),
    .B(_3702_),
    .Y(_3969_));
 sky130_fd_sc_hd__xnor2_1 _4815_ (.A(_3945_),
    .B(_3969_),
    .Y(_3970_));
 sky130_fd_sc_hd__nor2_1 _4816_ (.A(_3816_),
    .B(_3726_),
    .Y(_3971_));
 sky130_fd_sc_hd__o22a_1 _4817_ (.A1(_3739_),
    .A2(_3604_),
    .B1(_3794_),
    .B2(_3735_),
    .X(_3972_));
 sky130_fd_sc_hd__and2b_1 _4818_ (.A_N(_3972_),
    .B(_3956_),
    .X(_3973_));
 sky130_fd_sc_hd__and2_1 _4819_ (.A(_3971_),
    .B(_3973_),
    .X(_3974_));
 sky130_fd_sc_hd__xnor2_1 _4820_ (.A(_3970_),
    .B(_3974_),
    .Y(_3975_));
 sky130_fd_sc_hd__nand2_1 _4821_ (.A(_3970_),
    .B(_3974_),
    .Y(_3976_));
 sky130_fd_sc_hd__o21ai_1 _4822_ (.A1(_3968_),
    .A2(_3975_),
    .B1(_3976_),
    .Y(_3977_));
 sky130_fd_sc_hd__xnor2_1 _4823_ (.A(_3967_),
    .B(_3977_),
    .Y(_3978_));
 sky130_fd_sc_hd__and2b_1 _4824_ (.A_N(_3967_),
    .B(_3977_),
    .X(_3979_));
 sky130_fd_sc_hd__a21oi_1 _4825_ (.A1(_3965_),
    .A2(_3978_),
    .B1(_3979_),
    .Y(_3980_));
 sky130_fd_sc_hd__xnor2_1 _4826_ (.A(_3964_),
    .B(_3980_),
    .Y(_3981_));
 sky130_fd_sc_hd__or2_1 _4827_ (.A(_3964_),
    .B(_3980_),
    .X(_3982_));
 sky130_fd_sc_hd__o21a_1 _4828_ (.A1(_3963_),
    .A2(_3981_),
    .B1(_3982_),
    .X(_3983_));
 sky130_fd_sc_hd__xnor2_1 _4829_ (.A(_3955_),
    .B(_3983_),
    .Y(_3984_));
 sky130_fd_sc_hd__o32a_1 _4830_ (.A1(_2540_),
    .A2(_3615_),
    .A3(_3984_),
    .B1(_3983_),
    .B2(_3955_),
    .X(_3985_));
 sky130_fd_sc_hd__buf_6 _4831_ (.A(_3894_),
    .X(_3986_));
 sky130_fd_sc_hd__nand2_1 _4832_ (.A(_3901_),
    .B(_3986_),
    .Y(_3987_));
 sky130_fd_sc_hd__clkbuf_4 _4833_ (.A(_3853_),
    .X(_3988_));
 sky130_fd_sc_hd__nor3_4 _4834_ (.A(\posit_add.in1[14] ),
    .B(_3013_),
    .C(_2584_),
    .Y(_3989_));
 sky130_fd_sc_hd__o22a_1 _4835_ (.A1(_3828_),
    .A2(_3988_),
    .B1(_3989_),
    .B2(_3845_),
    .X(_3990_));
 sky130_fd_sc_hd__a21o_1 _4836_ (.A1(_3893_),
    .A2(_3854_),
    .B1(_3990_),
    .X(_3991_));
 sky130_fd_sc_hd__xor2_1 _4837_ (.A(_3987_),
    .B(_3991_),
    .X(_3992_));
 sky130_fd_sc_hd__and2_1 _4838_ (.A(_3818_),
    .B(_3842_),
    .X(_3993_));
 sky130_fd_sc_hd__nand2_1 _4839_ (.A(_3992_),
    .B(_3993_),
    .Y(_3994_));
 sky130_fd_sc_hd__or2_1 _4840_ (.A(_3992_),
    .B(_3993_),
    .X(_3995_));
 sky130_fd_sc_hd__nand2_1 _4841_ (.A(_3994_),
    .B(_3995_),
    .Y(_3996_));
 sky130_fd_sc_hd__nor2_1 _4842_ (.A(_3875_),
    .B(_3879_),
    .Y(_3997_));
 sky130_fd_sc_hd__a31o_1 _4843_ (.A1(_3881_),
    .A2(_3883_),
    .A3(_3880_),
    .B1(_3997_),
    .X(_3998_));
 sky130_fd_sc_hd__or3_1 _4844_ (.A(_3827_),
    .B(_3771_),
    .C(_3871_),
    .X(_3999_));
 sky130_fd_sc_hd__o21ai_1 _4845_ (.A1(_3827_),
    .A2(_3771_),
    .B1(_3871_),
    .Y(_4000_));
 sky130_fd_sc_hd__nor2_1 _4846_ (.A(_3763_),
    .B(_3817_),
    .Y(_4001_));
 sky130_fd_sc_hd__and3_1 _4847_ (.A(_3999_),
    .B(_4000_),
    .C(_4001_),
    .X(_4002_));
 sky130_fd_sc_hd__a21oi_1 _4848_ (.A1(_3999_),
    .A2(_4000_),
    .B1(_4001_),
    .Y(_4003_));
 sky130_fd_sc_hd__or2_1 _4849_ (.A(_4002_),
    .B(_4003_),
    .X(_4004_));
 sky130_fd_sc_hd__or3_1 _4850_ (.A(_3829_),
    .B(_3839_),
    .C(_4004_),
    .X(_4005_));
 sky130_fd_sc_hd__o21ai_1 _4851_ (.A1(_3829_),
    .A2(_3839_),
    .B1(_4004_),
    .Y(_4006_));
 sky130_fd_sc_hd__and2_1 _4852_ (.A(_4005_),
    .B(_4006_),
    .X(_4007_));
 sky130_fd_sc_hd__xnor2_1 _4853_ (.A(_3998_),
    .B(_4007_),
    .Y(_4008_));
 sky130_fd_sc_hd__xnor2_1 _4854_ (.A(_3996_),
    .B(_4008_),
    .Y(_4009_));
 sky130_fd_sc_hd__nand2_1 _4855_ (.A(_3860_),
    .B(_3888_),
    .Y(_4010_));
 sky130_fd_sc_hd__xnor2_1 _4856_ (.A(_4009_),
    .B(_4010_),
    .Y(_4011_));
 sky130_fd_sc_hd__and2_1 _4857_ (.A(_3929_),
    .B(_3931_),
    .X(_4012_));
 sky130_fd_sc_hd__and2b_1 _4858_ (.A_N(_3886_),
    .B(_3873_),
    .X(_4013_));
 sky130_fd_sc_hd__a21o_1 _4859_ (.A1(_3856_),
    .A2(_3885_),
    .B1(_4013_),
    .X(_4014_));
 sky130_fd_sc_hd__or4_2 _4860_ (.A(_1352_),
    .B(_1374_),
    .C(_1396_),
    .D(_1407_),
    .X(_4015_));
 sky130_fd_sc_hd__nor2_8 _4861_ (.A(\posit_add.in2[14] ),
    .B(_4015_),
    .Y(_4016_));
 sky130_fd_sc_hd__buf_4 _4862_ (.A(_4016_),
    .X(_4017_));
 sky130_fd_sc_hd__nor2_2 _4863_ (.A(_4017_),
    .B(_3725_),
    .Y(_4018_));
 sky130_fd_sc_hd__xor2_1 _4864_ (.A(_4018_),
    .B(_3927_),
    .X(_4019_));
 sky130_fd_sc_hd__or3_1 _4865_ (.A(_3701_),
    .B(_3930_),
    .C(_4019_),
    .X(_4020_));
 sky130_fd_sc_hd__o21ai_1 _4866_ (.A1(_3701_),
    .A2(_3930_),
    .B1(_4019_),
    .Y(_4021_));
 sky130_fd_sc_hd__nand2_1 _4867_ (.A(_4020_),
    .B(_4021_),
    .Y(_4022_));
 sky130_fd_sc_hd__xnor2_1 _4868_ (.A(_4022_),
    .B(_3928_),
    .Y(_4023_));
 sky130_fd_sc_hd__nor2_1 _4869_ (.A(_3719_),
    .B(_3795_),
    .Y(_4024_));
 sky130_fd_sc_hd__xnor2_1 _4870_ (.A(_4023_),
    .B(_4024_),
    .Y(_4025_));
 sky130_fd_sc_hd__xor2_1 _4871_ (.A(_4014_),
    .B(_4025_),
    .X(_4026_));
 sky130_fd_sc_hd__xnor2_1 _4872_ (.A(_4012_),
    .B(_4026_),
    .Y(_4027_));
 sky130_fd_sc_hd__xnor2_2 _4873_ (.A(_4011_),
    .B(_4027_),
    .Y(_4028_));
 sky130_fd_sc_hd__and2b_1 _4874_ (.A_N(_3890_),
    .B(_3913_),
    .X(_4029_));
 sky130_fd_sc_hd__o21bai_2 _4875_ (.A1(_3914_),
    .A2(_3936_),
    .B1_N(_4029_),
    .Y(_4030_));
 sky130_fd_sc_hd__xnor2_2 _4876_ (.A(_4028_),
    .B(_4030_),
    .Y(_4031_));
 sky130_fd_sc_hd__o21ba_1 _4877_ (.A1(_3935_),
    .A2(_3728_),
    .B1_N(_3933_),
    .X(_4032_));
 sky130_fd_sc_hd__xnor2_2 _4878_ (.A(_4031_),
    .B(_4032_),
    .Y(_4033_));
 sky130_fd_sc_hd__or2b_1 _4879_ (.A(_3937_),
    .B_N(_3953_),
    .X(_4034_));
 sky130_fd_sc_hd__a21boi_1 _4880_ (.A1(_3807_),
    .A2(_3954_),
    .B1_N(_4034_),
    .Y(_4035_));
 sky130_fd_sc_hd__xor2_1 _4881_ (.A(_4033_),
    .B(_4035_),
    .X(_4036_));
 sky130_fd_sc_hd__clkbuf_4 _4882_ (.A(_3750_),
    .X(_4037_));
 sky130_fd_sc_hd__nor2_1 _4883_ (.A(_2540_),
    .B(_4037_),
    .Y(_4038_));
 sky130_fd_sc_hd__xor2_1 _4884_ (.A(_4036_),
    .B(_4038_),
    .X(_4039_));
 sky130_fd_sc_hd__or2b_1 _4885_ (.A(_3985_),
    .B_N(_4039_),
    .X(_4040_));
 sky130_fd_sc_hd__or2b_1 _4886_ (.A(_4039_),
    .B_N(_3985_),
    .X(_4041_));
 sky130_fd_sc_hd__nand2_1 _4887_ (.A(_4040_),
    .B(_4041_),
    .Y(_4042_));
 sky130_fd_sc_hd__a31oi_2 _4888_ (.A1(_1990_),
    .A2(_2320_),
    .A3(_2419_),
    .B1(_2496_),
    .Y(_4043_));
 sky130_fd_sc_hd__nor2_1 _4889_ (.A(_3729_),
    .B(_4043_),
    .Y(_4044_));
 sky130_fd_sc_hd__buf_4 _4890_ (.A(_4044_),
    .X(_4045_));
 sky130_fd_sc_hd__nand2_1 _4891_ (.A(_4045_),
    .B(_3986_),
    .Y(_4046_));
 sky130_fd_sc_hd__xnor2_1 _4892_ (.A(_3984_),
    .B(_4046_),
    .Y(_4047_));
 sky130_fd_sc_hd__xor2_2 _4893_ (.A(_3963_),
    .B(_3981_),
    .X(_4048_));
 sky130_fd_sc_hd__xnor2_1 _4894_ (.A(_3965_),
    .B(_3978_),
    .Y(_4049_));
 sky130_fd_sc_hd__a32o_1 _4895_ (.A1(_3722_),
    .A2(_3754_),
    .A3(_3878_),
    .B1(_3868_),
    .B2(_3776_),
    .X(_4050_));
 sky130_fd_sc_hd__o31a_1 _4896_ (.A1(_3792_),
    .A2(_3755_),
    .A3(_3959_),
    .B1(_4050_),
    .X(_4051_));
 sky130_fd_sc_hd__and4_1 _4897_ (.A(_3892_),
    .B(_3832_),
    .C(_3943_),
    .D(_3868_),
    .X(_4052_));
 sky130_fd_sc_hd__xor2_1 _4898_ (.A(_4051_),
    .B(_4052_),
    .X(_4053_));
 sky130_fd_sc_hd__and3_1 _4899_ (.A(_3878_),
    .B(_3907_),
    .C(_3789_),
    .X(_4054_));
 sky130_fd_sc_hd__nand2_1 _4900_ (.A(_4051_),
    .B(_4052_),
    .Y(_4055_));
 sky130_fd_sc_hd__a21bo_1 _4901_ (.A1(_4053_),
    .A2(_4054_),
    .B1_N(_4055_),
    .X(_4056_));
 sky130_fd_sc_hd__xnor2_1 _4902_ (.A(_3968_),
    .B(_3975_),
    .Y(_4057_));
 sky130_fd_sc_hd__xnor2_1 _4903_ (.A(_3971_),
    .B(_3973_),
    .Y(_4058_));
 sky130_fd_sc_hd__xnor2_1 _4904_ (.A(_4053_),
    .B(_4054_),
    .Y(_4059_));
 sky130_fd_sc_hd__or2_1 _4905_ (.A(_4058_),
    .B(_4059_),
    .X(_4060_));
 sky130_fd_sc_hd__xor2_1 _4906_ (.A(_4057_),
    .B(_4060_),
    .X(_4061_));
 sky130_fd_sc_hd__nor2_1 _4907_ (.A(_4057_),
    .B(_4060_),
    .Y(_4062_));
 sky130_fd_sc_hd__a21o_1 _4908_ (.A1(_4056_),
    .A2(_4061_),
    .B1(_4062_),
    .X(_4063_));
 sky130_fd_sc_hd__and2b_1 _4909_ (.A_N(_4049_),
    .B(_4063_),
    .X(_4064_));
 sky130_fd_sc_hd__xnor2_1 _4910_ (.A(_4048_),
    .B(_4064_),
    .Y(_4065_));
 sky130_fd_sc_hd__or3_1 _4911_ (.A(_2540_),
    .B(_3817_),
    .C(_4065_),
    .X(_4066_));
 sky130_fd_sc_hd__a21bo_1 _4912_ (.A1(_4048_),
    .A2(_4064_),
    .B1_N(_4066_),
    .X(_4067_));
 sky130_fd_sc_hd__xnor2_1 _4913_ (.A(_4047_),
    .B(_4067_),
    .Y(_4068_));
 sky130_fd_sc_hd__o21ai_1 _4914_ (.A1(_2540_),
    .A2(_3817_),
    .B1(_4065_),
    .Y(_4069_));
 sky130_fd_sc_hd__nand2_1 _4915_ (.A(_4066_),
    .B(_4069_),
    .Y(_4070_));
 sky130_fd_sc_hd__xor2_1 _4916_ (.A(_4049_),
    .B(_4063_),
    .X(_4071_));
 sky130_fd_sc_hd__xnor2_1 _4917_ (.A(_4056_),
    .B(_4061_),
    .Y(_4072_));
 sky130_fd_sc_hd__nor2_1 _4918_ (.A(_3739_),
    .B(_3702_),
    .Y(_4073_));
 sky130_fd_sc_hd__and3_1 _4919_ (.A(_3892_),
    .B(_3883_),
    .C(_4073_),
    .X(_4074_));
 sky130_fd_sc_hd__o32a_1 _4920_ (.A1(_3772_),
    .A2(_3771_),
    .A3(_3882_),
    .B1(_3702_),
    .B2(_3792_),
    .X(_4075_));
 sky130_fd_sc_hd__a31oi_2 _4921_ (.A1(_3878_),
    .A2(_3907_),
    .A3(_3789_),
    .B1(_4075_),
    .Y(_4076_));
 sky130_fd_sc_hd__xnor2_1 _4922_ (.A(_4074_),
    .B(_4076_),
    .Y(_4077_));
 sky130_fd_sc_hd__or3_1 _4923_ (.A(_3793_),
    .B(_3725_),
    .C(_3959_),
    .X(_4078_));
 sky130_fd_sc_hd__nand2_1 _4924_ (.A(_4074_),
    .B(_4076_),
    .Y(_4079_));
 sky130_fd_sc_hd__o21a_1 _4925_ (.A1(_4077_),
    .A2(_4078_),
    .B1(_4079_),
    .X(_4080_));
 sky130_fd_sc_hd__xor2_1 _4926_ (.A(_4058_),
    .B(_4059_),
    .X(_4081_));
 sky130_fd_sc_hd__o22a_1 _4927_ (.A1(_3845_),
    .A2(_3817_),
    .B1(_3930_),
    .B2(_3828_),
    .X(_4082_));
 sky130_fd_sc_hd__or2_1 _4928_ (.A(_4052_),
    .B(_4082_),
    .X(_4083_));
 sky130_fd_sc_hd__xor2_1 _4929_ (.A(_4077_),
    .B(_4078_),
    .X(_4084_));
 sky130_fd_sc_hd__and2b_1 _4930_ (.A_N(_4083_),
    .B(_4084_),
    .X(_4085_));
 sky130_fd_sc_hd__xnor2_1 _4931_ (.A(_4081_),
    .B(_4085_),
    .Y(_4086_));
 sky130_fd_sc_hd__nand2_1 _4932_ (.A(_4081_),
    .B(_4085_),
    .Y(_4087_));
 sky130_fd_sc_hd__o21a_1 _4933_ (.A1(_4080_),
    .A2(_4086_),
    .B1(_4087_),
    .X(_4088_));
 sky130_fd_sc_hd__buf_4 _4934_ (.A(_3883_),
    .X(_4089_));
 sky130_fd_sc_hd__nand2_1 _4935_ (.A(_4045_),
    .B(_4089_),
    .Y(_4090_));
 sky130_fd_sc_hd__nor2_1 _4936_ (.A(_4072_),
    .B(_4088_),
    .Y(_4091_));
 sky130_fd_sc_hd__xnor2_1 _4937_ (.A(_4071_),
    .B(_4091_),
    .Y(_4092_));
 sky130_fd_sc_hd__or2b_1 _4938_ (.A(_4090_),
    .B_N(_4092_),
    .X(_4093_));
 sky130_fd_sc_hd__o31a_1 _4939_ (.A1(_4071_),
    .A2(_4072_),
    .A3(_4088_),
    .B1(_4093_),
    .X(_4094_));
 sky130_fd_sc_hd__nand2_1 _4940_ (.A(_4070_),
    .B(_4094_),
    .Y(_4095_));
 sky130_fd_sc_hd__xnor2_1 _4941_ (.A(_4090_),
    .B(_4092_),
    .Y(_4096_));
 sky130_fd_sc_hd__nor2_1 _4942_ (.A(_2540_),
    .B(_3930_),
    .Y(_4097_));
 sky130_fd_sc_hd__and2_1 _4943_ (.A(_4072_),
    .B(_4088_),
    .X(_4098_));
 sky130_fd_sc_hd__or2_1 _4944_ (.A(_4091_),
    .B(_4098_),
    .X(_4099_));
 sky130_fd_sc_hd__xnor2_1 _4945_ (.A(_4080_),
    .B(_4086_),
    .Y(_4100_));
 sky130_fd_sc_hd__or4_1 _4946_ (.A(_3828_),
    .B(_3845_),
    .C(_3930_),
    .D(_3726_),
    .X(_4101_));
 sky130_fd_sc_hd__o21ai_1 _4947_ (.A1(_3793_),
    .A2(_3726_),
    .B1(_3959_),
    .Y(_4102_));
 sky130_fd_sc_hd__and2_1 _4948_ (.A(_4078_),
    .B(_4102_),
    .X(_4103_));
 sky130_fd_sc_hd__or2b_1 _4949_ (.A(_4101_),
    .B_N(_4103_),
    .X(_4104_));
 sky130_fd_sc_hd__o22a_1 _4950_ (.A1(_3845_),
    .A2(_3795_),
    .B1(_3702_),
    .B2(_3828_),
    .X(_4105_));
 sky130_fd_sc_hd__nor2_1 _4951_ (.A(_4074_),
    .B(_4105_),
    .Y(_4106_));
 sky130_fd_sc_hd__xnor2_1 _4952_ (.A(_4101_),
    .B(_4103_),
    .Y(_4107_));
 sky130_fd_sc_hd__nand2_1 _4953_ (.A(_4106_),
    .B(_4107_),
    .Y(_4108_));
 sky130_fd_sc_hd__xnor2_1 _4954_ (.A(_4083_),
    .B(_4084_),
    .Y(_4109_));
 sky130_fd_sc_hd__a21boi_1 _4955_ (.A1(_4104_),
    .A2(_4108_),
    .B1_N(_4109_),
    .Y(_4110_));
 sky130_fd_sc_hd__and2b_1 _4956_ (.A_N(_4100_),
    .B(_4110_),
    .X(_4111_));
 sky130_fd_sc_hd__xnor2_1 _4957_ (.A(_4099_),
    .B(_4111_),
    .Y(_4112_));
 sky130_fd_sc_hd__and2b_1 _4958_ (.A_N(_4099_),
    .B(_4111_),
    .X(_4113_));
 sky130_fd_sc_hd__a21oi_1 _4959_ (.A1(_4097_),
    .A2(_4112_),
    .B1(_4113_),
    .Y(_4114_));
 sky130_fd_sc_hd__xnor2_1 _4960_ (.A(_4096_),
    .B(_4114_),
    .Y(_4115_));
 sky130_fd_sc_hd__xnor2_1 _4961_ (.A(_4109_),
    .B(_4108_),
    .Y(_4116_));
 sky130_fd_sc_hd__xnor2_2 _4962_ (.A(_4104_),
    .B(_4116_),
    .Y(_4117_));
 sky130_fd_sc_hd__xnor2_1 _4963_ (.A(_4106_),
    .B(_4107_),
    .Y(_4118_));
 sky130_fd_sc_hd__or2_1 _4964_ (.A(_3771_),
    .B(_3703_),
    .X(_4119_));
 sky130_fd_sc_hd__a22o_1 _4965_ (.A1(_3832_),
    .A2(_3868_),
    .B1(_3804_),
    .B2(_3893_),
    .X(_4120_));
 sky130_fd_sc_hd__nand2_1 _4966_ (.A(_4101_),
    .B(_4120_),
    .Y(_4121_));
 sky130_fd_sc_hd__xor2_1 _4967_ (.A(_4119_),
    .B(_4121_),
    .X(_4122_));
 sky130_fd_sc_hd__or4b_1 _4968_ (.A(_3845_),
    .B(_3726_),
    .C(_4119_),
    .D_N(_4122_),
    .X(_4123_));
 sky130_fd_sc_hd__nor2_1 _4969_ (.A(_4118_),
    .B(_4123_),
    .Y(_4124_));
 sky130_fd_sc_hd__nand2_1 _4970_ (.A(_4117_),
    .B(_4124_),
    .Y(_4125_));
 sky130_fd_sc_hd__buf_4 _4971_ (.A(_3726_),
    .X(_4126_));
 sky130_fd_sc_hd__or3_1 _4972_ (.A(_4119_),
    .B(_4118_),
    .C(_4121_),
    .X(_4127_));
 sky130_fd_sc_hd__inv_2 _4973_ (.A(_4127_),
    .Y(_4128_));
 sky130_fd_sc_hd__or2_1 _4974_ (.A(_4128_),
    .B(_4124_),
    .X(_4129_));
 sky130_fd_sc_hd__xnor2_1 _4975_ (.A(_4117_),
    .B(_4129_),
    .Y(_4130_));
 sky130_fd_sc_hd__or3_1 _4976_ (.A(_2529_),
    .B(_4126_),
    .C(_4130_),
    .X(_4131_));
 sky130_fd_sc_hd__or2_1 _4977_ (.A(_2529_),
    .B(_3703_),
    .X(_4132_));
 sky130_fd_sc_hd__xnor2_1 _4978_ (.A(_4100_),
    .B(_4110_),
    .Y(_4133_));
 sky130_fd_sc_hd__nand2_1 _4979_ (.A(_4117_),
    .B(_4128_),
    .Y(_4134_));
 sky130_fd_sc_hd__xor2_1 _4980_ (.A(_4133_),
    .B(_4134_),
    .X(_4135_));
 sky130_fd_sc_hd__nor2_1 _4981_ (.A(_4132_),
    .B(_4135_),
    .Y(_4136_));
 sky130_fd_sc_hd__and2_1 _4982_ (.A(_4132_),
    .B(_4135_),
    .X(_4137_));
 sky130_fd_sc_hd__or2_1 _4983_ (.A(_4136_),
    .B(_4137_),
    .X(_4138_));
 sky130_fd_sc_hd__a21o_1 _4984_ (.A1(_4125_),
    .A2(_4131_),
    .B1(_4138_),
    .X(_4139_));
 sky130_fd_sc_hd__inv_2 _4985_ (.A(_4139_),
    .Y(_4140_));
 sky130_fd_sc_hd__xnor2_1 _4986_ (.A(_4097_),
    .B(_4112_),
    .Y(_4141_));
 sky130_fd_sc_hd__a31o_1 _4987_ (.A1(_4133_),
    .A2(_4117_),
    .A3(_4128_),
    .B1(_4136_),
    .X(_4142_));
 sky130_fd_sc_hd__xnor2_1 _4988_ (.A(_4141_),
    .B(_4142_),
    .Y(_4143_));
 sky130_fd_sc_hd__and2b_1 _4989_ (.A_N(_4141_),
    .B(_4142_),
    .X(_4144_));
 sky130_fd_sc_hd__a21o_1 _4990_ (.A1(_4140_),
    .A2(_4143_),
    .B1(_4144_),
    .X(_4145_));
 sky130_fd_sc_hd__and2b_1 _4991_ (.A_N(_4114_),
    .B(_4096_),
    .X(_4146_));
 sky130_fd_sc_hd__a21o_1 _4992_ (.A1(_4115_),
    .A2(_4145_),
    .B1(_4146_),
    .X(_4147_));
 sky130_fd_sc_hd__nor2_1 _4993_ (.A(_4070_),
    .B(_4094_),
    .Y(_4148_));
 sky130_fd_sc_hd__a21o_1 _4994_ (.A1(_4095_),
    .A2(_4147_),
    .B1(_4148_),
    .X(_4149_));
 sky130_fd_sc_hd__and2b_1 _4995_ (.A_N(_4047_),
    .B(_4067_),
    .X(_4150_));
 sky130_fd_sc_hd__a21oi_1 _4996_ (.A1(_4068_),
    .A2(_4149_),
    .B1(_4150_),
    .Y(_4151_));
 sky130_fd_sc_hd__xor2_1 _4997_ (.A(_4042_),
    .B(_4151_),
    .X(_4152_));
 sky130_fd_sc_hd__buf_4 _4998_ (.A(_3838_),
    .X(_4153_));
 sky130_fd_sc_hd__a32o_1 _4999_ (.A1(_3929_),
    .A2(_3931_),
    .A3(_4026_),
    .B1(_4025_),
    .B2(_4014_),
    .X(_4154_));
 sky130_fd_sc_hd__nand2_1 _5000_ (.A(_3998_),
    .B(_4007_),
    .Y(_4155_));
 sky130_fd_sc_hd__nor2_1 _5001_ (.A(_3719_),
    .B(_3817_),
    .Y(_4156_));
 sky130_fd_sc_hd__nor2_2 _5002_ (.A(_4016_),
    .B(_3702_),
    .Y(_4157_));
 sky130_fd_sc_hd__nor2_1 _5003_ (.A(_3924_),
    .B(_3930_),
    .Y(_4158_));
 sky130_fd_sc_hd__xor2_1 _5004_ (.A(_4157_),
    .B(_4158_),
    .X(_4159_));
 sky130_fd_sc_hd__or3b_1 _5005_ (.A(_3701_),
    .B(_3795_),
    .C_N(_4159_),
    .X(_4160_));
 sky130_fd_sc_hd__a21o_1 _5006_ (.A1(_3802_),
    .A2(_3883_),
    .B1(_4159_),
    .X(_4161_));
 sky130_fd_sc_hd__and2_1 _5007_ (.A(_4160_),
    .B(_4161_),
    .X(_4162_));
 sky130_fd_sc_hd__o31a_1 _5008_ (.A1(_4017_),
    .A2(_3726_),
    .A3(_3927_),
    .B1(_4020_),
    .X(_4163_));
 sky130_fd_sc_hd__xnor2_1 _5009_ (.A(_4162_),
    .B(_4163_),
    .Y(_4164_));
 sky130_fd_sc_hd__xnor2_1 _5010_ (.A(_4156_),
    .B(_4164_),
    .Y(_4165_));
 sky130_fd_sc_hd__a21oi_1 _5011_ (.A1(_4005_),
    .A2(_4155_),
    .B1(_4165_),
    .Y(_4166_));
 sky130_fd_sc_hd__and3_1 _5012_ (.A(_4005_),
    .B(_4155_),
    .C(_4165_),
    .X(_4167_));
 sky130_fd_sc_hd__or2_1 _5013_ (.A(_4166_),
    .B(_4167_),
    .X(_4168_));
 sky130_fd_sc_hd__o32a_1 _5014_ (.A1(_3800_),
    .A2(_3795_),
    .A3(_4023_),
    .B1(_3928_),
    .B2(_4022_),
    .X(_4169_));
 sky130_fd_sc_hd__xnor2_1 _5015_ (.A(_4168_),
    .B(_4169_),
    .Y(_4170_));
 sky130_fd_sc_hd__or2_1 _5016_ (.A(_3996_),
    .B(_4008_),
    .X(_4171_));
 sky130_fd_sc_hd__nand2_1 _5017_ (.A(_3893_),
    .B(_3854_),
    .Y(_4172_));
 sky130_fd_sc_hd__nand2_1 _5018_ (.A(_3881_),
    .B(_3894_),
    .Y(_4173_));
 sky130_fd_sc_hd__or3_2 _5019_ (.A(\posit_add.in1[14] ),
    .B(_3013_),
    .C(_2584_),
    .X(_4174_));
 sky130_fd_sc_hd__and4_1 _5020_ (.A(_3776_),
    .B(_3878_),
    .C(_3855_),
    .D(_4174_),
    .X(_4175_));
 sky130_fd_sc_hd__o22a_1 _5021_ (.A1(_3793_),
    .A2(_3988_),
    .B1(_3989_),
    .B2(_3771_),
    .X(_4176_));
 sky130_fd_sc_hd__nor2_1 _5022_ (.A(_4175_),
    .B(_4176_),
    .Y(_4177_));
 sky130_fd_sc_hd__xnor2_1 _5023_ (.A(_4173_),
    .B(_4177_),
    .Y(_4178_));
 sky130_fd_sc_hd__xnor2_1 _5024_ (.A(_4172_),
    .B(_4178_),
    .Y(_4179_));
 sky130_fd_sc_hd__a21bo_1 _5025_ (.A1(_4000_),
    .A2(_4001_),
    .B1_N(_3999_),
    .X(_4180_));
 sky130_fd_sc_hd__xnor2_1 _5026_ (.A(_4179_),
    .B(_4180_),
    .Y(_4181_));
 sky130_fd_sc_hd__or2_1 _5027_ (.A(_3827_),
    .B(_3816_),
    .X(_4182_));
 sky130_fd_sc_hd__or3_1 _5028_ (.A(_3828_),
    .B(_3750_),
    .C(_4182_),
    .X(_4183_));
 sky130_fd_sc_hd__o21ai_1 _5029_ (.A1(_3816_),
    .A2(_4037_),
    .B1(_3829_),
    .Y(_4184_));
 sky130_fd_sc_hd__and2_1 _5030_ (.A(_4183_),
    .B(_4184_),
    .X(_4185_));
 sky130_fd_sc_hd__nor2_1 _5031_ (.A(_3987_),
    .B(_3991_),
    .Y(_4186_));
 sky130_fd_sc_hd__nand2_1 _5032_ (.A(_4185_),
    .B(_4186_),
    .Y(_4187_));
 sky130_fd_sc_hd__or2_1 _5033_ (.A(_4185_),
    .B(_4186_),
    .X(_4188_));
 sky130_fd_sc_hd__nand2_1 _5034_ (.A(_4187_),
    .B(_4188_),
    .Y(_4189_));
 sky130_fd_sc_hd__xnor2_1 _5035_ (.A(_4181_),
    .B(_4189_),
    .Y(_4190_));
 sky130_fd_sc_hd__a21oi_1 _5036_ (.A1(_3994_),
    .A2(_4171_),
    .B1(_4190_),
    .Y(_4191_));
 sky130_fd_sc_hd__and3_1 _5037_ (.A(_4190_),
    .B(_3994_),
    .C(_4171_),
    .X(_4192_));
 sky130_fd_sc_hd__nor2_1 _5038_ (.A(_4191_),
    .B(_4192_),
    .Y(_4193_));
 sky130_fd_sc_hd__xnor2_1 _5039_ (.A(_4170_),
    .B(_4193_),
    .Y(_4194_));
 sky130_fd_sc_hd__and3_1 _5040_ (.A(_4009_),
    .B(_3860_),
    .C(_3888_),
    .X(_4195_));
 sky130_fd_sc_hd__and2b_1 _5041_ (.A_N(_4009_),
    .B(_4010_),
    .X(_4196_));
 sky130_fd_sc_hd__o21ba_1 _5042_ (.A1(_4195_),
    .A2(_4027_),
    .B1_N(_4196_),
    .X(_4197_));
 sky130_fd_sc_hd__xnor2_1 _5043_ (.A(_4194_),
    .B(_4197_),
    .Y(_4198_));
 sky130_fd_sc_hd__xnor2_1 _5044_ (.A(_4154_),
    .B(_4198_),
    .Y(_4199_));
 sky130_fd_sc_hd__nor2_1 _5045_ (.A(_4031_),
    .B(_4032_),
    .Y(_4200_));
 sky130_fd_sc_hd__a21oi_1 _5046_ (.A1(_4028_),
    .A2(_4030_),
    .B1(_4200_),
    .Y(_4201_));
 sky130_fd_sc_hd__xor2_1 _5047_ (.A(_4199_),
    .B(_4201_),
    .X(_4202_));
 sky130_fd_sc_hd__and3_1 _5048_ (.A(_4045_),
    .B(_4153_),
    .C(_4202_),
    .X(_4203_));
 sky130_fd_sc_hd__a21oi_1 _5049_ (.A1(_4045_),
    .A2(_4153_),
    .B1(_4202_),
    .Y(_4204_));
 sky130_fd_sc_hd__nor2_1 _5050_ (.A(_4203_),
    .B(_4204_),
    .Y(_4205_));
 sky130_fd_sc_hd__o2bb2a_1 _5051_ (.A1_N(_4036_),
    .A2_N(_4038_),
    .B1(_4033_),
    .B2(_4035_),
    .X(_4206_));
 sky130_fd_sc_hd__xnor2_1 _5052_ (.A(_4205_),
    .B(_4206_),
    .Y(_4207_));
 sky130_fd_sc_hd__o21ai_1 _5053_ (.A1(_4042_),
    .A2(_4151_),
    .B1(_4040_),
    .Y(_4208_));
 sky130_fd_sc_hd__xor2_1 _5054_ (.A(_4207_),
    .B(_4208_),
    .X(_4209_));
 sky130_fd_sc_hd__buf_4 _5055_ (.A(_4017_),
    .X(_4210_));
 sky130_fd_sc_hd__or2_1 _5056_ (.A(_4210_),
    .B(_3615_),
    .X(_4211_));
 sky130_fd_sc_hd__or2_1 _5057_ (.A(_3925_),
    .B(_4037_),
    .X(_4212_));
 sky130_fd_sc_hd__nor2_1 _5058_ (.A(_4210_),
    .B(_3615_),
    .Y(_4213_));
 sky130_fd_sc_hd__xnor2_1 _5059_ (.A(_4213_),
    .B(_4212_),
    .Y(_4214_));
 sky130_fd_sc_hd__and3_1 _5060_ (.A(_3802_),
    .B(_3838_),
    .C(_4214_),
    .X(_4215_));
 sky130_fd_sc_hd__o21ba_1 _5061_ (.A1(_4211_),
    .A2(_4212_),
    .B1_N(_4215_),
    .X(_4216_));
 sky130_fd_sc_hd__buf_6 _5062_ (.A(_3855_),
    .X(_4217_));
 sky130_fd_sc_hd__nand2_1 _5063_ (.A(_3802_),
    .B(_4217_),
    .Y(_4218_));
 sky130_fd_sc_hd__or2_1 _5064_ (.A(_4210_),
    .B(_3840_),
    .X(_4219_));
 sky130_fd_sc_hd__or2_1 _5065_ (.A(_4210_),
    .B(_4037_),
    .X(_4220_));
 sky130_fd_sc_hd__o22a_1 _5066_ (.A1(_3917_),
    .A2(_3922_),
    .B1(_3769_),
    .B2(_1748_),
    .X(_4221_));
 sky130_fd_sc_hd__buf_4 _5067_ (.A(_4221_),
    .X(_4222_));
 sky130_fd_sc_hd__nand2_1 _5068_ (.A(_4222_),
    .B(_3838_),
    .Y(_4223_));
 sky130_fd_sc_hd__nand2_1 _5069_ (.A(_4220_),
    .B(_4223_),
    .Y(_4224_));
 sky130_fd_sc_hd__o21ai_1 _5070_ (.A1(_4219_),
    .A2(_4212_),
    .B1(_4224_),
    .Y(_4225_));
 sky130_fd_sc_hd__xor2_1 _5071_ (.A(_4218_),
    .B(_4225_),
    .X(_4226_));
 sky130_fd_sc_hd__and2b_1 _5072_ (.A_N(_4216_),
    .B(_4226_),
    .X(_4227_));
 sky130_fd_sc_hd__buf_4 _5073_ (.A(_3827_),
    .X(_4228_));
 sky130_fd_sc_hd__nor2_1 _5074_ (.A(_4228_),
    .B(_3800_),
    .Y(_4229_));
 sky130_fd_sc_hd__xnor2_1 _5075_ (.A(_4226_),
    .B(_4216_),
    .Y(_4230_));
 sky130_fd_sc_hd__and2_1 _5076_ (.A(_4229_),
    .B(_4230_),
    .X(_4231_));
 sky130_fd_sc_hd__buf_4 _5077_ (.A(_3989_),
    .X(_4232_));
 sky130_fd_sc_hd__nor2_1 _5078_ (.A(_4228_),
    .B(_3701_),
    .Y(_4233_));
 sky130_fd_sc_hd__nor2_1 _5079_ (.A(_3988_),
    .B(_4223_),
    .Y(_4234_));
 sky130_fd_sc_hd__nor2_1 _5080_ (.A(_4210_),
    .B(_3840_),
    .Y(_4235_));
 sky130_fd_sc_hd__a21oi_1 _5081_ (.A1(_4222_),
    .A2(_3855_),
    .B1(_4235_),
    .Y(_4236_));
 sky130_fd_sc_hd__nor2_1 _5082_ (.A(_4234_),
    .B(_4236_),
    .Y(_4237_));
 sky130_fd_sc_hd__xnor2_1 _5083_ (.A(_4233_),
    .B(_4237_),
    .Y(_4238_));
 sky130_fd_sc_hd__o22a_1 _5084_ (.A1(_4220_),
    .A2(_4223_),
    .B1(_4225_),
    .B2(_4218_),
    .X(_4239_));
 sky130_fd_sc_hd__or2_1 _5085_ (.A(_4238_),
    .B(_4239_),
    .X(_4240_));
 sky130_fd_sc_hd__nand2_1 _5086_ (.A(_4238_),
    .B(_4239_),
    .Y(_4241_));
 sky130_fd_sc_hd__nand2_1 _5087_ (.A(_4240_),
    .B(_4241_),
    .Y(_4242_));
 sky130_fd_sc_hd__or3_1 _5088_ (.A(_3800_),
    .B(_4232_),
    .C(_4242_),
    .X(_4243_));
 sky130_fd_sc_hd__o21ai_1 _5089_ (.A1(_3800_),
    .A2(_4232_),
    .B1(_4242_),
    .Y(_4244_));
 sky130_fd_sc_hd__and2_1 _5090_ (.A(_4243_),
    .B(_4244_),
    .X(_4245_));
 sky130_fd_sc_hd__o21a_1 _5091_ (.A1(_4227_),
    .A2(_4231_),
    .B1(_4245_),
    .X(_4246_));
 sky130_fd_sc_hd__nand2_1 _5092_ (.A(_4240_),
    .B(_4243_),
    .Y(_4247_));
 sky130_fd_sc_hd__and2_1 _5093_ (.A(_4233_),
    .B(_4237_),
    .X(_4248_));
 sky130_fd_sc_hd__nor2_1 _5094_ (.A(_3701_),
    .B(_4232_),
    .Y(_4249_));
 sky130_fd_sc_hd__buf_4 _5095_ (.A(_4210_),
    .X(_4250_));
 sky130_fd_sc_hd__or2_2 _5096_ (.A(_4250_),
    .B(_3988_),
    .X(_4251_));
 sky130_fd_sc_hd__nor2_1 _5097_ (.A(_4228_),
    .B(_3925_),
    .Y(_4252_));
 sky130_fd_sc_hd__xnor2_1 _5098_ (.A(_4251_),
    .B(_4252_),
    .Y(_4253_));
 sky130_fd_sc_hd__nand2_1 _5099_ (.A(_4249_),
    .B(_4253_),
    .Y(_4254_));
 sky130_fd_sc_hd__or2_1 _5100_ (.A(_4249_),
    .B(_4253_),
    .X(_4255_));
 sky130_fd_sc_hd__and2_1 _5101_ (.A(_4254_),
    .B(_4255_),
    .X(_4256_));
 sky130_fd_sc_hd__o21ai_2 _5102_ (.A1(_4234_),
    .A2(_4248_),
    .B1(_4256_),
    .Y(_0075_));
 sky130_fd_sc_hd__or3_1 _5103_ (.A(_4234_),
    .B(_4248_),
    .C(_4256_),
    .X(_0076_));
 sky130_fd_sc_hd__nand2_1 _5104_ (.A(_0075_),
    .B(_0076_),
    .Y(_0077_));
 sky130_fd_sc_hd__xnor2_1 _5105_ (.A(_4247_),
    .B(_0077_),
    .Y(_0078_));
 sky130_fd_sc_hd__nand2_1 _5106_ (.A(_4246_),
    .B(_0078_),
    .Y(_0079_));
 sky130_fd_sc_hd__buf_4 _5107_ (.A(_4228_),
    .X(_0080_));
 sky130_fd_sc_hd__o31a_1 _5108_ (.A1(_0080_),
    .A2(_3925_),
    .A3(_4251_),
    .B1(_4254_),
    .X(_0081_));
 sky130_fd_sc_hd__buf_4 _5109_ (.A(_4232_),
    .X(_0082_));
 sky130_fd_sc_hd__or2_1 _5110_ (.A(_4228_),
    .B(_4250_),
    .X(_0083_));
 sky130_fd_sc_hd__o21a_1 _5111_ (.A1(_3925_),
    .A2(_0082_),
    .B1(_0083_),
    .X(_0084_));
 sky130_fd_sc_hd__or2_1 _5112_ (.A(_4252_),
    .B(_0084_),
    .X(_0085_));
 sky130_fd_sc_hd__xnor2_1 _5113_ (.A(_0081_),
    .B(_0085_),
    .Y(_0086_));
 sky130_fd_sc_hd__a21o_1 _5114_ (.A1(_4240_),
    .A2(_4243_),
    .B1(_0077_),
    .X(_0087_));
 sky130_fd_sc_hd__nand2_1 _5115_ (.A(_0075_),
    .B(_0087_),
    .Y(_0088_));
 sky130_fd_sc_hd__xor2_1 _5116_ (.A(_0086_),
    .B(_0088_),
    .X(_0089_));
 sky130_fd_sc_hd__nor2_1 _5117_ (.A(_0079_),
    .B(_0089_),
    .Y(_0090_));
 sky130_fd_sc_hd__or2_1 _5118_ (.A(_0087_),
    .B(_0086_),
    .X(_0091_));
 sky130_fd_sc_hd__or2_4 _5119_ (.A(_4210_),
    .B(_3989_),
    .X(_0092_));
 sky130_fd_sc_hd__o21bai_1 _5120_ (.A1(_4254_),
    .A2(_0084_),
    .B1_N(_4252_),
    .Y(_0093_));
 sky130_fd_sc_hd__o21a_1 _5121_ (.A1(_0092_),
    .A2(_0093_),
    .B1(_0075_),
    .X(_0094_));
 sky130_fd_sc_hd__nor2_1 _5122_ (.A(_0091_),
    .B(_0094_),
    .Y(_0095_));
 sky130_fd_sc_hd__nor3_1 _5123_ (.A(_0092_),
    .B(_0075_),
    .C(_0093_),
    .Y(_0096_));
 sky130_fd_sc_hd__o21a_1 _5124_ (.A1(_0094_),
    .A2(_0096_),
    .B1(_0091_),
    .X(_0097_));
 sky130_fd_sc_hd__nor2_1 _5125_ (.A(_0095_),
    .B(_0097_),
    .Y(_0098_));
 sky130_fd_sc_hd__xor2_1 _5126_ (.A(_0090_),
    .B(_0098_),
    .X(_0099_));
 sky130_fd_sc_hd__or2_1 _5127_ (.A(_4246_),
    .B(_0078_),
    .X(_0100_));
 sky130_fd_sc_hd__and2_1 _5128_ (.A(_0079_),
    .B(_0100_),
    .X(_0101_));
 sky130_fd_sc_hd__xnor2_1 _5129_ (.A(_4229_),
    .B(_4230_),
    .Y(_0102_));
 sky130_fd_sc_hd__a21oi_1 _5130_ (.A1(_3802_),
    .A2(_3838_),
    .B1(_4214_),
    .Y(_0103_));
 sky130_fd_sc_hd__nor2_1 _5131_ (.A(_4215_),
    .B(_0103_),
    .Y(_0104_));
 sky130_fd_sc_hd__or2_2 _5132_ (.A(_4017_),
    .B(_3755_),
    .X(_0105_));
 sky130_fd_sc_hd__or3_1 _5133_ (.A(_3925_),
    .B(_3615_),
    .C(_0105_),
    .X(_0106_));
 sky130_fd_sc_hd__o21ai_1 _5134_ (.A1(_3925_),
    .A2(_3615_),
    .B1(_0105_),
    .Y(_0107_));
 sky130_fd_sc_hd__nand2_1 _5135_ (.A(_0106_),
    .B(_0107_),
    .Y(_0108_));
 sky130_fd_sc_hd__or3_1 _5136_ (.A(_3701_),
    .B(_3750_),
    .C(_0108_),
    .X(_0109_));
 sky130_fd_sc_hd__nand2_1 _5137_ (.A(_0106_),
    .B(_0109_),
    .Y(_0110_));
 sky130_fd_sc_hd__a2bb2o_1 _5138_ (.A1_N(_3716_),
    .A2_N(_3711_),
    .B1(_3710_),
    .B2(_3690_),
    .X(_0111_));
 sky130_fd_sc_hd__clkbuf_4 _5139_ (.A(_0111_),
    .X(_0112_));
 sky130_fd_sc_hd__buf_4 _5140_ (.A(_0112_),
    .X(_0113_));
 sky130_fd_sc_hd__nand2_1 _5141_ (.A(_0113_),
    .B(_4217_),
    .Y(_0114_));
 sky130_fd_sc_hd__xor2_1 _5142_ (.A(_0104_),
    .B(_0110_),
    .X(_0115_));
 sky130_fd_sc_hd__clkinv_2 _5143_ (.A(_0115_),
    .Y(_0116_));
 sky130_fd_sc_hd__o2bb2a_1 _5144_ (.A1_N(_0104_),
    .A2_N(_0110_),
    .B1(_0114_),
    .B2(_0116_),
    .X(_0117_));
 sky130_fd_sc_hd__nor2_1 _5145_ (.A(_0102_),
    .B(_0117_),
    .Y(_0118_));
 sky130_fd_sc_hd__and2_1 _5146_ (.A(_0102_),
    .B(_0117_),
    .X(_0119_));
 sky130_fd_sc_hd__or2_1 _5147_ (.A(_0118_),
    .B(_0119_),
    .X(_0120_));
 sky130_fd_sc_hd__buf_4 _5148_ (.A(_4174_),
    .X(_0121_));
 sky130_fd_sc_hd__and3_1 _5149_ (.A(_3881_),
    .B(_0121_),
    .C(_4182_),
    .X(_0122_));
 sky130_fd_sc_hd__or2b_1 _5150_ (.A(_0120_),
    .B_N(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__or2_1 _5151_ (.A(_3827_),
    .B(_3763_),
    .X(_0124_));
 sky130_fd_sc_hd__or3_1 _5152_ (.A(_3816_),
    .B(_3989_),
    .C(_0124_),
    .X(_0125_));
 sky130_fd_sc_hd__nor3_1 _5153_ (.A(_4227_),
    .B(_4231_),
    .C(_4245_),
    .Y(_0126_));
 sky130_fd_sc_hd__or2_1 _5154_ (.A(_4246_),
    .B(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__a21oi_1 _5155_ (.A1(_0123_),
    .A2(_0125_),
    .B1(_0127_),
    .Y(_0128_));
 sky130_fd_sc_hd__and3_1 _5156_ (.A(_0127_),
    .B(_0123_),
    .C(_0125_),
    .X(_0129_));
 sky130_fd_sc_hd__nor2_1 _5157_ (.A(_0128_),
    .B(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__a21o_1 _5158_ (.A1(_0118_),
    .A2(_0130_),
    .B1(_0128_),
    .X(_0131_));
 sky130_fd_sc_hd__nand2_1 _5159_ (.A(_0101_),
    .B(_0131_),
    .Y(_0132_));
 sky130_fd_sc_hd__xnor2_1 _5160_ (.A(_0101_),
    .B(_0131_),
    .Y(_0133_));
 sky130_fd_sc_hd__xnor2_1 _5161_ (.A(_0118_),
    .B(_0130_),
    .Y(_0134_));
 sky130_fd_sc_hd__xor2_1 _5162_ (.A(_0120_),
    .B(_0122_),
    .X(_0135_));
 sky130_fd_sc_hd__o21ai_1 _5163_ (.A1(_3816_),
    .A2(_4232_),
    .B1(_0124_),
    .Y(_0136_));
 sky130_fd_sc_hd__and4_1 _5164_ (.A(_3881_),
    .B(_3776_),
    .C(_3838_),
    .D(_0121_),
    .X(_0137_));
 sky130_fd_sc_hd__nand2_1 _5165_ (.A(_3855_),
    .B(_0137_),
    .Y(_0138_));
 sky130_fd_sc_hd__a21o_1 _5166_ (.A1(_3881_),
    .A2(_3855_),
    .B1(_0137_),
    .X(_0139_));
 sky130_fd_sc_hd__nand2_1 _5167_ (.A(_0138_),
    .B(_0139_),
    .Y(_0140_));
 sky130_fd_sc_hd__o2bb2a_1 _5168_ (.A1_N(_0125_),
    .A2_N(_0136_),
    .B1(_0140_),
    .B2(_4182_),
    .X(_0141_));
 sky130_fd_sc_hd__xnor2_1 _5169_ (.A(_0114_),
    .B(_0115_),
    .Y(_0142_));
 sky130_fd_sc_hd__xnor2_1 _5170_ (.A(_0138_),
    .B(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__o21ai_1 _5171_ (.A1(_3701_),
    .A2(_4037_),
    .B1(_0108_),
    .Y(_0144_));
 sky130_fd_sc_hd__nand2_1 _5172_ (.A(_0109_),
    .B(_0144_),
    .Y(_0145_));
 sky130_fd_sc_hd__nand2_1 _5173_ (.A(_3802_),
    .B(_3986_),
    .Y(_0146_));
 sky130_fd_sc_hd__buf_4 _5174_ (.A(_3943_),
    .X(_0147_));
 sky130_fd_sc_hd__nor2_1 _5175_ (.A(_4017_),
    .B(_3795_),
    .Y(_0148_));
 sky130_fd_sc_hd__a21oi_1 _5176_ (.A1(_4222_),
    .A2(_0147_),
    .B1(_0148_),
    .Y(_0149_));
 sky130_fd_sc_hd__or3_1 _5177_ (.A(_3925_),
    .B(_0105_),
    .C(_3795_),
    .X(_0150_));
 sky130_fd_sc_hd__o21a_1 _5178_ (.A1(_0146_),
    .A2(_0149_),
    .B1(_0150_),
    .X(_0151_));
 sky130_fd_sc_hd__xnor2_1 _5179_ (.A(_0145_),
    .B(_0151_),
    .Y(_0152_));
 sky130_fd_sc_hd__and3b_1 _5180_ (.A_N(_0152_),
    .B(_3838_),
    .C(_0113_),
    .X(_0153_));
 sky130_fd_sc_hd__o21ba_1 _5181_ (.A1(_0145_),
    .A2(_0151_),
    .B1_N(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__xnor2_1 _5182_ (.A(_0143_),
    .B(_0154_),
    .Y(_0155_));
 sky130_fd_sc_hd__or2b_1 _5183_ (.A(_0141_),
    .B_N(_0155_),
    .X(_0156_));
 sky130_fd_sc_hd__or2b_1 _5184_ (.A(_0138_),
    .B_N(_0142_),
    .X(_0157_));
 sky130_fd_sc_hd__or2b_1 _5185_ (.A(_0154_),
    .B_N(_0143_),
    .X(_0158_));
 sky130_fd_sc_hd__and2_1 _5186_ (.A(_0157_),
    .B(_0158_),
    .X(_0159_));
 sky130_fd_sc_hd__xnor2_1 _5187_ (.A(_0135_),
    .B(_0156_),
    .Y(_0160_));
 sky130_fd_sc_hd__or2_1 _5188_ (.A(_0159_),
    .B(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__o21ai_1 _5189_ (.A1(_0135_),
    .A2(_0156_),
    .B1(_0161_),
    .Y(_0162_));
 sky130_fd_sc_hd__or2b_1 _5190_ (.A(_0134_),
    .B_N(_0162_),
    .X(_0163_));
 sky130_fd_sc_hd__xor2_1 _5191_ (.A(_0134_),
    .B(_0162_),
    .X(_0164_));
 sky130_fd_sc_hd__nand2_1 _5192_ (.A(_3901_),
    .B(_3838_),
    .Y(_0165_));
 sky130_fd_sc_hd__nand2_1 _5193_ (.A(_3893_),
    .B(_0121_),
    .Y(_0166_));
 sky130_fd_sc_hd__or2_1 _5194_ (.A(_0165_),
    .B(_0166_),
    .X(_0167_));
 sky130_fd_sc_hd__o22a_1 _5195_ (.A1(_3763_),
    .A2(_3840_),
    .B1(_3989_),
    .B2(_3793_),
    .X(_0168_));
 sky130_fd_sc_hd__or4_2 _5196_ (.A(_0124_),
    .B(_0137_),
    .C(_0168_),
    .D(_3875_),
    .X(_0169_));
 sky130_fd_sc_hd__o22ai_1 _5197_ (.A1(_0137_),
    .A2(_0168_),
    .B1(_3875_),
    .B2(_0124_),
    .Y(_0170_));
 sky130_fd_sc_hd__nand2_1 _5198_ (.A(_0169_),
    .B(_0170_),
    .Y(_0171_));
 sky130_fd_sc_hd__o21a_1 _5199_ (.A1(_3816_),
    .A2(_3988_),
    .B1(_0167_),
    .X(_0172_));
 sky130_fd_sc_hd__o22a_1 _5200_ (.A1(_3988_),
    .A2(_0167_),
    .B1(_0171_),
    .B2(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__xor2_1 _5201_ (.A(_4182_),
    .B(_0140_),
    .X(_0174_));
 sky130_fd_sc_hd__and2b_1 _5202_ (.A_N(_0173_),
    .B(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__o21a_1 _5203_ (.A1(_3800_),
    .A2(_3840_),
    .B1(_0152_),
    .X(_0176_));
 sky130_fd_sc_hd__nor2_1 _5204_ (.A(_0153_),
    .B(_0176_),
    .Y(_0177_));
 sky130_fd_sc_hd__xnor2_1 _5205_ (.A(_0169_),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__nor2_1 _5206_ (.A(_3800_),
    .B(_4037_),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _5207_ (.A(_0150_),
    .Y(_0180_));
 sky130_fd_sc_hd__nor2_1 _5208_ (.A(_0180_),
    .B(_0149_),
    .Y(_0181_));
 sky130_fd_sc_hd__xnor2_1 _5209_ (.A(_0146_),
    .B(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__nor2_1 _5210_ (.A(_3701_),
    .B(_3817_),
    .Y(_0183_));
 sky130_fd_sc_hd__nor2_2 _5211_ (.A(_4017_),
    .B(_3930_),
    .Y(_0184_));
 sky130_fd_sc_hd__and3_1 _5212_ (.A(_4222_),
    .B(_3883_),
    .C(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__a21oi_1 _5213_ (.A1(_4222_),
    .A2(_3883_),
    .B1(_0184_),
    .Y(_0186_));
 sky130_fd_sc_hd__nor2_1 _5214_ (.A(_0185_),
    .B(_0186_),
    .Y(_0187_));
 sky130_fd_sc_hd__a21oi_1 _5215_ (.A1(_0183_),
    .A2(_0187_),
    .B1(_0185_),
    .Y(_0188_));
 sky130_fd_sc_hd__xnor2_1 _5216_ (.A(_0182_),
    .B(_0188_),
    .Y(_0189_));
 sky130_fd_sc_hd__or2b_1 _5217_ (.A(_0188_),
    .B_N(_0182_),
    .X(_0190_));
 sky130_fd_sc_hd__a21bo_1 _5218_ (.A1(_0179_),
    .A2(_0189_),
    .B1_N(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__xnor2_1 _5219_ (.A(_0178_),
    .B(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__and2b_1 _5220_ (.A_N(_0174_),
    .B(_0173_),
    .X(_0193_));
 sky130_fd_sc_hd__or2_1 _5221_ (.A(_0175_),
    .B(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__nor2_1 _5222_ (.A(_0192_),
    .B(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__xnor2_1 _5223_ (.A(_0155_),
    .B(_0141_),
    .Y(_0196_));
 sky130_fd_sc_hd__o21a_1 _5224_ (.A1(_0175_),
    .A2(_0195_),
    .B1(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__nor3_1 _5225_ (.A(_0196_),
    .B(_0175_),
    .C(_0195_),
    .Y(_0198_));
 sky130_fd_sc_hd__or2_1 _5226_ (.A(_0197_),
    .B(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__or3_1 _5227_ (.A(_0153_),
    .B(_0169_),
    .C(_0176_),
    .X(_0200_));
 sky130_fd_sc_hd__a21bo_1 _5228_ (.A1(_0178_),
    .A2(_0191_),
    .B1_N(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__and2b_1 _5229_ (.A_N(_0199_),
    .B(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__nand2_1 _5230_ (.A(_0159_),
    .B(_0160_),
    .Y(_0203_));
 sky130_fd_sc_hd__and2_1 _5231_ (.A(_0161_),
    .B(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__o21ai_1 _5232_ (.A1(_0197_),
    .A2(_0202_),
    .B1(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__nor2_1 _5233_ (.A(_0164_),
    .B(_0205_),
    .Y(_0206_));
 sky130_fd_sc_hd__and2_1 _5234_ (.A(_0164_),
    .B(_0205_),
    .X(_0207_));
 sky130_fd_sc_hd__or2_1 _5235_ (.A(_0206_),
    .B(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__inv_2 _5236_ (.A(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__xor2_1 _5237_ (.A(_0165_),
    .B(_0166_),
    .X(_0210_));
 sky130_fd_sc_hd__or4b_1 _5238_ (.A(_3828_),
    .B(_4037_),
    .C(_4182_),
    .D_N(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__and3_1 _5239_ (.A(_3881_),
    .B(_3986_),
    .C(_4177_),
    .X(_0212_));
 sky130_fd_sc_hd__o22a_1 _5240_ (.A1(_3827_),
    .A2(_3793_),
    .B1(_3750_),
    .B2(_3763_),
    .X(_0213_));
 sky130_fd_sc_hd__o21ba_1 _5241_ (.A1(_0124_),
    .A2(_3875_),
    .B1_N(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__o21ai_1 _5242_ (.A1(_4175_),
    .A2(_0212_),
    .B1(_0214_),
    .Y(_0215_));
 sky130_fd_sc_hd__or3_1 _5243_ (.A(_0214_),
    .B(_4175_),
    .C(_0212_),
    .X(_0216_));
 sky130_fd_sc_hd__and2_1 _5244_ (.A(_0215_),
    .B(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__inv_4 _5245_ (.A(_4228_),
    .Y(_0218_));
 sky130_fd_sc_hd__a31o_1 _5246_ (.A1(_0218_),
    .A2(_3901_),
    .A3(_3844_),
    .B1(_0210_),
    .X(_0219_));
 sky130_fd_sc_hd__nand2_1 _5247_ (.A(_0211_),
    .B(_0219_),
    .Y(_0220_));
 sky130_fd_sc_hd__inv_2 _5248_ (.A(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__nand2_1 _5249_ (.A(_0217_),
    .B(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__o21ba_1 _5250_ (.A1(_3988_),
    .A2(_0167_),
    .B1_N(_0172_),
    .X(_0223_));
 sky130_fd_sc_hd__xor2_1 _5251_ (.A(_0171_),
    .B(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__a21o_1 _5252_ (.A1(_0211_),
    .A2(_0222_),
    .B1(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__xnor2_1 _5253_ (.A(_0179_),
    .B(_0189_),
    .Y(_0226_));
 sky130_fd_sc_hd__nor2_1 _5254_ (.A(_0215_),
    .B(_0226_),
    .Y(_0227_));
 sky130_fd_sc_hd__and2_1 _5255_ (.A(_0215_),
    .B(_0226_),
    .X(_0228_));
 sky130_fd_sc_hd__nor2_1 _5256_ (.A(_0227_),
    .B(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__xnor2_1 _5257_ (.A(_0183_),
    .B(_0187_),
    .Y(_0230_));
 sky130_fd_sc_hd__a21bo_1 _5258_ (.A1(_4157_),
    .A2(_4158_),
    .B1_N(_4160_),
    .X(_0231_));
 sky130_fd_sc_hd__xor2_1 _5259_ (.A(_0230_),
    .B(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__or2b_1 _5260_ (.A(_0230_),
    .B_N(_0231_),
    .X(_0233_));
 sky130_fd_sc_hd__o31ai_2 _5261_ (.A1(_3800_),
    .A2(_3615_),
    .A3(_0232_),
    .B1(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__xor2_1 _5262_ (.A(_0229_),
    .B(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__nand3_1 _5263_ (.A(_0224_),
    .B(_0211_),
    .C(_0222_),
    .Y(_0236_));
 sky130_fd_sc_hd__and2_1 _5264_ (.A(_0225_),
    .B(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__nand2_1 _5265_ (.A(_0235_),
    .B(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__nand2_1 _5266_ (.A(_0192_),
    .B(_0194_),
    .Y(_0239_));
 sky130_fd_sc_hd__or2b_1 _5267_ (.A(_0195_),
    .B_N(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__a21oi_1 _5268_ (.A1(_0225_),
    .A2(_0238_),
    .B1(_0240_),
    .Y(_0241_));
 sky130_fd_sc_hd__and3_1 _5269_ (.A(_0240_),
    .B(_0225_),
    .C(_0238_),
    .X(_0242_));
 sky130_fd_sc_hd__or2_1 _5270_ (.A(_0241_),
    .B(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__a21o_1 _5271_ (.A1(_0229_),
    .A2(_0234_),
    .B1(_0227_),
    .X(_0244_));
 sky130_fd_sc_hd__and2b_1 _5272_ (.A_N(_0243_),
    .B(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__xnor2_1 _5273_ (.A(_0201_),
    .B(_0199_),
    .Y(_0246_));
 sky130_fd_sc_hd__o21ai_2 _5274_ (.A1(_0241_),
    .A2(_0245_),
    .B1(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__or3_1 _5275_ (.A(_0204_),
    .B(_0197_),
    .C(_0202_),
    .X(_0248_));
 sky130_fd_sc_hd__and2_1 _5276_ (.A(_0205_),
    .B(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__xor2_1 _5277_ (.A(_0247_),
    .B(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__or2_1 _5278_ (.A(_0235_),
    .B(_0237_),
    .X(_0251_));
 sky130_fd_sc_hd__nand2_1 _5279_ (.A(_0238_),
    .B(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__or2_1 _5280_ (.A(_4181_),
    .B(_4189_),
    .X(_0253_));
 sky130_fd_sc_hd__xnor2_1 _5281_ (.A(_0217_),
    .B(_0221_),
    .Y(_0254_));
 sky130_fd_sc_hd__a21o_1 _5282_ (.A1(_4187_),
    .A2(_0253_),
    .B1(_0254_),
    .X(_0255_));
 sky130_fd_sc_hd__and3_1 _5283_ (.A(_3893_),
    .B(_3854_),
    .C(_4178_),
    .X(_0256_));
 sky130_fd_sc_hd__a21o_1 _5284_ (.A1(_4179_),
    .A2(_4180_),
    .B1(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__nor2_1 _5285_ (.A(_3800_),
    .B(_3615_),
    .Y(_0258_));
 sky130_fd_sc_hd__xnor2_1 _5286_ (.A(_0258_),
    .B(_0232_),
    .Y(_0259_));
 sky130_fd_sc_hd__xnor2_1 _5287_ (.A(_0257_),
    .B(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hd__and2b_1 _5288_ (.A_N(_4163_),
    .B(_4162_),
    .X(_0261_));
 sky130_fd_sc_hd__a21oi_1 _5289_ (.A1(_4156_),
    .A2(_4164_),
    .B1(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__or2_1 _5290_ (.A(_0260_),
    .B(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__nand2_1 _5291_ (.A(_0260_),
    .B(_0262_),
    .Y(_0264_));
 sky130_fd_sc_hd__nand2_1 _5292_ (.A(_0263_),
    .B(_0264_),
    .Y(_0265_));
 sky130_fd_sc_hd__nand3_1 _5293_ (.A(_0254_),
    .B(_4187_),
    .C(_0253_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand2_1 _5294_ (.A(_0255_),
    .B(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__or2_1 _5295_ (.A(_0265_),
    .B(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__and2_1 _5296_ (.A(_0255_),
    .B(_0268_),
    .X(_0269_));
 sky130_fd_sc_hd__xnor2_1 _5297_ (.A(_0252_),
    .B(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__a21bo_1 _5298_ (.A1(_0257_),
    .A2(_0259_),
    .B1_N(_0263_),
    .X(_0271_));
 sky130_fd_sc_hd__and2b_1 _5299_ (.A_N(_0270_),
    .B(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__o21ba_1 _5300_ (.A1(_0252_),
    .A2(_0269_),
    .B1_N(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__xnor2_1 _5301_ (.A(_0244_),
    .B(_0243_),
    .Y(_0274_));
 sky130_fd_sc_hd__or2b_1 _5302_ (.A(_0273_),
    .B_N(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__xnor2_1 _5303_ (.A(_0274_),
    .B(_0273_),
    .Y(_0276_));
 sky130_fd_sc_hd__or3b_1 _5304_ (.A(_2540_),
    .B(_4232_),
    .C_N(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__or3_1 _5305_ (.A(_0246_),
    .B(_0241_),
    .C(_0245_),
    .X(_0278_));
 sky130_fd_sc_hd__nand2_1 _5306_ (.A(_0247_),
    .B(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__a21oi_1 _5307_ (.A1(_0275_),
    .A2(_0277_),
    .B1(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__and3_1 _5308_ (.A(_0279_),
    .B(_0275_),
    .C(_0277_),
    .X(_0281_));
 sky130_fd_sc_hd__nor2_1 _5309_ (.A(_0280_),
    .B(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__a21o_1 _5310_ (.A1(_4045_),
    .A2(_0121_),
    .B1(_0276_),
    .X(_0283_));
 sky130_fd_sc_hd__nand2_1 _5311_ (.A(_0277_),
    .B(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__or2_1 _5312_ (.A(_4228_),
    .B(_2540_),
    .X(_0285_));
 sky130_fd_sc_hd__xor2_1 _5313_ (.A(_0271_),
    .B(_0270_),
    .X(_0286_));
 sky130_fd_sc_hd__and2b_1 _5314_ (.A_N(_4170_),
    .B(_4193_),
    .X(_0287_));
 sky130_fd_sc_hd__nor2_1 _5315_ (.A(_4191_),
    .B(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__nand2_1 _5316_ (.A(_0265_),
    .B(_0267_),
    .Y(_0289_));
 sky130_fd_sc_hd__and2_1 _5317_ (.A(_0268_),
    .B(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__or2b_1 _5318_ (.A(_0288_),
    .B_N(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__o21ba_1 _5319_ (.A1(_4168_),
    .A2(_4169_),
    .B1_N(_4166_),
    .X(_0292_));
 sky130_fd_sc_hd__xnor2_1 _5320_ (.A(_0290_),
    .B(_0288_),
    .Y(_0293_));
 sky130_fd_sc_hd__or2b_1 _5321_ (.A(_0292_),
    .B_N(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__and2_1 _5322_ (.A(_0291_),
    .B(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__xnor2_1 _5323_ (.A(_0286_),
    .B(_0295_),
    .Y(_0296_));
 sky130_fd_sc_hd__or2_1 _5324_ (.A(_0286_),
    .B(_0295_),
    .X(_0297_));
 sky130_fd_sc_hd__o21ai_1 _5325_ (.A1(_0285_),
    .A2(_0296_),
    .B1(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__or2b_1 _5326_ (.A(_0284_),
    .B_N(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__or2b_1 _5327_ (.A(_0298_),
    .B_N(_0284_),
    .X(_0300_));
 sky130_fd_sc_hd__nand2_1 _5328_ (.A(_0299_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__xnor2_1 _5329_ (.A(_0285_),
    .B(_0296_),
    .Y(_0302_));
 sky130_fd_sc_hd__clkbuf_4 _5330_ (.A(_3988_),
    .X(_0303_));
 sky130_fd_sc_hd__xnor2_1 _5331_ (.A(_0292_),
    .B(_0293_),
    .Y(_0304_));
 sky130_fd_sc_hd__o21a_1 _5332_ (.A1(_4191_),
    .A2(_4192_),
    .B1(_4170_),
    .X(_0305_));
 sky130_fd_sc_hd__nand2_1 _5333_ (.A(_4154_),
    .B(_4198_),
    .Y(_0306_));
 sky130_fd_sc_hd__o31a_1 _5334_ (.A1(_0287_),
    .A2(_0305_),
    .A3(_4197_),
    .B1(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__xor2_1 _5335_ (.A(_0304_),
    .B(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__or2b_1 _5336_ (.A(_0307_),
    .B_N(_0304_),
    .X(_0309_));
 sky130_fd_sc_hd__o31a_1 _5337_ (.A1(_2540_),
    .A2(_0303_),
    .A3(_0308_),
    .B1(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__nor2_1 _5338_ (.A(_0302_),
    .B(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__and2_1 _5339_ (.A(_0302_),
    .B(_0310_),
    .X(_0312_));
 sky130_fd_sc_hd__nor2_1 _5340_ (.A(_0311_),
    .B(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__o21ba_1 _5341_ (.A1(_4199_),
    .A2(_4201_),
    .B1_N(_4203_),
    .X(_0314_));
 sky130_fd_sc_hd__nor2_1 _5342_ (.A(_2540_),
    .B(_3988_),
    .Y(_0315_));
 sky130_fd_sc_hd__xnor2_1 _5343_ (.A(_0315_),
    .B(_0308_),
    .Y(_0316_));
 sky130_fd_sc_hd__or2b_1 _5344_ (.A(_0314_),
    .B_N(_0316_),
    .X(_0317_));
 sky130_fd_sc_hd__or2b_1 _5345_ (.A(_0316_),
    .B_N(_0314_),
    .X(_0318_));
 sky130_fd_sc_hd__nand2_1 _5346_ (.A(_0317_),
    .B(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__and2b_1 _5347_ (.A_N(_4206_),
    .B(_4205_),
    .X(_0320_));
 sky130_fd_sc_hd__a21oi_1 _5348_ (.A1(_4207_),
    .A2(_4208_),
    .B1(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__o21ai_1 _5349_ (.A1(_0319_),
    .A2(_0321_),
    .B1(_0317_),
    .Y(_0322_));
 sky130_fd_sc_hd__a21oi_1 _5350_ (.A1(_0313_),
    .A2(_0322_),
    .B1(_0311_),
    .Y(_0323_));
 sky130_fd_sc_hd__o21ai_1 _5351_ (.A1(_0301_),
    .A2(_0323_),
    .B1(_0299_),
    .Y(_0324_));
 sky130_fd_sc_hd__a21oi_1 _5352_ (.A1(_0282_),
    .A2(_0324_),
    .B1(_0280_),
    .Y(_0325_));
 sky130_fd_sc_hd__and2b_1 _5353_ (.A_N(_0247_),
    .B(_0249_),
    .X(_0326_));
 sky130_fd_sc_hd__o21bai_1 _5354_ (.A1(_0250_),
    .A2(_0325_),
    .B1_N(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__a21oi_1 _5355_ (.A1(_0209_),
    .A2(_0327_),
    .B1(_0206_),
    .Y(_0328_));
 sky130_fd_sc_hd__xor2_1 _5356_ (.A(_0133_),
    .B(_0163_),
    .X(_0329_));
 sky130_fd_sc_hd__and2b_1 _5357_ (.A_N(_0328_),
    .B(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__o21bai_1 _5358_ (.A1(_0133_),
    .A2(_0163_),
    .B1_N(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__a21oi_1 _5359_ (.A1(_0079_),
    .A2(_0132_),
    .B1(_0089_),
    .Y(_0332_));
 sky130_fd_sc_hd__a31oi_1 _5360_ (.A1(_0079_),
    .A2(_0089_),
    .A3(_0132_),
    .B1(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__a2bb2o_1 _5361_ (.A1_N(_0089_),
    .A2_N(_0132_),
    .B1(_0331_),
    .B2(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__or3_1 _5362_ (.A(_0093_),
    .B(_0096_),
    .C(_0095_),
    .X(_0335_));
 sky130_fd_sc_hd__a21o_1 _5363_ (.A1(_0090_),
    .A2(_0098_),
    .B1(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__a21o_2 _5364_ (.A1(_0099_),
    .A2(_0334_),
    .B1(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__clkbuf_4 _5365_ (.A(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _5366_ (.A0(_4152_),
    .A1(_4209_),
    .S(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__xor2_1 _5367_ (.A(_0319_),
    .B(_0321_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _5368_ (.A0(_4209_),
    .A1(_0340_),
    .S(_0338_),
    .X(_0341_));
 sky130_fd_sc_hd__xnor2_1 _5369_ (.A(_1781_),
    .B(_2452_),
    .Y(_0342_));
 sky130_fd_sc_hd__a211o_1 _5370_ (.A1(_3068_),
    .A2(_3296_),
    .B1(_3328_),
    .C1(_3035_),
    .X(_0343_));
 sky130_fd_sc_hd__nand2_1 _5371_ (.A(_3328_),
    .B(_3318_),
    .Y(_0344_));
 sky130_fd_sc_hd__nand2_1 _5372_ (.A(_0343_),
    .B(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__nor2_1 _5373_ (.A(_0342_),
    .B(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__inv_2 _5374_ (.A(_1781_),
    .Y(_0347_));
 sky130_fd_sc_hd__xnor2_2 _5375_ (.A(_0347_),
    .B(_2452_),
    .Y(_0348_));
 sky130_fd_sc_hd__and2_1 _5376_ (.A(_0343_),
    .B(_0344_),
    .X(_0349_));
 sky130_fd_sc_hd__nor2_2 _5377_ (.A(_0348_),
    .B(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__or2_2 _5378_ (.A(_0346_),
    .B(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__a211o_1 _5379_ (.A1(_3079_),
    .A2(_3296_),
    .B1(_3101_),
    .C1(_3046_),
    .X(_0352_));
 sky130_fd_sc_hd__o21a_1 _5380_ (.A1(_2727_),
    .A2(_3530_),
    .B1(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _5381_ (.A0(_3068_),
    .A1(_0353_),
    .S(_3446_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _5382_ (.A0(_3850_),
    .A1(_0354_),
    .S(_3156_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_4 _5383_ (.A0(_3754_),
    .A1(_0355_),
    .S(_3721_),
    .X(_0356_));
 sky130_fd_sc_hd__nand3_1 _5384_ (.A(_3736_),
    .B(_3659_),
    .C(_3671_),
    .Y(_0357_));
 sky130_fd_sc_hd__or2_1 _5385_ (.A(_1484_),
    .B(_2452_),
    .X(_0358_));
 sky130_fd_sc_hd__o21ai_1 _5386_ (.A1(_1583_),
    .A2(_3635_),
    .B1(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__nor2_1 _5387_ (.A(_3830_),
    .B(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__a211o_1 _5388_ (.A1(_1451_),
    .A2(_3830_),
    .B1(_0360_),
    .C1(_3736_),
    .X(_0361_));
 sky130_fd_sc_hd__nor2_1 _5389_ (.A(_1748_),
    .B(_2507_),
    .Y(_0362_));
 sky130_fd_sc_hd__a31o_2 _5390_ (.A1(_0357_),
    .A2(_1748_),
    .A3(_0361_),
    .B1(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__or2b_1 _5391_ (.A(_0356_),
    .B_N(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__a21oi_4 _5392_ (.A1(_3690_),
    .A2(_3716_),
    .B1(_3774_),
    .Y(_0365_));
 sky130_fd_sc_hd__and3_1 _5393_ (.A(_1748_),
    .B(_3706_),
    .C(_3708_),
    .X(_0366_));
 sky130_fd_sc_hd__a211o_1 _5394_ (.A1(_1484_),
    .A2(_3830_),
    .B1(_3729_),
    .C1(_3736_),
    .X(_0367_));
 sky130_fd_sc_hd__a21oi_1 _5395_ (.A1(_2309_),
    .A2(_3920_),
    .B1(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__a221oi_4 _5396_ (.A1(_3729_),
    .A2(_0365_),
    .B1(_0366_),
    .B2(_3736_),
    .C1(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__clkinv_2 _5397_ (.A(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__a211o_1 _5398_ (.A1(_2760_),
    .A2(_3307_),
    .B1(_3822_),
    .C1(_3477_),
    .X(_0371_));
 sky130_fd_sc_hd__o21a_1 _5399_ (.A1(_3101_),
    .A2(_3446_),
    .B1(_3145_),
    .X(_0372_));
 sky130_fd_sc_hd__a32oi_4 _5400_ (.A1(_3520_),
    .A2(_3833_),
    .A3(_3834_),
    .B1(_0371_),
    .B2(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__mux2_4 _5401_ (.A0(_3882_),
    .A1(_0373_),
    .S(_3721_),
    .X(_0374_));
 sky130_fd_sc_hd__xnor2_4 _5402_ (.A(_0370_),
    .B(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__a21oi_2 _5403_ (.A1(_3741_),
    .A2(_3743_),
    .B1(_3156_),
    .Y(_0376_));
 sky130_fd_sc_hd__o211a_1 _5404_ (.A1(_2727_),
    .A2(_3530_),
    .B1(_0352_),
    .C1(_3488_),
    .X(_0377_));
 sky130_fd_sc_hd__o211a_1 _5405_ (.A1(_3819_),
    .A2(_3530_),
    .B1(_3848_),
    .C1(_3446_),
    .X(_0378_));
 sky130_fd_sc_hd__o31ai_4 _5406_ (.A1(_3520_),
    .A2(_0377_),
    .A3(_0378_),
    .B1(_3721_),
    .Y(_0379_));
 sky130_fd_sc_hd__nand4_2 _5407_ (.A(_3594_),
    .B(_3156_),
    .C(_3746_),
    .D(_3748_),
    .Y(_0380_));
 sky130_fd_sc_hd__a211o_1 _5408_ (.A1(_1605_),
    .A2(_3635_),
    .B1(_3651_),
    .C1(_3830_),
    .X(_0381_));
 sky130_fd_sc_hd__o21a_1 _5409_ (.A1(_2309_),
    .A2(_0359_),
    .B1(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__a21o_1 _5410_ (.A1(_3757_),
    .A2(_3758_),
    .B1(_3690_),
    .X(_0383_));
 sky130_fd_sc_hd__o21ai_1 _5411_ (.A1(_3736_),
    .A2(_0382_),
    .B1(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__mux2_2 _5412_ (.A0(_0384_),
    .A1(_3733_),
    .S(_3729_),
    .X(_0385_));
 sky130_fd_sc_hd__o211a_1 _5413_ (.A1(_0376_),
    .A2(_0379_),
    .B1(_0380_),
    .C1(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__inv_2 _5414_ (.A(_0385_),
    .Y(_0387_));
 sky130_fd_sc_hd__o21ai_4 _5415_ (.A1(_0376_),
    .A2(_0379_),
    .B1(_0380_),
    .Y(_0388_));
 sky130_fd_sc_hd__and2_1 _5416_ (.A(_0387_),
    .B(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__or2_2 _5417_ (.A(_0386_),
    .B(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__inv_2 _5418_ (.A(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__a21o_1 _5419_ (.A1(_0391_),
    .A2(_0337_),
    .B1(_0389_),
    .X(_0392_));
 sky130_fd_sc_hd__nor2_1 _5420_ (.A(_0369_),
    .B(_0374_),
    .Y(_0393_));
 sky130_fd_sc_hd__a21o_1 _5421_ (.A1(_0375_),
    .A2(_0392_),
    .B1(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__and2b_1 _5422_ (.A_N(_0363_),
    .B(_0356_),
    .X(_0395_));
 sky130_fd_sc_hd__a21o_1 _5423_ (.A1(_0364_),
    .A2(_0394_),
    .B1(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__xnor2_2 _5424_ (.A(_0351_),
    .B(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__inv_2 _5425_ (.A(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__nand2_2 _5426_ (.A(_3328_),
    .B(_1781_),
    .Y(_0399_));
 sky130_fd_sc_hd__nor2_1 _5427_ (.A(_0347_),
    .B(_4210_),
    .Y(_0400_));
 sky130_fd_sc_hd__a21oi_1 _5428_ (.A1(_3328_),
    .A2(_0121_),
    .B1(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__inv_2 _5429_ (.A(_1946_),
    .Y(_0402_));
 sky130_fd_sc_hd__a21o_1 _5430_ (.A1(_0347_),
    .A2(_0402_),
    .B1(_1748_),
    .X(_0403_));
 sky130_fd_sc_hd__a31o_1 _5431_ (.A1(_3690_),
    .A2(_3830_),
    .A3(_3635_),
    .B1(_0347_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _5432_ (.A0(_3729_),
    .A1(_0403_),
    .S(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__o21ai_1 _5433_ (.A1(_3328_),
    .A2(_2826_),
    .B1(_3772_),
    .Y(_0406_));
 sky130_fd_sc_hd__a21o_1 _5434_ (.A1(_3424_),
    .A2(_3530_),
    .B1(_2980_),
    .X(_0407_));
 sky130_fd_sc_hd__inv_2 _5435_ (.A(_0343_),
    .Y(_0408_));
 sky130_fd_sc_hd__nand2_1 _5436_ (.A(_3424_),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__xnor2_2 _5437_ (.A(_3167_),
    .B(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__a21o_1 _5438_ (.A1(_0407_),
    .A2(_0410_),
    .B1(_2980_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _5439_ (.A0(_3772_),
    .A1(_0406_),
    .S(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__nor2_1 _5440_ (.A(_0405_),
    .B(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__and2_1 _5441_ (.A(_0405_),
    .B(_0412_),
    .X(_0414_));
 sky130_fd_sc_hd__or2_1 _5442_ (.A(_0413_),
    .B(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__inv_2 _5443_ (.A(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__xnor2_1 _5444_ (.A(_0407_),
    .B(_0410_),
    .Y(_0417_));
 sky130_fd_sc_hd__nand2_1 _5445_ (.A(_3830_),
    .B(_3635_),
    .Y(_0418_));
 sky130_fd_sc_hd__or2_1 _5446_ (.A(_1781_),
    .B(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__xnor2_1 _5447_ (.A(_3690_),
    .B(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__nand2_1 _5448_ (.A(_1781_),
    .B(_0418_),
    .Y(_0421_));
 sky130_fd_sc_hd__mux2_1 _5449_ (.A0(_3736_),
    .A1(_0420_),
    .S(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__nor2_1 _5450_ (.A(_0417_),
    .B(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__and2_1 _5451_ (.A(_0417_),
    .B(_0422_),
    .X(_0424_));
 sky130_fd_sc_hd__nor2_2 _5452_ (.A(_0423_),
    .B(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__xnor2_1 _5453_ (.A(_3830_),
    .B(_0348_),
    .Y(_0426_));
 sky130_fd_sc_hd__o21a_1 _5454_ (.A1(_3488_),
    .A2(_0408_),
    .B1(_0409_),
    .X(_0427_));
 sky130_fd_sc_hd__clkinv_2 _5455_ (.A(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__mux2_1 _5456_ (.A0(_3488_),
    .A1(_0428_),
    .S(_0344_),
    .X(_0429_));
 sky130_fd_sc_hd__or2_1 _5457_ (.A(_0426_),
    .B(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__nand2_1 _5458_ (.A(_0426_),
    .B(_0429_),
    .Y(_0431_));
 sky130_fd_sc_hd__and2_1 _5459_ (.A(_0430_),
    .B(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_4 _5460_ (.A(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__nand2_1 _5461_ (.A(_0348_),
    .B(_0349_),
    .Y(_0434_));
 sky130_fd_sc_hd__a21oi_4 _5462_ (.A1(_0434_),
    .A2(_0396_),
    .B1(_0350_),
    .Y(_0435_));
 sky130_fd_sc_hd__and2b_1 _5463_ (.A_N(_0426_),
    .B(_0429_),
    .X(_0436_));
 sky130_fd_sc_hd__o21bai_2 _5464_ (.A1(_0433_),
    .A2(_0435_),
    .B1_N(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__a21o_1 _5465_ (.A1(_0425_),
    .A2(_0437_),
    .B1(_0423_),
    .X(_0438_));
 sky130_fd_sc_hd__a21o_1 _5466_ (.A1(_0416_),
    .A2(_0438_),
    .B1(_0413_),
    .X(_0439_));
 sky130_fd_sc_hd__o32a_4 _5467_ (.A1(_4250_),
    .A2(_0082_),
    .A3(_0399_),
    .B1(_0401_),
    .B2(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__xnor2_1 _5468_ (.A(_0398_),
    .B(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__xor2_4 _5469_ (.A(_0356_),
    .B(_0363_),
    .X(_0442_));
 sky130_fd_sc_hd__xnor2_2 _5470_ (.A(_0442_),
    .B(_0394_),
    .Y(_0443_));
 sky130_fd_sc_hd__xor2_2 _5471_ (.A(_0375_),
    .B(_0392_),
    .X(_0444_));
 sky130_fd_sc_hd__xnor2_2 _5472_ (.A(_0390_),
    .B(_0337_),
    .Y(_0445_));
 sky130_fd_sc_hd__or4_2 _5473_ (.A(_0397_),
    .B(_0443_),
    .C(_0444_),
    .D(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__inv_2 _5474_ (.A(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__inv_2 _5475_ (.A(_0425_),
    .Y(_0448_));
 sky130_fd_sc_hd__xnor2_2 _5476_ (.A(_0448_),
    .B(_0437_),
    .Y(_0449_));
 sky130_fd_sc_hd__xor2_4 _5477_ (.A(_0433_),
    .B(_0435_),
    .X(_0450_));
 sky130_fd_sc_hd__clkinv_2 _5478_ (.A(_0440_),
    .Y(_0451_));
 sky130_fd_sc_hd__o21a_1 _5479_ (.A1(_0446_),
    .A2(_0450_),
    .B1(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__xnor2_1 _5480_ (.A(_0449_),
    .B(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__or2_1 _5481_ (.A(_0447_),
    .B(_0440_),
    .X(_0454_));
 sky130_fd_sc_hd__xnor2_2 _5482_ (.A(_0450_),
    .B(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__or4b_1 _5483_ (.A(_0447_),
    .B(_0453_),
    .C(_0441_),
    .D_N(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__xnor2_2 _5484_ (.A(_0416_),
    .B(_0438_),
    .Y(_0457_));
 sky130_fd_sc_hd__nor3_2 _5485_ (.A(_0446_),
    .B(_0450_),
    .C(_0449_),
    .Y(_0458_));
 sky130_fd_sc_hd__or2_1 _5486_ (.A(_0440_),
    .B(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__xnor2_1 _5487_ (.A(_0457_),
    .B(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__nor2_1 _5488_ (.A(_0092_),
    .B(_0399_),
    .Y(_0461_));
 sky130_fd_sc_hd__or2_1 _5489_ (.A(_0461_),
    .B(_0401_),
    .X(_0462_));
 sky130_fd_sc_hd__a21bo_1 _5490_ (.A1(_0457_),
    .A2(_0458_),
    .B1_N(_0461_),
    .X(_0463_));
 sky130_fd_sc_hd__nand3_1 _5491_ (.A(_0462_),
    .B(_0439_),
    .C(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__nor2_1 _5492_ (.A(_0461_),
    .B(_0401_),
    .Y(_0465_));
 sky130_fd_sc_hd__a2111o_1 _5493_ (.A1(_0457_),
    .A2(_0458_),
    .B1(_0465_),
    .C1(_0439_),
    .D1(_0440_),
    .X(_0466_));
 sky130_fd_sc_hd__nand2_2 _5494_ (.A(_0464_),
    .B(_0466_),
    .Y(_0467_));
 sky130_fd_sc_hd__o21bai_2 _5495_ (.A1(_0456_),
    .A2(_0460_),
    .B1_N(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__or2_2 _5496_ (.A(_0441_),
    .B(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_4 _5497_ (.A(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _5498_ (.A0(_0339_),
    .A1(_0341_),
    .S(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__or2b_1 _5499_ (.A(_4148_),
    .B_N(_4095_),
    .X(_0472_));
 sky130_fd_sc_hd__xnor2_1 _5500_ (.A(_0472_),
    .B(_4147_),
    .Y(_0473_));
 sky130_fd_sc_hd__xor2_1 _5501_ (.A(_4068_),
    .B(_4149_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _5502_ (.A0(_0473_),
    .A1(_0474_),
    .S(_0338_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _5503_ (.A0(_0474_),
    .A1(_4152_),
    .S(_0337_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _5504_ (.A0(_0475_),
    .A1(_0476_),
    .S(_0469_),
    .X(_0477_));
 sky130_fd_sc_hd__nor2_1 _5505_ (.A(_0447_),
    .B(_0441_),
    .Y(_0478_));
 sky130_fd_sc_hd__xor2_2 _5506_ (.A(_0478_),
    .B(_0455_),
    .X(_0479_));
 sky130_fd_sc_hd__nor2_4 _5507_ (.A(_0468_),
    .B(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__mux2_1 _5508_ (.A0(_0471_),
    .A1(_0477_),
    .S(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__xor2_1 _5509_ (.A(_0301_),
    .B(_0323_),
    .X(_0482_));
 sky130_fd_sc_hd__xor2_1 _5510_ (.A(_0282_),
    .B(_0324_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _5511_ (.A0(_0482_),
    .A1(_0483_),
    .S(_0338_),
    .X(_0484_));
 sky130_fd_sc_hd__xor2_1 _5512_ (.A(_0250_),
    .B(_0325_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _5513_ (.A0(_0483_),
    .A1(_0485_),
    .S(_0338_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _5514_ (.A0(_0484_),
    .A1(_0486_),
    .S(_0470_),
    .X(_0487_));
 sky130_fd_sc_hd__xor2_1 _5515_ (.A(_0313_),
    .B(_0322_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _5516_ (.A0(_0340_),
    .A1(_0488_),
    .S(_0337_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _5517_ (.A0(_0488_),
    .A1(_0482_),
    .S(_0337_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _5518_ (.A0(_0489_),
    .A1(_0490_),
    .S(_0469_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _5519_ (.A0(_0487_),
    .A1(_0491_),
    .S(_0480_),
    .X(_0492_));
 sky130_fd_sc_hd__a21bo_1 _5520_ (.A1(_0478_),
    .A2(_0455_),
    .B1_N(_0453_),
    .X(_0493_));
 sky130_fd_sc_hd__a21o_2 _5521_ (.A1(_0456_),
    .A2(_0493_),
    .B1(_0468_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _5522_ (.A0(_0481_),
    .A1(_0492_),
    .S(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__clkinv_2 _5523_ (.A(_0495_),
    .Y(_0496_));
 sky130_fd_sc_hd__and2b_1 _5524_ (.A_N(_0329_),
    .B(_0328_),
    .X(_0497_));
 sky130_fd_sc_hd__nor2_1 _5525_ (.A(_0330_),
    .B(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__xor2_1 _5526_ (.A(_0331_),
    .B(_0333_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _5527_ (.A0(_0498_),
    .A1(_0499_),
    .S(_0338_),
    .X(_0500_));
 sky130_fd_sc_hd__or2_1 _5528_ (.A(_0099_),
    .B(_0334_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _5529_ (.A0(_0499_),
    .A1(_0501_),
    .S(_0336_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _5530_ (.A0(_0500_),
    .A1(_0502_),
    .S(_0470_),
    .X(_0503_));
 sky130_fd_sc_hd__xnor2_1 _5531_ (.A(_0208_),
    .B(_0327_),
    .Y(_0504_));
 sky130_fd_sc_hd__mux2_1 _5532_ (.A0(_0485_),
    .A1(_0504_),
    .S(_0338_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _5533_ (.A0(_0504_),
    .A1(_0498_),
    .S(_0337_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _5534_ (.A0(_0505_),
    .A1(_0506_),
    .S(_0469_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _5535_ (.A0(_0503_),
    .A1(_0507_),
    .S(_0480_),
    .X(_0508_));
 sky130_fd_sc_hd__inv_2 _5536_ (.A(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__buf_2 _5537_ (.A(_0470_),
    .X(_0510_));
 sky130_fd_sc_hd__nand2_1 _5538_ (.A(_0440_),
    .B(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__o21ai_1 _5539_ (.A1(_0443_),
    .A2(_0510_),
    .B1(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__or2b_1 _5540_ (.A(_0444_),
    .B_N(_0510_),
    .X(_0513_));
 sky130_fd_sc_hd__o21ai_1 _5541_ (.A1(_0445_),
    .A2(_0510_),
    .B1(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__clkbuf_4 _5542_ (.A(_0480_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _5543_ (.A0(_0512_),
    .A1(_0514_),
    .S(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _5544_ (.A0(_0509_),
    .A1(_0516_),
    .S(_0494_),
    .X(_0517_));
 sky130_fd_sc_hd__nand2_1 _5545_ (.A(_0456_),
    .B(_0460_),
    .Y(_0518_));
 sky130_fd_sc_hd__or2_2 _5546_ (.A(_0518_),
    .B(_0467_),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _5547_ (.A0(_0496_),
    .A1(_0517_),
    .S(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__nor2_4 _5548_ (.A(_0518_),
    .B(_0467_),
    .Y(_0521_));
 sky130_fd_sc_hd__mux2_1 _5549_ (.A0(_0502_),
    .A1(_0445_),
    .S(_0510_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _5550_ (.A0(_0506_),
    .A1(_0500_),
    .S(_0510_),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _5551_ (.A0(_0522_),
    .A1(_0523_),
    .S(_0515_),
    .X(_0524_));
 sky130_fd_sc_hd__o31ai_1 _5552_ (.A1(_0397_),
    .A2(_0440_),
    .A3(_0468_),
    .B1(_0511_),
    .Y(_0525_));
 sky130_fd_sc_hd__mux2_1 _5553_ (.A0(_0444_),
    .A1(_0443_),
    .S(_0510_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _5554_ (.A0(_0525_),
    .A1(_0526_),
    .S(_0515_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _5555_ (.A0(_0524_),
    .A1(_0527_),
    .S(_0494_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _5556_ (.A0(_0486_),
    .A1(_0505_),
    .S(_0470_),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _5557_ (.A0(_0490_),
    .A1(_0484_),
    .S(_0470_),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _5558_ (.A0(_0529_),
    .A1(_0530_),
    .S(_0480_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _5559_ (.A0(_0341_),
    .A1(_0489_),
    .S(_0470_),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_1 _5560_ (.A0(_0476_),
    .A1(_0339_),
    .S(_0470_),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _5561_ (.A0(_0532_),
    .A1(_0533_),
    .S(_0480_),
    .X(_0534_));
 sky130_fd_sc_hd__inv_2 _5562_ (.A(_0494_),
    .Y(_0535_));
 sky130_fd_sc_hd__mux2_1 _5563_ (.A0(_0531_),
    .A1(_0534_),
    .S(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__or2_1 _5564_ (.A(_0519_),
    .B(_0536_),
    .X(_0537_));
 sky130_fd_sc_hd__o21ai_1 _5565_ (.A1(_0521_),
    .A2(_0528_),
    .B1(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hd__xor2_1 _5566_ (.A(_4115_),
    .B(_4145_),
    .X(_0539_));
 sky130_fd_sc_hd__mux2_1 _5567_ (.A0(_0539_),
    .A1(_0473_),
    .S(_0338_),
    .X(_0540_));
 sky130_fd_sc_hd__mux2_1 _5568_ (.A0(_0540_),
    .A1(_0475_),
    .S(_0470_),
    .X(_0541_));
 sky130_fd_sc_hd__xnor2_1 _5569_ (.A(_4139_),
    .B(_4143_),
    .Y(_0542_));
 sky130_fd_sc_hd__mux2_1 _5570_ (.A0(_0542_),
    .A1(_0539_),
    .S(_0338_),
    .X(_0543_));
 sky130_fd_sc_hd__mux2_1 _5571_ (.A0(_0543_),
    .A1(_0540_),
    .S(_0470_),
    .X(_0544_));
 sky130_fd_sc_hd__o21ba_1 _5572_ (.A1(_0541_),
    .A2(_0544_),
    .B1_N(_0515_),
    .X(_0545_));
 sky130_fd_sc_hd__and3_1 _5573_ (.A(_4138_),
    .B(_4125_),
    .C(_4131_),
    .X(_0546_));
 sky130_fd_sc_hd__nor2_1 _5574_ (.A(_4140_),
    .B(_0546_),
    .Y(_0547_));
 sky130_fd_sc_hd__clkbuf_4 _5575_ (.A(_4126_),
    .X(_0548_));
 sky130_fd_sc_hd__o21ai_1 _5576_ (.A1(_2540_),
    .A2(_0548_),
    .B1(_4130_),
    .Y(_0549_));
 sky130_fd_sc_hd__o211a_1 _5577_ (.A1(_4119_),
    .A2(_4121_),
    .B1(_4123_),
    .C1(_4118_),
    .X(_0550_));
 sky130_fd_sc_hd__nor2_1 _5578_ (.A(_3845_),
    .B(_0548_),
    .Y(_0551_));
 sky130_fd_sc_hd__a2111oi_1 _5579_ (.A1(_3878_),
    .A2(_3804_),
    .B1(_4073_),
    .C1(_0551_),
    .D1(_4122_),
    .Y(_0552_));
 sky130_fd_sc_hd__o21ai_1 _5580_ (.A1(_4129_),
    .A2(_0550_),
    .B1(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__a21o_1 _5581_ (.A1(_4131_),
    .A2(_0549_),
    .B1(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__a211o_1 _5582_ (.A1(_0338_),
    .A2(_0542_),
    .B1(_0547_),
    .C1(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__a21o_1 _5583_ (.A1(_0510_),
    .A2(_0543_),
    .B1(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__buf_2 _5584_ (.A(_0494_),
    .X(_0557_));
 sky130_fd_sc_hd__o21ai_1 _5585_ (.A1(_0545_),
    .A2(_0556_),
    .B1(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__mux2_1 _5586_ (.A0(_0491_),
    .A1(_0471_),
    .S(_0480_),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_1 _5587_ (.A0(_0477_),
    .A1(_0544_),
    .S(_0480_),
    .X(_0560_));
 sky130_fd_sc_hd__mux2_1 _5588_ (.A0(_0559_),
    .A1(_0560_),
    .S(_0535_),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_1 _5589_ (.A0(_0533_),
    .A1(_0541_),
    .S(_0480_),
    .X(_0562_));
 sky130_fd_sc_hd__and2_1 _5590_ (.A(_0535_),
    .B(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _5591_ (.A0(_0530_),
    .A1(_0532_),
    .S(_0480_),
    .X(_0564_));
 sky130_fd_sc_hd__and2_1 _5592_ (.A(_0494_),
    .B(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__or4_1 _5593_ (.A(_0519_),
    .B(_0561_),
    .C(_0563_),
    .D(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _5594_ (.A0(_0507_),
    .A1(_0487_),
    .S(_0515_),
    .X(_0567_));
 sky130_fd_sc_hd__clkinv_2 _5595_ (.A(_0514_),
    .Y(_0568_));
 sky130_fd_sc_hd__mux2_1 _5596_ (.A0(_0568_),
    .A1(_0503_),
    .S(_0515_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_1 _5597_ (.A0(_0567_),
    .A1(_0569_),
    .S(_0494_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _5598_ (.A0(_0523_),
    .A1(_0529_),
    .S(_0515_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _5599_ (.A0(_0526_),
    .A1(_0522_),
    .S(_0515_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_1 _5600_ (.A0(_0571_),
    .A1(_0572_),
    .S(_0557_),
    .X(_0573_));
 sky130_fd_sc_hd__nand2_1 _5601_ (.A(_0535_),
    .B(_0479_),
    .Y(_0574_));
 sky130_fd_sc_hd__inv_2 _5602_ (.A(_0574_),
    .Y(_0575_));
 sky130_fd_sc_hd__mux2_1 _5603_ (.A0(_0555_),
    .A1(_0543_),
    .S(_0510_),
    .X(_0576_));
 sky130_fd_sc_hd__or2_1 _5604_ (.A(_0494_),
    .B(_0556_),
    .X(_0577_));
 sky130_fd_sc_hd__a21o_1 _5605_ (.A1(_0574_),
    .A2(_0577_),
    .B1(_0545_),
    .X(_0578_));
 sky130_fd_sc_hd__or4_1 _5606_ (.A(_0535_),
    .B(_0481_),
    .C(_0534_),
    .D(_0562_),
    .X(_0579_));
 sky130_fd_sc_hd__a22o_1 _5607_ (.A1(_0575_),
    .A2(_0576_),
    .B1(_0578_),
    .B2(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__or4_1 _5608_ (.A(_0521_),
    .B(_0570_),
    .C(_0573_),
    .D(_0580_),
    .X(_0581_));
 sky130_fd_sc_hd__a32o_1 _5609_ (.A1(_0510_),
    .A2(_0555_),
    .A3(_0575_),
    .B1(_0560_),
    .B2(_0557_),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _5610_ (.A0(_0567_),
    .A1(_0559_),
    .S(_0535_),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _5611_ (.A0(_0531_),
    .A1(_0524_),
    .S(_0494_),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_1 _5612_ (.A0(_0571_),
    .A1(_0564_),
    .S(_0535_),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_1 _5613_ (.A0(_0492_),
    .A1(_0508_),
    .S(_0494_),
    .X(_0586_));
 sky130_fd_sc_hd__or4_1 _5614_ (.A(_0495_),
    .B(_0586_),
    .C(_0561_),
    .D(_0536_),
    .X(_0587_));
 sky130_fd_sc_hd__or4_1 _5615_ (.A(_0521_),
    .B(_0563_),
    .C(_0565_),
    .D(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__or4_1 _5616_ (.A(_0583_),
    .B(_0584_),
    .C(_0585_),
    .D(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__o31a_1 _5617_ (.A1(_0519_),
    .A2(_0580_),
    .A3(_0582_),
    .B1(_0589_),
    .X(_0590_));
 sky130_fd_sc_hd__a21oi_1 _5618_ (.A1(_0566_),
    .A2(_0581_),
    .B1(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__a32o_1 _5619_ (.A1(_0441_),
    .A2(_0455_),
    .A3(_0518_),
    .B1(_0519_),
    .B2(_0557_),
    .X(_0592_));
 sky130_fd_sc_hd__a31o_1 _5620_ (.A1(_0538_),
    .A2(_0558_),
    .A3(_0591_),
    .B1(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__and2b_1 _5621_ (.A_N(_0520_),
    .B(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__or3_1 _5622_ (.A(_0592_),
    .B(_0538_),
    .C(_0520_),
    .X(_0595_));
 sky130_fd_sc_hd__o21ai_1 _5623_ (.A1(_0593_),
    .A2(_0520_),
    .B1(_0538_),
    .Y(_0596_));
 sky130_fd_sc_hd__and2_1 _5624_ (.A(_0595_),
    .B(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__a21oi_1 _5625_ (.A1(_1330_),
    .A2(_0594_),
    .B1(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__or3b_4 _5626_ (.A(_0092_),
    .B(\cmd[7] ),
    .C_N(\cmd[6] ),
    .X(_0599_));
 sky130_fd_sc_hd__clkbuf_4 _5627_ (.A(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__buf_2 _5628_ (.A(_1319_),
    .X(_0601_));
 sky130_fd_sc_hd__and3b_1 _5629_ (.A_N(_0538_),
    .B(_0594_),
    .C(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__or2_1 _5630_ (.A(_0356_),
    .B(_0363_),
    .X(_0603_));
 sky130_fd_sc_hd__a21oi_4 _5631_ (.A1(_1737_),
    .A2(_2507_),
    .B1(_3775_),
    .Y(_0604_));
 sky130_fd_sc_hd__a21o_1 _5632_ (.A1(_3814_),
    .A2(_0604_),
    .B1(_3699_),
    .X(_0605_));
 sky130_fd_sc_hd__a21o_1 _5633_ (.A1(_3699_),
    .A2(_3814_),
    .B1(_0112_),
    .X(_0606_));
 sky130_fd_sc_hd__o2bb2a_2 _5634_ (.A1_N(_3759_),
    .A2_N(_3760_),
    .B1(_3898_),
    .B2(_3899_),
    .X(_0607_));
 sky130_fd_sc_hd__nor2_1 _5635_ (.A(_0112_),
    .B(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__a21o_2 _5636_ (.A1(_1748_),
    .A2(_2507_),
    .B1(_3775_),
    .X(_0609_));
 sky130_fd_sc_hd__a31o_1 _5637_ (.A1(_3865_),
    .A2(_3900_),
    .A3(_0609_),
    .B1(_3801_),
    .X(_0610_));
 sky130_fd_sc_hd__a32o_1 _5638_ (.A1(_3762_),
    .A2(_0605_),
    .A3(_0606_),
    .B1(_0608_),
    .B2(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__nand2_1 _5639_ (.A(_3900_),
    .B(_0609_),
    .Y(_0612_));
 sky130_fd_sc_hd__nor2_2 _5640_ (.A(_0112_),
    .B(_3864_),
    .Y(_0613_));
 sky130_fd_sc_hd__or3_2 _5641_ (.A(_4043_),
    .B(_3898_),
    .C(_3899_),
    .X(_0614_));
 sky130_fd_sc_hd__o2111a_1 _5642_ (.A1(_3900_),
    .A2(_0609_),
    .B1(_0614_),
    .C1(_3864_),
    .D1(_3718_),
    .X(_0615_));
 sky130_fd_sc_hd__nand2_2 _5643_ (.A(_2507_),
    .B(_3775_),
    .Y(_0616_));
 sky130_fd_sc_hd__a221oi_1 _5644_ (.A1(_0616_),
    .A2(_0607_),
    .B1(_0614_),
    .B2(_3864_),
    .C1(_3718_),
    .Y(_0617_));
 sky130_fd_sc_hd__a2111o_1 _5645_ (.A1(_0612_),
    .A2(_0613_),
    .B1(_0615_),
    .C1(_0617_),
    .D1(_3801_),
    .X(_0618_));
 sky130_fd_sc_hd__a22o_2 _5646_ (.A1(_3811_),
    .A2(_3812_),
    .B1(_3775_),
    .B2(_2507_),
    .X(_0619_));
 sky130_fd_sc_hd__and2_1 _5647_ (.A(_3865_),
    .B(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__nor2_1 _5648_ (.A(_3865_),
    .B(_0619_),
    .Y(_0621_));
 sky130_fd_sc_hd__a21o_1 _5649_ (.A1(_3717_),
    .A2(_0607_),
    .B1(_3699_),
    .X(_0622_));
 sky130_fd_sc_hd__o31a_1 _5650_ (.A1(_0620_),
    .A2(_0621_),
    .A3(_0622_),
    .B1(_3923_),
    .X(_0623_));
 sky130_fd_sc_hd__a22o_2 _5651_ (.A1(_4221_),
    .A2(_0611_),
    .B1(_0618_),
    .B2(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__nand2_1 _5652_ (.A(_3901_),
    .B(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__a21oi_2 _5653_ (.A1(_3864_),
    .A2(_0619_),
    .B1(_0112_),
    .Y(_0626_));
 sky130_fd_sc_hd__o21ai_4 _5654_ (.A1(_3699_),
    .A2(_0626_),
    .B1(_3923_),
    .Y(_0627_));
 sky130_fd_sc_hd__a211o_1 _5655_ (.A1(_3864_),
    .A2(_0619_),
    .B1(_3699_),
    .C1(_0111_),
    .X(_0628_));
 sky130_fd_sc_hd__a211o_1 _5656_ (.A1(_0616_),
    .A2(_0607_),
    .B1(_3801_),
    .C1(_3717_),
    .X(_0629_));
 sky130_fd_sc_hd__o311a_1 _5657_ (.A1(_3761_),
    .A2(_3813_),
    .A3(_0604_),
    .B1(_3717_),
    .C1(_3699_),
    .X(_0630_));
 sky130_fd_sc_hd__a31o_2 _5658_ (.A1(_3923_),
    .A2(_0628_),
    .A3(_0629_),
    .B1(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__or4b_1 _5659_ (.A(_3792_),
    .B(_0627_),
    .C(_3735_),
    .D_N(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__o21a_2 _5660_ (.A1(_3700_),
    .A2(_0626_),
    .B1(_3923_),
    .X(_0633_));
 sky130_fd_sc_hd__buf_2 _5661_ (.A(_0631_),
    .X(_0634_));
 sky130_fd_sc_hd__a22o_1 _5662_ (.A1(_0633_),
    .A2(_3892_),
    .B1(_0634_),
    .B2(_3775_),
    .X(_0636_));
 sky130_fd_sc_hd__nand2_1 _5663_ (.A(_0632_),
    .B(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__xnor2_1 _5664_ (.A(_0625_),
    .B(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__or4b_1 _5665_ (.A(_0627_),
    .B(_3734_),
    .C(_3770_),
    .D_N(_0631_),
    .X(_0639_));
 sky130_fd_sc_hd__a22o_1 _5666_ (.A1(_0633_),
    .A2(_3878_),
    .B1(_0631_),
    .B2(_3892_),
    .X(_0640_));
 sky130_fd_sc_hd__nand4_1 _5667_ (.A(_4045_),
    .B(_0639_),
    .C(_0624_),
    .D(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__nand2_1 _5668_ (.A(_0639_),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__or2b_1 _5669_ (.A(_0638_),
    .B_N(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__xnor2_1 _5670_ (.A(_0642_),
    .B(_0638_),
    .Y(_0644_));
 sky130_fd_sc_hd__a21oi_1 _5671_ (.A1(_0619_),
    .A2(_0614_),
    .B1(_3761_),
    .Y(_0645_));
 sky130_fd_sc_hd__a31o_1 _5672_ (.A1(_1990_),
    .A2(_3713_),
    .A3(_3715_),
    .B1(_3774_),
    .X(_0647_));
 sky130_fd_sc_hd__a221o_1 _5673_ (.A1(_4043_),
    .A2(_0647_),
    .B1(_3811_),
    .B2(_3812_),
    .C1(_3678_),
    .X(_0648_));
 sky130_fd_sc_hd__a21oi_1 _5674_ (.A1(_0616_),
    .A2(_0648_),
    .B1(_3865_),
    .Y(_0649_));
 sky130_fd_sc_hd__a21o_1 _5675_ (.A1(_3900_),
    .A2(_0609_),
    .B1(_3717_),
    .X(_0650_));
 sky130_fd_sc_hd__nor2_1 _5676_ (.A(_3900_),
    .B(_0609_),
    .Y(_0651_));
 sky130_fd_sc_hd__o32a_1 _5677_ (.A1(_0112_),
    .A2(_0645_),
    .A3(_0649_),
    .B1(_0650_),
    .B2(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__o211a_1 _5678_ (.A1(_3813_),
    .A2(_0604_),
    .B1(_0619_),
    .C1(_3761_),
    .X(_0653_));
 sky130_fd_sc_hd__o31ai_1 _5679_ (.A1(_3718_),
    .A2(_0645_),
    .A3(_0653_),
    .B1(_3699_),
    .Y(_0654_));
 sky130_fd_sc_hd__o21a_1 _5680_ (.A1(_3813_),
    .A2(_0604_),
    .B1(_0619_),
    .X(_0655_));
 sky130_fd_sc_hd__or3_1 _5681_ (.A(_2507_),
    .B(_3864_),
    .C(_3813_),
    .X(_0656_));
 sky130_fd_sc_hd__a21oi_1 _5682_ (.A1(_0604_),
    .A2(_0607_),
    .B1(_0112_),
    .Y(_0658_));
 sky130_fd_sc_hd__o211a_1 _5683_ (.A1(_3762_),
    .A2(_0655_),
    .B1(_0656_),
    .C1(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__o22a_1 _5684_ (.A1(_3700_),
    .A2(_0652_),
    .B1(_0654_),
    .B2(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__a21oi_1 _5685_ (.A1(_3814_),
    .A2(_3791_),
    .B1(_2518_),
    .Y(_0661_));
 sky130_fd_sc_hd__o21a_1 _5686_ (.A1(_0651_),
    .A2(_0661_),
    .B1(_0613_),
    .X(_0662_));
 sky130_fd_sc_hd__nand2_1 _5687_ (.A(_0616_),
    .B(_0609_),
    .Y(_0663_));
 sky130_fd_sc_hd__nor2_1 _5688_ (.A(_0613_),
    .B(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__nor2_1 _5689_ (.A(_4043_),
    .B(_3791_),
    .Y(_0665_));
 sky130_fd_sc_hd__or2_1 _5690_ (.A(_0665_),
    .B(_0648_),
    .X(_0666_));
 sky130_fd_sc_hd__a21o_1 _5691_ (.A1(_0616_),
    .A2(_0609_),
    .B1(_3814_),
    .X(_0667_));
 sky130_fd_sc_hd__a211oi_1 _5692_ (.A1(_0666_),
    .A2(_0667_),
    .B1(_3718_),
    .C1(_3865_),
    .Y(_0669_));
 sky130_fd_sc_hd__mux2_1 _5693_ (.A0(_0365_),
    .A1(_3791_),
    .S(_3813_),
    .X(_0670_));
 sky130_fd_sc_hd__a21o_1 _5694_ (.A1(_0616_),
    .A2(_0609_),
    .B1(_3717_),
    .X(_0671_));
 sky130_fd_sc_hd__o2111a_1 _5695_ (.A1(_3900_),
    .A2(_4044_),
    .B1(_0647_),
    .C1(_3717_),
    .D1(_3761_),
    .X(_0672_));
 sky130_fd_sc_hd__a311o_1 _5696_ (.A1(_3865_),
    .A2(_0670_),
    .A3(_0671_),
    .B1(_0672_),
    .C1(_3801_),
    .X(_0673_));
 sky130_fd_sc_hd__o32a_1 _5697_ (.A1(_3700_),
    .A2(_0662_),
    .A3(_0664_),
    .B1(_0669_),
    .B2(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _5698_ (.A0(_0660_),
    .A1(_0674_),
    .S(_3924_),
    .X(_0675_));
 sky130_fd_sc_hd__buf_2 _5699_ (.A(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__nor2_1 _5700_ (.A(_3719_),
    .B(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__o221a_1 _5701_ (.A1(_0112_),
    .A2(_3865_),
    .B1(_3791_),
    .B2(_0614_),
    .C1(_0619_),
    .X(_0678_));
 sky130_fd_sc_hd__a21oi_1 _5702_ (.A1(_0613_),
    .A2(_0648_),
    .B1(_0678_),
    .Y(_0680_));
 sky130_fd_sc_hd__nand2_1 _5703_ (.A(_3814_),
    .B(_3791_),
    .Y(_0681_));
 sky130_fd_sc_hd__and3_1 _5704_ (.A(_3717_),
    .B(_3864_),
    .C(_0614_),
    .X(_0682_));
 sky130_fd_sc_hd__a32o_1 _5705_ (.A1(_0681_),
    .A2(_0613_),
    .A3(_0663_),
    .B1(_0666_),
    .B2(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__o22a_1 _5706_ (.A1(_3700_),
    .A2(_0680_),
    .B1(_0683_),
    .B2(_0654_),
    .X(_0684_));
 sky130_fd_sc_hd__nand2_1 _5707_ (.A(_3762_),
    .B(_3900_),
    .Y(_0685_));
 sky130_fd_sc_hd__a31o_1 _5708_ (.A1(_3718_),
    .A2(_0612_),
    .A3(_0685_),
    .B1(_0617_),
    .X(_0686_));
 sky130_fd_sc_hd__and2_2 _5709_ (.A(_0604_),
    .B(_0607_),
    .X(_0687_));
 sky130_fd_sc_hd__a21oi_1 _5710_ (.A1(_3814_),
    .A2(_0604_),
    .B1(_3762_),
    .Y(_0688_));
 sky130_fd_sc_hd__a211o_1 _5711_ (.A1(_3864_),
    .A2(_0619_),
    .B1(_0607_),
    .C1(_0112_),
    .X(_0689_));
 sky130_fd_sc_hd__o311a_1 _5712_ (.A1(_3718_),
    .A2(_0687_),
    .A3(_0688_),
    .B1(_0689_),
    .C1(_3801_),
    .X(_0691_));
 sky130_fd_sc_hd__a211o_1 _5713_ (.A1(_3700_),
    .A2(_0686_),
    .B1(_0691_),
    .C1(_3923_),
    .X(_0692_));
 sky130_fd_sc_hd__o21a_1 _5714_ (.A1(_4222_),
    .A2(_0684_),
    .B1(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__and2b_1 _5715_ (.A_N(_0630_),
    .B(_0622_),
    .X(_0694_));
 sky130_fd_sc_hd__and3_1 _5716_ (.A(_0111_),
    .B(_3864_),
    .C(_0619_),
    .X(_0695_));
 sky130_fd_sc_hd__o31a_1 _5717_ (.A1(_3699_),
    .A2(_0626_),
    .A3(_0695_),
    .B1(_3923_),
    .X(_0696_));
 sky130_fd_sc_hd__nor2_1 _5718_ (.A(_3762_),
    .B(_0614_),
    .Y(_0697_));
 sky130_fd_sc_hd__nand2_1 _5719_ (.A(_3699_),
    .B(_3718_),
    .Y(_0698_));
 sky130_fd_sc_hd__o22a_1 _5720_ (.A1(_0629_),
    .A2(_0697_),
    .B1(_0688_),
    .B2(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__a2bb2o_1 _5721_ (.A1_N(_3923_),
    .A2_N(_0694_),
    .B1(_0696_),
    .B2(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__clkbuf_4 _5722_ (.A(_0700_),
    .X(_0702_));
 sky130_fd_sc_hd__nor2_1 _5723_ (.A(_2529_),
    .B(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__or3b_1 _5724_ (.A(_3762_),
    .B(_0693_),
    .C_N(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__o21ai_1 _5725_ (.A1(_4222_),
    .A2(_0684_),
    .B1(_0692_),
    .Y(_0705_));
 sky130_fd_sc_hd__clkbuf_4 _5726_ (.A(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__a21o_1 _5727_ (.A1(_3866_),
    .A2(_0706_),
    .B1(_0703_),
    .X(_0707_));
 sky130_fd_sc_hd__nand3_1 _5728_ (.A(_0677_),
    .B(_0704_),
    .C(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__a21o_1 _5729_ (.A1(_0704_),
    .A2(_0707_),
    .B1(_0677_),
    .X(_0709_));
 sky130_fd_sc_hd__nand3_1 _5730_ (.A(_0644_),
    .B(_0708_),
    .C(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__o21ai_1 _5731_ (.A1(_0625_),
    .A2(_0637_),
    .B1(_0632_),
    .Y(_0711_));
 sky130_fd_sc_hd__nand2_1 _5732_ (.A(_3866_),
    .B(_0624_),
    .Y(_0713_));
 sky130_fd_sc_hd__nand2_1 _5733_ (.A(_3775_),
    .B(_0634_),
    .Y(_0714_));
 sky130_fd_sc_hd__nand2_1 _5734_ (.A(_4045_),
    .B(_0633_),
    .Y(_0715_));
 sky130_fd_sc_hd__a22o_1 _5735_ (.A1(_3775_),
    .A2(_0633_),
    .B1(_0631_),
    .B2(_4044_),
    .X(_0716_));
 sky130_fd_sc_hd__o21ai_1 _5736_ (.A1(_0714_),
    .A2(_0715_),
    .B1(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__xor2_1 _5737_ (.A(_0713_),
    .B(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__xor2_1 _5738_ (.A(_0711_),
    .B(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__nor2_1 _5739_ (.A(_3700_),
    .B(_0676_),
    .Y(_0720_));
 sky130_fd_sc_hd__or4_2 _5740_ (.A(_3719_),
    .B(_3815_),
    .C(_0702_),
    .D(_0693_),
    .X(_0721_));
 sky130_fd_sc_hd__inv_2 _5741_ (.A(_0700_),
    .Y(_0722_));
 sky130_fd_sc_hd__a22o_1 _5742_ (.A1(_3901_),
    .A2(_0722_),
    .B1(_0705_),
    .B2(_0113_),
    .X(_0724_));
 sky130_fd_sc_hd__nand3_1 _5743_ (.A(_0720_),
    .B(_0721_),
    .C(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__a21o_1 _5744_ (.A1(_0721_),
    .A2(_0724_),
    .B1(_0720_),
    .X(_0726_));
 sky130_fd_sc_hd__and3_1 _5745_ (.A(_0719_),
    .B(_0725_),
    .C(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__a21oi_1 _5746_ (.A1(_0725_),
    .A2(_0726_),
    .B1(_0719_),
    .Y(_0728_));
 sky130_fd_sc_hd__a211oi_1 _5747_ (.A1(_0643_),
    .A2(_0710_),
    .B1(_0727_),
    .C1(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__o211a_1 _5748_ (.A1(_0727_),
    .A2(_0728_),
    .B1(_0643_),
    .C1(_0710_),
    .X(_0730_));
 sky130_fd_sc_hd__a21boi_1 _5749_ (.A1(_0677_),
    .A2(_0707_),
    .B1_N(_0704_),
    .Y(_0731_));
 sky130_fd_sc_hd__a21o_1 _5750_ (.A1(_0647_),
    .A2(_4044_),
    .B1(_3814_),
    .X(_0732_));
 sky130_fd_sc_hd__a21o_1 _5751_ (.A1(_0666_),
    .A2(_0732_),
    .B1(_3762_),
    .X(_0733_));
 sky130_fd_sc_hd__a211o_1 _5752_ (.A1(_0365_),
    .A2(_3901_),
    .B1(_2529_),
    .C1(_3866_),
    .X(_0734_));
 sky130_fd_sc_hd__a21oi_1 _5753_ (.A1(_0616_),
    .A2(_0648_),
    .B1(_3762_),
    .Y(_0735_));
 sky130_fd_sc_hd__o21a_1 _5754_ (.A1(_0687_),
    .A2(_0735_),
    .B1(_3718_),
    .X(_0736_));
 sky130_fd_sc_hd__a311o_1 _5755_ (.A1(_0113_),
    .A2(_0733_),
    .A3(_0734_),
    .B1(_0736_),
    .C1(_4222_),
    .X(_0737_));
 sky130_fd_sc_hd__or3_1 _5756_ (.A(_0365_),
    .B(_3900_),
    .C(_2518_),
    .X(_0738_));
 sky130_fd_sc_hd__a211oi_1 _5757_ (.A1(_2507_),
    .A2(_3815_),
    .B1(_0670_),
    .C1(_3866_),
    .Y(_0739_));
 sky130_fd_sc_hd__a31o_1 _5758_ (.A1(_3866_),
    .A2(_0667_),
    .A3(_0738_),
    .B1(_0739_),
    .X(_0740_));
 sky130_fd_sc_hd__a21o_1 _5759_ (.A1(_0666_),
    .A2(_0667_),
    .B1(_3865_),
    .X(_0741_));
 sky130_fd_sc_hd__a21o_1 _5760_ (.A1(_0732_),
    .A2(_0738_),
    .B1(_3762_),
    .X(_0742_));
 sky130_fd_sc_hd__and3_1 _5761_ (.A(_0113_),
    .B(_0741_),
    .C(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__a211o_1 _5762_ (.A1(_3719_),
    .A2(_0740_),
    .B1(_0743_),
    .C1(_3924_),
    .X(_0745_));
 sky130_fd_sc_hd__nor2_1 _5763_ (.A(_3866_),
    .B(_0670_),
    .Y(_0746_));
 sky130_fd_sc_hd__a21o_1 _5764_ (.A1(_3814_),
    .A2(_2518_),
    .B1(_0365_),
    .X(_0747_));
 sky130_fd_sc_hd__a21o_1 _5765_ (.A1(_3865_),
    .A2(_0747_),
    .B1(_0112_),
    .X(_0748_));
 sky130_fd_sc_hd__o221a_1 _5766_ (.A1(_3718_),
    .A2(_3775_),
    .B1(_0746_),
    .B2(_0748_),
    .C1(_3924_),
    .X(_0749_));
 sky130_fd_sc_hd__a22o_1 _5767_ (.A1(_2507_),
    .A2(_3815_),
    .B1(_3792_),
    .B2(_0732_),
    .X(_0750_));
 sky130_fd_sc_hd__nand2_1 _5768_ (.A(_3814_),
    .B(_0665_),
    .Y(_0751_));
 sky130_fd_sc_hd__a221o_1 _5769_ (.A1(_0113_),
    .A2(_0663_),
    .B1(_0751_),
    .B2(_0615_),
    .C1(_3924_),
    .X(_0752_));
 sky130_fd_sc_hd__a21oi_1 _5770_ (.A1(_0613_),
    .A2(_0750_),
    .B1(_0752_),
    .Y(_0753_));
 sky130_fd_sc_hd__o21a_2 _5771_ (.A1(_0749_),
    .A2(_0753_),
    .B1(_3802_),
    .X(_0754_));
 sky130_fd_sc_hd__a31oi_4 _5772_ (.A1(_3700_),
    .A2(_0737_),
    .A3(_0745_),
    .B1(_0754_),
    .Y(_0755_));
 sky130_fd_sc_hd__nor2_1 _5773_ (.A(_3924_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__xor2_1 _5774_ (.A(_0731_),
    .B(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__xnor2_1 _5775_ (.A(_3735_),
    .B(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__or3_1 _5776_ (.A(_0729_),
    .B(_0730_),
    .C(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__and2b_1 _5777_ (.A_N(_0729_),
    .B(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__a21o_1 _5778_ (.A1(_0711_),
    .A2(_0718_),
    .B1(_0727_),
    .X(_0761_));
 sky130_fd_sc_hd__clkbuf_4 _5779_ (.A(_0624_),
    .X(_0762_));
 sky130_fd_sc_hd__nor2_1 _5780_ (.A(_0714_),
    .B(_0715_),
    .Y(_0763_));
 sky130_fd_sc_hd__a31o_1 _5781_ (.A1(_3866_),
    .A2(_0762_),
    .A3(_0716_),
    .B1(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__nand2_1 _5782_ (.A(_0113_),
    .B(_0762_),
    .Y(_0766_));
 sky130_fd_sc_hd__nand2_1 _5783_ (.A(_3901_),
    .B(_0634_),
    .Y(_0767_));
 sky130_fd_sc_hd__xor2_1 _5784_ (.A(_0715_),
    .B(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__xnor2_2 _5785_ (.A(_0766_),
    .B(_0768_),
    .Y(_0769_));
 sky130_fd_sc_hd__xnor2_1 _5786_ (.A(_0764_),
    .B(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__or2_1 _5787_ (.A(_3924_),
    .B(_0660_),
    .X(_0771_));
 sky130_fd_sc_hd__nor2_1 _5788_ (.A(_3763_),
    .B(_0702_),
    .Y(_0772_));
 sky130_fd_sc_hd__clkbuf_4 _5789_ (.A(_0693_),
    .X(_0773_));
 sky130_fd_sc_hd__nor2_1 _5790_ (.A(_3700_),
    .B(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__xnor2_1 _5791_ (.A(_0772_),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__xnor2_1 _5792_ (.A(_0771_),
    .B(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__xor2_1 _5793_ (.A(_0770_),
    .B(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__xnor2_1 _5794_ (.A(_0761_),
    .B(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__or2_2 _5795_ (.A(_4016_),
    .B(_0755_),
    .X(_0779_));
 sky130_fd_sc_hd__a21o_1 _5796_ (.A1(_0721_),
    .A2(_0725_),
    .B1(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__nand3_1 _5797_ (.A(_0721_),
    .B(_0725_),
    .C(_0779_),
    .Y(_0781_));
 sky130_fd_sc_hd__nand2_1 _5798_ (.A(_0780_),
    .B(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__xnor2_1 _5799_ (.A(_3792_),
    .B(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__xnor2_1 _5800_ (.A(_0778_),
    .B(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__xnor2_1 _5801_ (.A(_0760_),
    .B(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__buf_2 _5802_ (.A(_0755_),
    .X(_0787_));
 sky130_fd_sc_hd__or3_1 _5803_ (.A(_3924_),
    .B(_0731_),
    .C(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__o21ai_1 _5804_ (.A1(_3735_),
    .A2(_0757_),
    .B1(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__or2b_1 _5805_ (.A(_0785_),
    .B_N(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__o21a_1 _5806_ (.A1(_0760_),
    .A2(_0784_),
    .B1(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__or2b_1 _5807_ (.A(_0766_),
    .B_N(_0768_),
    .X(_0792_));
 sky130_fd_sc_hd__o21a_1 _5808_ (.A1(_0715_),
    .A2(_0767_),
    .B1(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__nand2_1 _5809_ (.A(_3802_),
    .B(_0762_),
    .Y(_0794_));
 sky130_fd_sc_hd__clkbuf_4 _5810_ (.A(_0633_),
    .X(_0795_));
 sky130_fd_sc_hd__a22o_1 _5811_ (.A1(_3901_),
    .A2(_0795_),
    .B1(_0634_),
    .B2(_3866_),
    .X(_0796_));
 sky130_fd_sc_hd__or4b_1 _5812_ (.A(_3763_),
    .B(_3815_),
    .C(_0627_),
    .D_N(_0634_),
    .X(_0798_));
 sky130_fd_sc_hd__nand2_1 _5813_ (.A(_0796_),
    .B(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__xnor2_1 _5814_ (.A(_0794_),
    .B(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__xnor2_1 _5815_ (.A(_0793_),
    .B(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__buf_2 _5816_ (.A(_0676_),
    .X(_0802_));
 sky130_fd_sc_hd__or2_2 _5817_ (.A(_4016_),
    .B(_0802_),
    .X(_0803_));
 sky130_fd_sc_hd__o21a_1 _5818_ (.A1(_3719_),
    .A2(_0702_),
    .B1(_0692_),
    .X(_0804_));
 sky130_fd_sc_hd__a41o_1 _5819_ (.A1(_4222_),
    .A2(_3700_),
    .A3(_0113_),
    .A4(_0706_),
    .B1(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__xnor2_1 _5820_ (.A(_0803_),
    .B(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__o2bb2ai_1 _5821_ (.A1_N(_0772_),
    .A2_N(_0774_),
    .B1(_0775_),
    .B2(_0771_),
    .Y(_0807_));
 sky130_fd_sc_hd__xnor2_1 _5822_ (.A(_0806_),
    .B(_0807_),
    .Y(_0809_));
 sky130_fd_sc_hd__xnor2_1 _5823_ (.A(_0801_),
    .B(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__nor2_1 _5824_ (.A(_0770_),
    .B(_0776_),
    .Y(_0811_));
 sky130_fd_sc_hd__a21oi_1 _5825_ (.A1(_0764_),
    .A2(_0769_),
    .B1(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__xnor2_1 _5826_ (.A(_2529_),
    .B(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__xnor2_1 _5827_ (.A(_0810_),
    .B(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__o21ai_1 _5828_ (.A1(_3792_),
    .A2(_0782_),
    .B1(_0780_),
    .Y(_0815_));
 sky130_fd_sc_hd__nand2_1 _5829_ (.A(_0761_),
    .B(_0777_),
    .Y(_0816_));
 sky130_fd_sc_hd__o21a_1 _5830_ (.A1(_0778_),
    .A2(_0783_),
    .B1(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__xnor2_1 _5831_ (.A(_0815_),
    .B(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__xnor2_1 _5832_ (.A(_0814_),
    .B(_0818_),
    .Y(_0820_));
 sky130_fd_sc_hd__xnor2_1 _5833_ (.A(_0791_),
    .B(_0820_),
    .Y(_0821_));
 sky130_fd_sc_hd__nor2_1 _5834_ (.A(_3763_),
    .B(_0676_),
    .Y(_0822_));
 sky130_fd_sc_hd__or2_1 _5835_ (.A(_3792_),
    .B(_0700_),
    .X(_0823_));
 sky130_fd_sc_hd__o21ai_1 _5836_ (.A1(_3815_),
    .A2(_0693_),
    .B1(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__or3_1 _5837_ (.A(_3815_),
    .B(_0693_),
    .C(_0823_),
    .X(_0825_));
 sky130_fd_sc_hd__a21boi_1 _5838_ (.A1(_0822_),
    .A2(_0824_),
    .B1_N(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__and2b_1 _5839_ (.A_N(_0826_),
    .B(_0754_),
    .X(_0827_));
 sky130_fd_sc_hd__xor2_1 _5840_ (.A(_0754_),
    .B(_0826_),
    .X(_0828_));
 sky130_fd_sc_hd__nor2_1 _5841_ (.A(_3770_),
    .B(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__or4b_1 _5842_ (.A(_0627_),
    .B(_3770_),
    .C(_3738_),
    .D_N(_0631_),
    .X(_0831_));
 sky130_fd_sc_hd__a22o_1 _5843_ (.A1(_3877_),
    .A2(_0631_),
    .B1(_3832_),
    .B2(_0633_),
    .X(_0832_));
 sky130_fd_sc_hd__nand4_1 _5844_ (.A(_3776_),
    .B(_0624_),
    .C(_0831_),
    .D(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__nand2_1 _5845_ (.A(_0831_),
    .B(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__a22o_1 _5846_ (.A1(_4045_),
    .A2(_0624_),
    .B1(_0640_),
    .B2(_0639_),
    .X(_0835_));
 sky130_fd_sc_hd__nand2_1 _5847_ (.A(_0641_),
    .B(_0835_),
    .Y(_0836_));
 sky130_fd_sc_hd__xnor2_1 _5848_ (.A(_0834_),
    .B(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__nand3_1 _5849_ (.A(_0822_),
    .B(_0825_),
    .C(_0824_),
    .Y(_0838_));
 sky130_fd_sc_hd__a21o_1 _5850_ (.A1(_0825_),
    .A2(_0824_),
    .B1(_0822_),
    .X(_0839_));
 sky130_fd_sc_hd__and3_1 _5851_ (.A(_0641_),
    .B(_0834_),
    .C(_0835_),
    .X(_0840_));
 sky130_fd_sc_hd__a31o_1 _5852_ (.A1(_0837_),
    .A2(_0838_),
    .A3(_0839_),
    .B1(_0840_),
    .X(_0842_));
 sky130_fd_sc_hd__a21o_1 _5853_ (.A1(_0708_),
    .A2(_0709_),
    .B1(_0644_),
    .X(_0843_));
 sky130_fd_sc_hd__and3_1 _5854_ (.A(_0710_),
    .B(_0842_),
    .C(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__a21oi_1 _5855_ (.A1(_0710_),
    .A2(_0843_),
    .B1(_0842_),
    .Y(_0845_));
 sky130_fd_sc_hd__xnor2_1 _5856_ (.A(_3770_),
    .B(_0828_),
    .Y(_0846_));
 sky130_fd_sc_hd__nor3_1 _5857_ (.A(_0844_),
    .B(_0845_),
    .C(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__o21ai_1 _5858_ (.A1(_0729_),
    .A2(_0730_),
    .B1(_0758_),
    .Y(_0848_));
 sky130_fd_sc_hd__o211ai_2 _5859_ (.A1(_0844_),
    .A2(_0847_),
    .B1(_0848_),
    .C1(_0759_),
    .Y(_0849_));
 sky130_fd_sc_hd__a211o_1 _5860_ (.A1(_0759_),
    .A2(_0848_),
    .B1(_0847_),
    .C1(_0844_),
    .X(_0850_));
 sky130_fd_sc_hd__o211a_1 _5861_ (.A1(_0827_),
    .A2(_0829_),
    .B1(_0849_),
    .C1(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__a211oi_1 _5862_ (.A1(_0849_),
    .A2(_0850_),
    .B1(_0827_),
    .C1(_0829_),
    .Y(_0852_));
 sky130_fd_sc_hd__nor2_1 _5863_ (.A(_0851_),
    .B(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__nor2_1 _5864_ (.A(_3815_),
    .B(_0676_),
    .Y(_0854_));
 sky130_fd_sc_hd__or2_1 _5865_ (.A(_3735_),
    .B(_0700_),
    .X(_0855_));
 sky130_fd_sc_hd__o21ai_1 _5866_ (.A1(_2529_),
    .A2(_0773_),
    .B1(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__or3_1 _5867_ (.A(_2529_),
    .B(_0693_),
    .C(_0855_),
    .X(_0857_));
 sky130_fd_sc_hd__a21bo_1 _5868_ (.A1(_0854_),
    .A2(_0856_),
    .B1_N(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__nor2_1 _5869_ (.A(_3719_),
    .B(_0755_),
    .Y(_0859_));
 sky130_fd_sc_hd__xnor2_1 _5870_ (.A(_0858_),
    .B(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__nand2_1 _5871_ (.A(_0858_),
    .B(_0859_),
    .Y(_0861_));
 sky130_fd_sc_hd__o21ai_1 _5872_ (.A1(_3738_),
    .A2(_0860_),
    .B1(_0861_),
    .Y(_0863_));
 sky130_fd_sc_hd__or3_1 _5873_ (.A(_0844_),
    .B(_0845_),
    .C(_0846_),
    .X(_0864_));
 sky130_fd_sc_hd__o21ai_1 _5874_ (.A1(_0844_),
    .A2(_0845_),
    .B1(_0846_),
    .Y(_0865_));
 sky130_fd_sc_hd__nand3_1 _5875_ (.A(_0837_),
    .B(_0838_),
    .C(_0839_),
    .Y(_0866_));
 sky130_fd_sc_hd__and4_1 _5876_ (.A(_3892_),
    .B(_0634_),
    .C(_0624_),
    .D(_3832_),
    .X(_0867_));
 sky130_fd_sc_hd__a22o_1 _5877_ (.A1(_3776_),
    .A2(_0624_),
    .B1(_0831_),
    .B2(_0832_),
    .X(_0868_));
 sky130_fd_sc_hd__and2_1 _5878_ (.A(_0833_),
    .B(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__xor2_1 _5879_ (.A(_0867_),
    .B(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__nand3_1 _5880_ (.A(_0854_),
    .B(_0856_),
    .C(_0857_),
    .Y(_0871_));
 sky130_fd_sc_hd__a21o_1 _5881_ (.A1(_0856_),
    .A2(_0857_),
    .B1(_0854_),
    .X(_0872_));
 sky130_fd_sc_hd__and2_1 _5882_ (.A(_0867_),
    .B(_0869_),
    .X(_0873_));
 sky130_fd_sc_hd__a31o_1 _5883_ (.A1(_0870_),
    .A2(_0871_),
    .A3(_0872_),
    .B1(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__a21o_1 _5884_ (.A1(_0838_),
    .A2(_0839_),
    .B1(_0837_),
    .X(_0875_));
 sky130_fd_sc_hd__and3_1 _5885_ (.A(_0866_),
    .B(_0874_),
    .C(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__a21oi_1 _5886_ (.A1(_0866_),
    .A2(_0875_),
    .B1(_0874_),
    .Y(_0877_));
 sky130_fd_sc_hd__xnor2_1 _5887_ (.A(_3738_),
    .B(_0860_),
    .Y(_0878_));
 sky130_fd_sc_hd__nor3_2 _5888_ (.A(_0876_),
    .B(_0877_),
    .C(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__a211o_1 _5889_ (.A1(_0864_),
    .A2(_0865_),
    .B1(_0879_),
    .C1(_0876_),
    .X(_0880_));
 sky130_fd_sc_hd__o211ai_1 _5890_ (.A1(_0876_),
    .A2(_0879_),
    .B1(_0865_),
    .C1(_0864_),
    .Y(_0881_));
 sky130_fd_sc_hd__a21boi_1 _5891_ (.A1(_0863_),
    .A2(_0880_),
    .B1_N(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__xnor2_2 _5892_ (.A(_0853_),
    .B(_0882_),
    .Y(_0884_));
 sky130_fd_sc_hd__or3_1 _5893_ (.A(_0693_),
    .B(_3738_),
    .C(_0855_),
    .X(_0885_));
 sky130_fd_sc_hd__nor2_1 _5894_ (.A(_3792_),
    .B(_0676_),
    .Y(_0886_));
 sky130_fd_sc_hd__a22o_1 _5895_ (.A1(_3892_),
    .A2(_0706_),
    .B1(_3832_),
    .B2(_0722_),
    .X(_0887_));
 sky130_fd_sc_hd__nand3_1 _5896_ (.A(_0885_),
    .B(_0886_),
    .C(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__nand2_1 _5897_ (.A(_0885_),
    .B(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__nor2_1 _5898_ (.A(_3815_),
    .B(_0787_),
    .Y(_0890_));
 sky130_fd_sc_hd__and2_1 _5899_ (.A(_0889_),
    .B(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__clkinv_2 _5900_ (.A(_0762_),
    .Y(_0892_));
 sky130_fd_sc_hd__o2bb2a_1 _5901_ (.A1_N(_0634_),
    .A2_N(_3832_),
    .B1(_0892_),
    .B2(_3735_),
    .X(_0893_));
 sky130_fd_sc_hd__nor2_1 _5902_ (.A(_0867_),
    .B(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__nor2_1 _5903_ (.A(_2529_),
    .B(_0676_),
    .Y(_0895_));
 sky130_fd_sc_hd__or3_1 _5904_ (.A(_3770_),
    .B(_0773_),
    .C(_0823_),
    .X(_0896_));
 sky130_fd_sc_hd__a22o_1 _5905_ (.A1(_3878_),
    .A2(_0722_),
    .B1(_0706_),
    .B2(_3776_),
    .X(_0897_));
 sky130_fd_sc_hd__nand3_1 _5906_ (.A(_0895_),
    .B(_0896_),
    .C(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__a21o_1 _5907_ (.A1(_0896_),
    .A2(_0897_),
    .B1(_0895_),
    .X(_0899_));
 sky130_fd_sc_hd__nand3_1 _5908_ (.A(_0894_),
    .B(_0898_),
    .C(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__a21o_1 _5909_ (.A1(_0898_),
    .A2(_0899_),
    .B1(_0894_),
    .X(_0901_));
 sky130_fd_sc_hd__nor2_1 _5910_ (.A(_3770_),
    .B(_0892_),
    .Y(_0902_));
 sky130_fd_sc_hd__a21o_1 _5911_ (.A1(_0885_),
    .A2(_0887_),
    .B1(_0886_),
    .X(_0903_));
 sky130_fd_sc_hd__and3_1 _5912_ (.A(_0888_),
    .B(_0902_),
    .C(_0903_),
    .X(_0905_));
 sky130_fd_sc_hd__a21o_1 _5913_ (.A1(_0900_),
    .A2(_0901_),
    .B1(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__xor2_1 _5914_ (.A(_0889_),
    .B(_0890_),
    .X(_0907_));
 sky130_fd_sc_hd__nand3_1 _5915_ (.A(_0905_),
    .B(_0900_),
    .C(_0901_),
    .Y(_0908_));
 sky130_fd_sc_hd__a21bo_1 _5916_ (.A1(_0906_),
    .A2(_0907_),
    .B1_N(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__nand2_1 _5917_ (.A(_0896_),
    .B(_0898_),
    .Y(_0910_));
 sky130_fd_sc_hd__nor2_1 _5918_ (.A(_3763_),
    .B(_0787_),
    .Y(_0911_));
 sky130_fd_sc_hd__xor2_1 _5919_ (.A(_0910_),
    .B(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__a21o_1 _5920_ (.A1(_0871_),
    .A2(_0872_),
    .B1(_0870_),
    .X(_0913_));
 sky130_fd_sc_hd__nand3_1 _5921_ (.A(_0870_),
    .B(_0871_),
    .C(_0872_),
    .Y(_0914_));
 sky130_fd_sc_hd__nand3b_2 _5922_ (.A_N(_0900_),
    .B(_0913_),
    .C(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__a21bo_1 _5923_ (.A1(_0914_),
    .A2(_0913_),
    .B1_N(_0900_),
    .X(_0916_));
 sky130_fd_sc_hd__nand3_2 _5924_ (.A(_0912_),
    .B(_0915_),
    .C(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__a21o_1 _5925_ (.A1(_0915_),
    .A2(_0916_),
    .B1(_0912_),
    .X(_0918_));
 sky130_fd_sc_hd__nand3_1 _5926_ (.A(_0909_),
    .B(_0917_),
    .C(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__a21o_1 _5927_ (.A1(_0917_),
    .A2(_0918_),
    .B1(_0909_),
    .X(_0920_));
 sky130_fd_sc_hd__nand3_1 _5928_ (.A(_0891_),
    .B(_0919_),
    .C(_0920_),
    .Y(_0921_));
 sky130_fd_sc_hd__a21o_1 _5929_ (.A1(_0919_),
    .A2(_0920_),
    .B1(_0891_),
    .X(_0922_));
 sky130_fd_sc_hd__nor2_1 _5930_ (.A(_3770_),
    .B(_0773_),
    .Y(_0923_));
 sky130_fd_sc_hd__nor2_1 _5931_ (.A(_3735_),
    .B(_0676_),
    .Y(_0924_));
 sky130_fd_sc_hd__nor2_1 _5932_ (.A(_2529_),
    .B(_0787_),
    .Y(_0926_));
 sky130_fd_sc_hd__and3_1 _5933_ (.A(_0923_),
    .B(_0924_),
    .C(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__nand3_1 _5934_ (.A(_0908_),
    .B(_0906_),
    .C(_0907_),
    .Y(_0928_));
 sky130_fd_sc_hd__a21o_1 _5935_ (.A1(_0908_),
    .A2(_0906_),
    .B1(_0907_),
    .X(_0929_));
 sky130_fd_sc_hd__a21oi_1 _5936_ (.A1(_0888_),
    .A2(_0903_),
    .B1(_0902_),
    .Y(_0930_));
 sky130_fd_sc_hd__nand2_1 _5937_ (.A(_0762_),
    .B(_3832_),
    .Y(_0931_));
 sky130_fd_sc_hd__xnor2_1 _5938_ (.A(_0923_),
    .B(_0924_),
    .Y(_0932_));
 sky130_fd_sc_hd__nor2_1 _5939_ (.A(_0931_),
    .B(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__o21bai_1 _5940_ (.A1(_0905_),
    .A2(_0930_),
    .B1_N(_0933_),
    .Y(_0934_));
 sky130_fd_sc_hd__nand2_1 _5941_ (.A(_0923_),
    .B(_0924_),
    .Y(_0935_));
 sky130_fd_sc_hd__xnor2_1 _5942_ (.A(_0935_),
    .B(_0926_),
    .Y(_0936_));
 sky130_fd_sc_hd__or3b_1 _5943_ (.A(_0905_),
    .B(_0930_),
    .C_N(_0933_),
    .X(_0937_));
 sky130_fd_sc_hd__a21bo_1 _5944_ (.A1(_0934_),
    .A2(_0936_),
    .B1_N(_0937_),
    .X(_0938_));
 sky130_fd_sc_hd__a21o_1 _5945_ (.A1(_0928_),
    .A2(_0929_),
    .B1(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__nand3_1 _5946_ (.A(_0928_),
    .B(_0938_),
    .C(_0929_),
    .Y(_0940_));
 sky130_fd_sc_hd__a21bo_1 _5947_ (.A1(_0927_),
    .A2(_0939_),
    .B1_N(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__a21o_1 _5948_ (.A1(_0921_),
    .A2(_0922_),
    .B1(_0941_),
    .X(_0942_));
 sky130_fd_sc_hd__nand3_1 _5949_ (.A(_0927_),
    .B(_0940_),
    .C(_0939_),
    .Y(_0943_));
 sky130_fd_sc_hd__a21o_1 _5950_ (.A1(_0940_),
    .A2(_0939_),
    .B1(_0927_),
    .X(_0944_));
 sky130_fd_sc_hd__nor2_1 _5951_ (.A(_0773_),
    .B(_3738_),
    .Y(_0945_));
 sky130_fd_sc_hd__nor2_1 _5952_ (.A(_3770_),
    .B(_0802_),
    .Y(_0947_));
 sky130_fd_sc_hd__nor2_1 _5953_ (.A(_3792_),
    .B(_0787_),
    .Y(_0948_));
 sky130_fd_sc_hd__and3_1 _5954_ (.A(_0945_),
    .B(_0947_),
    .C(_0948_),
    .X(_0949_));
 sky130_fd_sc_hd__and2_1 _5955_ (.A(_0931_),
    .B(_0932_),
    .X(_0950_));
 sky130_fd_sc_hd__nor2_1 _5956_ (.A(_0933_),
    .B(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__nand2_1 _5957_ (.A(_0945_),
    .B(_0947_),
    .Y(_0952_));
 sky130_fd_sc_hd__and2b_1 _5958_ (.A_N(_0948_),
    .B(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__nor2_1 _5959_ (.A(_0949_),
    .B(_0953_),
    .Y(_0954_));
 sky130_fd_sc_hd__and2_1 _5960_ (.A(_0951_),
    .B(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__nand3_1 _5961_ (.A(_0937_),
    .B(_0934_),
    .C(_0936_),
    .Y(_0956_));
 sky130_fd_sc_hd__a21o_1 _5962_ (.A1(_0937_),
    .A2(_0934_),
    .B1(_0936_),
    .X(_0957_));
 sky130_fd_sc_hd__and2_1 _5963_ (.A(_0956_),
    .B(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__o21a_1 _5964_ (.A1(_0949_),
    .A2(_0955_),
    .B1(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__and3_1 _5965_ (.A(_0943_),
    .B(_0944_),
    .C(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__and3_1 _5966_ (.A(_0921_),
    .B(_0922_),
    .C(_0941_),
    .X(_0961_));
 sky130_fd_sc_hd__a21oi_2 _5967_ (.A1(_0942_),
    .A2(_0960_),
    .B1(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__nand2_1 _5968_ (.A(_0910_),
    .B(_0911_),
    .Y(_0963_));
 sky130_fd_sc_hd__o21a_1 _5969_ (.A1(_0876_),
    .A2(_0877_),
    .B1(_0878_),
    .X(_0964_));
 sky130_fd_sc_hd__a211oi_1 _5970_ (.A1(_0915_),
    .A2(_0917_),
    .B1(_0964_),
    .C1(_0879_),
    .Y(_0965_));
 sky130_fd_sc_hd__o211a_1 _5971_ (.A1(_0879_),
    .A2(_0964_),
    .B1(_0917_),
    .C1(_0915_),
    .X(_0966_));
 sky130_fd_sc_hd__or3_1 _5972_ (.A(_0963_),
    .B(_0965_),
    .C(_0966_),
    .X(_0968_));
 sky130_fd_sc_hd__o21ai_1 _5973_ (.A1(_0965_),
    .A2(_0966_),
    .B1(_0963_),
    .Y(_0969_));
 sky130_fd_sc_hd__a21bo_1 _5974_ (.A1(_0891_),
    .A2(_0920_),
    .B1_N(_0919_),
    .X(_0970_));
 sky130_fd_sc_hd__and3_1 _5975_ (.A(_0968_),
    .B(_0969_),
    .C(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__a21oi_1 _5976_ (.A1(_0968_),
    .A2(_0969_),
    .B1(_0970_),
    .Y(_0972_));
 sky130_fd_sc_hd__or2_2 _5977_ (.A(_0971_),
    .B(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__a211o_1 _5978_ (.A1(_0915_),
    .A2(_0917_),
    .B1(_0964_),
    .C1(_0879_),
    .X(_0974_));
 sky130_fd_sc_hd__a21oi_1 _5979_ (.A1(_0881_),
    .A2(_0880_),
    .B1(_0863_),
    .Y(_0975_));
 sky130_fd_sc_hd__and3_1 _5980_ (.A(_0881_),
    .B(_0863_),
    .C(_0880_),
    .X(_0976_));
 sky130_fd_sc_hd__a211oi_1 _5981_ (.A1(_0974_),
    .A2(_0968_),
    .B1(_0975_),
    .C1(_0976_),
    .Y(_0977_));
 sky130_fd_sc_hd__o211a_1 _5982_ (.A1(_0976_),
    .A2(_0975_),
    .B1(_0968_),
    .C1(_0974_),
    .X(_0978_));
 sky130_fd_sc_hd__or2_1 _5983_ (.A(_0977_),
    .B(_0978_),
    .X(_0979_));
 sky130_fd_sc_hd__o21bai_1 _5984_ (.A1(_0971_),
    .A2(_0977_),
    .B1_N(_0978_),
    .Y(_0980_));
 sky130_fd_sc_hd__o31ai_4 _5985_ (.A1(_0962_),
    .A2(_0973_),
    .A3(_0979_),
    .B1(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__inv_2 _5986_ (.A(_0849_),
    .Y(_0982_));
 sky130_fd_sc_hd__xnor2_1 _5987_ (.A(_0789_),
    .B(_0785_),
    .Y(_0983_));
 sky130_fd_sc_hd__o21a_1 _5988_ (.A1(_0982_),
    .A2(_0851_),
    .B1(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__or3_1 _5989_ (.A(_0983_),
    .B(_0982_),
    .C(_0851_),
    .X(_0985_));
 sky130_fd_sc_hd__and2b_1 _5990_ (.A_N(_0984_),
    .B(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__and2b_1 _5991_ (.A_N(_0882_),
    .B(_0853_),
    .X(_0987_));
 sky130_fd_sc_hd__o21a_1 _5992_ (.A1(_0984_),
    .A2(_0987_),
    .B1(_0985_),
    .X(_0989_));
 sky130_fd_sc_hd__a31o_1 _5993_ (.A1(_0884_),
    .A2(_0981_),
    .A3(_0986_),
    .B1(_0989_),
    .X(_0990_));
 sky130_fd_sc_hd__xnor2_1 _5994_ (.A(_0821_),
    .B(_0990_),
    .Y(_0991_));
 sky130_fd_sc_hd__buf_2 _5995_ (.A(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__buf_2 _5996_ (.A(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__nor2_4 _5997_ (.A(_4016_),
    .B(_0992_),
    .Y(_0994_));
 sky130_fd_sc_hd__nand2_1 _5998_ (.A(_0795_),
    .B(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__or4_2 _5999_ (.A(_4016_),
    .B(_0892_),
    .C(_0702_),
    .D(_0991_),
    .X(_0996_));
 sky130_fd_sc_hd__a211oi_2 _6000_ (.A1(_0892_),
    .A2(_0702_),
    .B1(_0992_),
    .C1(_4016_),
    .Y(_0997_));
 sky130_fd_sc_hd__nand4_2 _6001_ (.A(_0634_),
    .B(_0994_),
    .C(_0996_),
    .D(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__and3_1 _6002_ (.A(_0995_),
    .B(_0996_),
    .C(_0998_),
    .X(_0999_));
 sky130_fd_sc_hd__clkbuf_2 _6003_ (.A(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__a21oi_1 _6004_ (.A1(_0996_),
    .A2(_0998_),
    .B1(_0995_),
    .Y(_1001_));
 sky130_fd_sc_hd__nor2_1 _6005_ (.A(_1000_),
    .B(_1001_),
    .Y(_1002_));
 sky130_fd_sc_hd__or3_1 _6006_ (.A(_4210_),
    .B(_0993_),
    .C(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__buf_2 _6007_ (.A(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__a22o_1 _6008_ (.A1(_0634_),
    .A2(_0994_),
    .B1(_0996_),
    .B2(_0997_),
    .X(_1005_));
 sky130_fd_sc_hd__or4_2 _6009_ (.A(_4017_),
    .B(_0802_),
    .C(_0773_),
    .D(_0992_),
    .X(_1006_));
 sky130_fd_sc_hd__inv_2 _6010_ (.A(_0802_),
    .Y(_1007_));
 sky130_fd_sc_hd__or3_2 _6011_ (.A(_4017_),
    .B(_0773_),
    .C(_0992_),
    .X(_1008_));
 sky130_fd_sc_hd__a21bo_1 _6012_ (.A1(_1007_),
    .A2(_0993_),
    .B1_N(_1008_),
    .X(_1010_));
 sky130_fd_sc_hd__nand4_1 _6013_ (.A(_0998_),
    .B(_1005_),
    .C(_1006_),
    .D(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__a22o_1 _6014_ (.A1(_0998_),
    .A2(_1005_),
    .B1(_1006_),
    .B2(_1010_),
    .X(_1012_));
 sky130_fd_sc_hd__nand2_1 _6015_ (.A(_1011_),
    .B(_1012_),
    .Y(_1013_));
 sky130_fd_sc_hd__and2_1 _6016_ (.A(_0998_),
    .B(_1005_),
    .X(_1014_));
 sky130_fd_sc_hd__clkbuf_2 _6017_ (.A(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__a21o_1 _6018_ (.A1(_0779_),
    .A2(_0803_),
    .B1(_0992_),
    .X(_1016_));
 sky130_fd_sc_hd__or3_2 _6019_ (.A(_0779_),
    .B(_0803_),
    .C(_0992_),
    .X(_1017_));
 sky130_fd_sc_hd__o21ai_1 _6020_ (.A1(_1008_),
    .A2(_1016_),
    .B1(_1017_),
    .Y(_1018_));
 sky130_fd_sc_hd__a31o_2 _6021_ (.A1(_3701_),
    .A2(_0737_),
    .A3(_0745_),
    .B1(_0754_),
    .X(_1019_));
 sky130_fd_sc_hd__nand2_1 _6022_ (.A(_1019_),
    .B(_0993_),
    .Y(_1020_));
 sky130_fd_sc_hd__o211a_1 _6023_ (.A1(_0803_),
    .A2(_0993_),
    .B1(_1008_),
    .C1(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__a21oi_1 _6024_ (.A1(_1006_),
    .A2(_1018_),
    .B1(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__nand2_1 _6025_ (.A(_1006_),
    .B(_1018_),
    .Y(_1023_));
 sky130_fd_sc_hd__a21bo_1 _6026_ (.A1(_1015_),
    .A2(_1022_),
    .B1_N(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__xnor2_1 _6027_ (.A(_1013_),
    .B(_1024_),
    .Y(_1025_));
 sky130_fd_sc_hd__xnor2_1 _6028_ (.A(_1004_),
    .B(_1025_),
    .Y(_1026_));
 sky130_fd_sc_hd__nor2_1 _6029_ (.A(_1015_),
    .B(_1022_),
    .Y(_1027_));
 sky130_fd_sc_hd__a21oi_1 _6030_ (.A1(_0779_),
    .A2(_0803_),
    .B1(_0992_),
    .Y(_1028_));
 sky130_fd_sc_hd__mux2_2 _6031_ (.A0(_1017_),
    .A1(_1028_),
    .S(_1008_),
    .X(_1029_));
 sky130_fd_sc_hd__nor2_2 _6032_ (.A(_0773_),
    .B(_1017_),
    .Y(_1031_));
 sky130_fd_sc_hd__a21o_1 _6033_ (.A1(_1015_),
    .A2(_1029_),
    .B1(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__nand2_1 _6034_ (.A(_1015_),
    .B(_1022_),
    .Y(_1033_));
 sky130_fd_sc_hd__a2bb2o_1 _6035_ (.A1_N(_1004_),
    .A2_N(_1027_),
    .B1(_1032_),
    .B2(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__and2_1 _6036_ (.A(_1026_),
    .B(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__xnor2_1 _6037_ (.A(_1026_),
    .B(_1034_),
    .Y(_1036_));
 sky130_fd_sc_hd__nor2_1 _6038_ (.A(_1000_),
    .B(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__a22oi_1 _6039_ (.A1(_0706_),
    .A2(_0993_),
    .B1(_0998_),
    .B2(_1005_),
    .Y(_1038_));
 sky130_fd_sc_hd__a21oi_1 _6040_ (.A1(_1006_),
    .A2(_1011_),
    .B1(_1038_),
    .Y(_1039_));
 sky130_fd_sc_hd__and2_1 _6041_ (.A(_1006_),
    .B(_1038_),
    .X(_1040_));
 sky130_fd_sc_hd__nor2_1 _6042_ (.A(_1039_),
    .B(_1040_),
    .Y(_1041_));
 sky130_fd_sc_hd__xnor2_1 _6043_ (.A(_1004_),
    .B(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__and3_1 _6044_ (.A(_1013_),
    .B(_1023_),
    .C(_1033_),
    .X(_1043_));
 sky130_fd_sc_hd__or2b_1 _6045_ (.A(_1013_),
    .B_N(_1024_),
    .X(_1044_));
 sky130_fd_sc_hd__o21a_1 _6046_ (.A1(_1004_),
    .A2(_1043_),
    .B1(_1044_),
    .X(_1045_));
 sky130_fd_sc_hd__xor2_1 _6047_ (.A(_1042_),
    .B(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__nor2_1 _6048_ (.A(_1000_),
    .B(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__and2_1 _6049_ (.A(_1000_),
    .B(_1046_),
    .X(_1048_));
 sky130_fd_sc_hd__nor2_1 _6050_ (.A(_1047_),
    .B(_1048_),
    .Y(_1049_));
 sky130_fd_sc_hd__o21ai_2 _6051_ (.A1(_1035_),
    .A2(_1037_),
    .B1(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__or2b_1 _6052_ (.A(_0978_),
    .B_N(_0971_),
    .X(_1052_));
 sky130_fd_sc_hd__o31a_1 _6053_ (.A1(_0962_),
    .A2(_0973_),
    .A3(_0979_),
    .B1(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__nor2_1 _6054_ (.A(_0971_),
    .B(_0972_),
    .Y(_1054_));
 sky130_fd_sc_hd__a21oi_1 _6055_ (.A1(_0943_),
    .A2(_0944_),
    .B1(_0959_),
    .Y(_1055_));
 sky130_fd_sc_hd__nor2_1 _6056_ (.A(_0960_),
    .B(_1055_),
    .Y(_1056_));
 sky130_fd_sc_hd__nand2_1 _6057_ (.A(_0949_),
    .B(_0958_),
    .Y(_1057_));
 sky130_fd_sc_hd__and3_1 _6058_ (.A(_0956_),
    .B(_0955_),
    .C(_0957_),
    .X(_1058_));
 sky130_fd_sc_hd__a21oi_1 _6059_ (.A1(_0956_),
    .A2(_0957_),
    .B1(_0955_),
    .Y(_1059_));
 sky130_fd_sc_hd__o21bai_1 _6060_ (.A1(_1058_),
    .A2(_1059_),
    .B1_N(_0949_),
    .Y(_1060_));
 sky130_fd_sc_hd__nor2_1 _6061_ (.A(_0951_),
    .B(_0954_),
    .Y(_1061_));
 sky130_fd_sc_hd__nor2_1 _6062_ (.A(_0955_),
    .B(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__or2_1 _6063_ (.A(_0945_),
    .B(_0947_),
    .X(_1063_));
 sky130_fd_sc_hd__and2_1 _6064_ (.A(_0952_),
    .B(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__and3_1 _6065_ (.A(_3892_),
    .B(_1019_),
    .C(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__and2_1 _6066_ (.A(_1062_),
    .B(_1065_),
    .X(_1066_));
 sky130_fd_sc_hd__a21o_1 _6067_ (.A1(_1057_),
    .A2(_1060_),
    .B1(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__or3b_1 _6068_ (.A(_0787_),
    .B(_3739_),
    .C_N(_0947_),
    .X(_1068_));
 sky130_fd_sc_hd__a21oi_1 _6069_ (.A1(_3892_),
    .A2(_1019_),
    .B1(_1064_),
    .Y(_1069_));
 sky130_fd_sc_hd__or2_1 _6070_ (.A(_1065_),
    .B(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__nor4_1 _6071_ (.A(_0955_),
    .B(_1061_),
    .C(_1068_),
    .D(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__and3_1 _6072_ (.A(_1057_),
    .B(_1060_),
    .C(_1066_),
    .X(_1073_));
 sky130_fd_sc_hd__a21o_1 _6073_ (.A1(_1067_),
    .A2(_1071_),
    .B1(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__and2_1 _6074_ (.A(_0942_),
    .B(_0960_),
    .X(_1075_));
 sky130_fd_sc_hd__a311o_1 _6075_ (.A1(_0942_),
    .A2(_1056_),
    .A3(_1074_),
    .B1(_0961_),
    .C1(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__nor2_1 _6076_ (.A(_0977_),
    .B(_0978_),
    .Y(_1077_));
 sky130_fd_sc_hd__a211o_1 _6077_ (.A1(_1054_),
    .A2(_1076_),
    .B1(_1077_),
    .C1(_0971_),
    .X(_1078_));
 sky130_fd_sc_hd__nand2_1 _6078_ (.A(_1056_),
    .B(_1074_),
    .Y(_1079_));
 sky130_fd_sc_hd__nor2_1 _6079_ (.A(_0961_),
    .B(_0960_),
    .Y(_1080_));
 sky130_fd_sc_hd__a211o_1 _6080_ (.A1(_0942_),
    .A2(_1080_),
    .B1(_1056_),
    .C1(_1074_),
    .X(_1081_));
 sky130_fd_sc_hd__and3b_1 _6081_ (.A_N(_1073_),
    .B(_1067_),
    .C(_1071_),
    .X(_1082_));
 sky130_fd_sc_hd__a21oi_1 _6082_ (.A1(_1057_),
    .A2(_1060_),
    .B1(_1066_),
    .Y(_1083_));
 sky130_fd_sc_hd__nor2_1 _6083_ (.A(_1062_),
    .B(_1065_),
    .Y(_1084_));
 sky130_fd_sc_hd__and2_1 _6084_ (.A(_1068_),
    .B(_1070_),
    .X(_1085_));
 sky130_fd_sc_hd__o221a_1 _6085_ (.A1(_1073_),
    .A2(_1083_),
    .B1(_1084_),
    .B2(_1066_),
    .C1(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__a21o_1 _6086_ (.A1(_3770_),
    .A2(_3739_),
    .B1(_0787_),
    .X(_1087_));
 sky130_fd_sc_hd__o221a_1 _6087_ (.A1(_0802_),
    .A2(_3739_),
    .B1(_1082_),
    .B2(_1086_),
    .C1(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__a21bo_1 _6088_ (.A1(_1079_),
    .A2(_1081_),
    .B1_N(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__xnor2_2 _6089_ (.A(_0973_),
    .B(_1076_),
    .Y(_1090_));
 sky130_fd_sc_hd__a211o_1 _6090_ (.A1(_1053_),
    .A2(_1078_),
    .B1(_1089_),
    .C1(_1090_),
    .X(_1091_));
 sky130_fd_sc_hd__xor2_2 _6091_ (.A(_0884_),
    .B(_0981_),
    .X(_1092_));
 sky130_fd_sc_hd__xnor2_1 _6092_ (.A(_1091_),
    .B(_1092_),
    .Y(_1094_));
 sky130_fd_sc_hd__buf_2 _6093_ (.A(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__and3_1 _6094_ (.A(_0762_),
    .B(_0722_),
    .C(_0994_),
    .X(_1096_));
 sky130_fd_sc_hd__buf_2 _6095_ (.A(_0634_),
    .X(_1097_));
 sky130_fd_sc_hd__a2111o_1 _6096_ (.A1(_1053_),
    .A2(_1078_),
    .B1(_1092_),
    .C1(_1090_),
    .D1(_1089_),
    .X(_1098_));
 sky130_fd_sc_hd__a21oi_1 _6097_ (.A1(_0884_),
    .A2(_0981_),
    .B1(_0987_),
    .Y(_1099_));
 sky130_fd_sc_hd__xnor2_2 _6098_ (.A(_1099_),
    .B(_0986_),
    .Y(_1100_));
 sky130_fd_sc_hd__a21oi_1 _6099_ (.A1(_1098_),
    .A2(_1100_),
    .B1(_4016_),
    .Y(_1101_));
 sky130_fd_sc_hd__buf_2 _6100_ (.A(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__and4_1 _6101_ (.A(_1097_),
    .B(_0996_),
    .C(_0997_),
    .D(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__or2_1 _6102_ (.A(_1096_),
    .B(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__nand2_1 _6103_ (.A(_0795_),
    .B(_1102_),
    .Y(_1105_));
 sky130_fd_sc_hd__xnor2_1 _6104_ (.A(_1104_),
    .B(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__xnor2_1 _6105_ (.A(_1095_),
    .B(_1106_),
    .Y(_1107_));
 sky130_fd_sc_hd__xnor2_1 _6106_ (.A(_1015_),
    .B(_1029_),
    .Y(_1108_));
 sky130_fd_sc_hd__a22o_1 _6107_ (.A1(_0996_),
    .A2(_0997_),
    .B1(_1102_),
    .B2(_1097_),
    .X(_1109_));
 sky130_fd_sc_hd__and2b_1 _6108_ (.A_N(_1103_),
    .B(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__a21oi_1 _6109_ (.A1(_1029_),
    .A2(_1110_),
    .B1(_1031_),
    .Y(_1111_));
 sky130_fd_sc_hd__nor2_1 _6110_ (.A(_1108_),
    .B(_1111_),
    .Y(_1112_));
 sky130_fd_sc_hd__nand2_1 _6111_ (.A(_1108_),
    .B(_1111_),
    .Y(_1113_));
 sky130_fd_sc_hd__or2b_1 _6112_ (.A(_1112_),
    .B_N(_1113_),
    .X(_1115_));
 sky130_fd_sc_hd__xor2_1 _6113_ (.A(_1107_),
    .B(_1115_),
    .X(_1116_));
 sky130_fd_sc_hd__a21o_1 _6114_ (.A1(_1008_),
    .A2(_1016_),
    .B1(_1031_),
    .X(_1117_));
 sky130_fd_sc_hd__or3_1 _6115_ (.A(_4017_),
    .B(_0892_),
    .C(_0992_),
    .X(_1118_));
 sky130_fd_sc_hd__a211o_1 _6116_ (.A1(_1098_),
    .A2(_1100_),
    .B1(_4017_),
    .C1(_0702_),
    .X(_1119_));
 sky130_fd_sc_hd__xnor2_1 _6117_ (.A(_1118_),
    .B(_1119_),
    .Y(_1120_));
 sky130_fd_sc_hd__or2b_1 _6118_ (.A(_1095_),
    .B_N(_1097_),
    .X(_1121_));
 sky130_fd_sc_hd__xnor2_1 _6119_ (.A(_1120_),
    .B(_1121_),
    .Y(_1122_));
 sky130_fd_sc_hd__o21ba_1 _6120_ (.A1(_1117_),
    .A2(_1122_),
    .B1_N(_1031_),
    .X(_1123_));
 sky130_fd_sc_hd__xnor2_1 _6121_ (.A(_1117_),
    .B(_1110_),
    .Y(_1124_));
 sky130_fd_sc_hd__or2b_1 _6122_ (.A(_1123_),
    .B_N(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__o211ai_1 _6123_ (.A1(_1090_),
    .A2(_1089_),
    .B1(_1078_),
    .C1(_1053_),
    .Y(_1126_));
 sky130_fd_sc_hd__and2_1 _6124_ (.A(_1091_),
    .B(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__buf_2 _6125_ (.A(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__o2bb2a_1 _6126_ (.A1_N(_1096_),
    .A2_N(_1102_),
    .B1(_1120_),
    .B2(_1121_),
    .X(_1129_));
 sky130_fd_sc_hd__nor2_1 _6127_ (.A(_0627_),
    .B(_1095_),
    .Y(_1130_));
 sky130_fd_sc_hd__xnor2_1 _6128_ (.A(_1129_),
    .B(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__xor2_1 _6129_ (.A(_1128_),
    .B(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__xnor2_1 _6130_ (.A(_1123_),
    .B(_1124_),
    .Y(_1133_));
 sky130_fd_sc_hd__nand2_1 _6131_ (.A(_1132_),
    .B(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__nand2_1 _6132_ (.A(_1125_),
    .B(_1134_),
    .Y(_1136_));
 sky130_fd_sc_hd__or2b_1 _6133_ (.A(_1116_),
    .B_N(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__xor2_1 _6134_ (.A(_1136_),
    .B(_1116_),
    .X(_1138_));
 sky130_fd_sc_hd__nand2_1 _6135_ (.A(_1128_),
    .B(_1131_),
    .Y(_1139_));
 sky130_fd_sc_hd__o31ai_2 _6136_ (.A1(_0627_),
    .A2(_1095_),
    .A3(_1129_),
    .B1(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__or2b_1 _6137_ (.A(_1138_),
    .B_N(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__and2b_1 _6138_ (.A_N(_1095_),
    .B(_1106_),
    .X(_1142_));
 sky130_fd_sc_hd__a31o_1 _6139_ (.A1(_0795_),
    .A2(_1102_),
    .A3(_1104_),
    .B1(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__xor2_1 _6140_ (.A(_1002_),
    .B(_1102_),
    .X(_1144_));
 sky130_fd_sc_hd__nand2_1 _6141_ (.A(_1015_),
    .B(_1031_),
    .Y(_1145_));
 sky130_fd_sc_hd__or3_1 _6142_ (.A(_1015_),
    .B(_1031_),
    .C(_1029_),
    .X(_1146_));
 sky130_fd_sc_hd__and2_1 _6143_ (.A(_1145_),
    .B(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__nand2_1 _6144_ (.A(_1144_),
    .B(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__or2_1 _6145_ (.A(_1144_),
    .B(_1147_),
    .X(_1149_));
 sky130_fd_sc_hd__and2_1 _6146_ (.A(_1148_),
    .B(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__a21o_1 _6147_ (.A1(_1107_),
    .A2(_1113_),
    .B1(_1112_),
    .X(_1151_));
 sky130_fd_sc_hd__xor2_1 _6148_ (.A(_1150_),
    .B(_1151_),
    .X(_1152_));
 sky130_fd_sc_hd__xnor2_1 _6149_ (.A(_1143_),
    .B(_1152_),
    .Y(_1153_));
 sky130_fd_sc_hd__a21oi_1 _6150_ (.A1(_1137_),
    .A2(_1141_),
    .B1(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__and3_1 _6151_ (.A(_1137_),
    .B(_1141_),
    .C(_1153_),
    .X(_1155_));
 sky130_fd_sc_hd__or2_1 _6152_ (.A(_1154_),
    .B(_1155_),
    .X(_1157_));
 sky130_fd_sc_hd__xor2_1 _6153_ (.A(_1140_),
    .B(_1138_),
    .X(_1158_));
 sky130_fd_sc_hd__or3_1 _6154_ (.A(_0892_),
    .B(_1095_),
    .C(_1119_),
    .X(_1159_));
 sky130_fd_sc_hd__a2bb2o_1 _6155_ (.A1_N(_0702_),
    .A2_N(_1095_),
    .B1(_1102_),
    .B2(_0762_),
    .X(_1160_));
 sky130_fd_sc_hd__and2_1 _6156_ (.A(_1097_),
    .B(_1128_),
    .X(_1161_));
 sky130_fd_sc_hd__nand3_1 _6157_ (.A(_1160_),
    .B(_1159_),
    .C(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__nand2_1 _6158_ (.A(_1159_),
    .B(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__clkbuf_4 _6159_ (.A(_1089_),
    .X(_1164_));
 sky130_fd_sc_hd__nor2_1 _6160_ (.A(_1090_),
    .B(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__and2_1 _6161_ (.A(_1090_),
    .B(_1089_),
    .X(_1166_));
 sky130_fd_sc_hd__or2_1 _6162_ (.A(_1165_),
    .B(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__buf_2 _6163_ (.A(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__nand2_1 _6164_ (.A(_0795_),
    .B(_1128_),
    .Y(_1169_));
 sky130_fd_sc_hd__xnor2_1 _6165_ (.A(_1163_),
    .B(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__and2b_1 _6166_ (.A_N(_1168_),
    .B(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__a31o_1 _6167_ (.A1(_0795_),
    .A2(_1128_),
    .A3(_1163_),
    .B1(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__xnor2_1 _6168_ (.A(_1168_),
    .B(_1170_),
    .Y(_1173_));
 sky130_fd_sc_hd__a21o_1 _6169_ (.A1(_1160_),
    .A2(_1159_),
    .B1(_1161_),
    .X(_1174_));
 sky130_fd_sc_hd__or3b_1 _6170_ (.A(_1016_),
    .B(_1008_),
    .C_N(_1017_),
    .X(_1175_));
 sky130_fd_sc_hd__and4_1 _6171_ (.A(_0706_),
    .B(_1017_),
    .C(_1028_),
    .D(_1101_),
    .X(_1176_));
 sky130_fd_sc_hd__a21o_1 _6172_ (.A1(_1175_),
    .A2(_1029_),
    .B1(_1176_),
    .X(_1178_));
 sky130_fd_sc_hd__and3_1 _6173_ (.A(_1162_),
    .B(_1174_),
    .C(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__nor2_1 _6174_ (.A(_1031_),
    .B(_1179_),
    .Y(_1180_));
 sky130_fd_sc_hd__xnor2_1 _6175_ (.A(_1029_),
    .B(_1122_),
    .Y(_1181_));
 sky130_fd_sc_hd__xnor2_1 _6176_ (.A(_1180_),
    .B(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__and2b_1 _6177_ (.A_N(_1180_),
    .B(_1181_),
    .X(_1183_));
 sky130_fd_sc_hd__a21oi_1 _6178_ (.A1(_1173_),
    .A2(_1182_),
    .B1(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__or2_1 _6179_ (.A(_1132_),
    .B(_1133_),
    .X(_1185_));
 sky130_fd_sc_hd__nand2_1 _6180_ (.A(_1134_),
    .B(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__xor2_1 _6181_ (.A(_1184_),
    .B(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__nor2_1 _6182_ (.A(_1184_),
    .B(_1186_),
    .Y(_1189_));
 sky130_fd_sc_hd__a21oi_1 _6183_ (.A1(_1172_),
    .A2(_1187_),
    .B1(_1189_),
    .Y(_1190_));
 sky130_fd_sc_hd__xnor2_1 _6184_ (.A(_1158_),
    .B(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__or2_1 _6185_ (.A(_0892_),
    .B(_1094_),
    .X(_1192_));
 sky130_fd_sc_hd__nand2_1 _6186_ (.A(_0722_),
    .B(_1127_),
    .Y(_1193_));
 sky130_fd_sc_hd__xnor2_1 _6187_ (.A(_1192_),
    .B(_1193_),
    .Y(_1194_));
 sky130_fd_sc_hd__or2b_1 _6188_ (.A(_1168_),
    .B_N(_1097_),
    .X(_1195_));
 sky130_fd_sc_hd__xor2_1 _6189_ (.A(_1194_),
    .B(_1195_),
    .X(_1196_));
 sky130_fd_sc_hd__nor2_1 _6190_ (.A(_0773_),
    .B(_1095_),
    .Y(_1197_));
 sky130_fd_sc_hd__nor2_1 _6191_ (.A(_0779_),
    .B(_0992_),
    .Y(_1198_));
 sky130_fd_sc_hd__a211o_1 _6192_ (.A1(_1098_),
    .A2(_1100_),
    .B1(_4016_),
    .C1(_0802_),
    .X(_1200_));
 sky130_fd_sc_hd__xnor2_1 _6193_ (.A(_1198_),
    .B(_1200_),
    .Y(_1201_));
 sky130_fd_sc_hd__and3_1 _6194_ (.A(_1007_),
    .B(_1198_),
    .C(_1101_),
    .X(_1202_));
 sky130_fd_sc_hd__a21o_1 _6195_ (.A1(_1197_),
    .A2(_1201_),
    .B1(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__a22o_1 _6196_ (.A1(_1017_),
    .A2(_1028_),
    .B1(_1102_),
    .B2(_0706_),
    .X(_1204_));
 sky130_fd_sc_hd__and2b_1 _6197_ (.A_N(_1176_),
    .B(_1204_),
    .X(_1205_));
 sky130_fd_sc_hd__xor2_1 _6198_ (.A(_1203_),
    .B(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__and2_1 _6199_ (.A(_1203_),
    .B(_1205_),
    .X(_1207_));
 sky130_fd_sc_hd__a21oi_1 _6200_ (.A1(_1196_),
    .A2(_1206_),
    .B1(_1207_),
    .Y(_1208_));
 sky130_fd_sc_hd__a21oi_1 _6201_ (.A1(_1162_),
    .A2(_1174_),
    .B1(_1178_),
    .Y(_1209_));
 sky130_fd_sc_hd__nor2_1 _6202_ (.A(_1179_),
    .B(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__xnor2_1 _6203_ (.A(_1208_),
    .B(_1210_),
    .Y(_1211_));
 sky130_fd_sc_hd__or2_1 _6204_ (.A(_1192_),
    .B(_1193_),
    .X(_1212_));
 sky130_fd_sc_hd__o21a_1 _6205_ (.A1(_1194_),
    .A2(_1195_),
    .B1(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__or2_1 _6206_ (.A(_0627_),
    .B(_1168_),
    .X(_1214_));
 sky130_fd_sc_hd__xor2_1 _6207_ (.A(_1213_),
    .B(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__xor2_1 _6208_ (.A(_1164_),
    .B(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__and2b_1 _6209_ (.A_N(_1208_),
    .B(_1210_),
    .X(_1217_));
 sky130_fd_sc_hd__a21o_1 _6210_ (.A1(_1211_),
    .A2(_1216_),
    .B1(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__xor2_1 _6211_ (.A(_1173_),
    .B(_1182_),
    .X(_1219_));
 sky130_fd_sc_hd__nand2_1 _6212_ (.A(_1218_),
    .B(_1219_),
    .Y(_1221_));
 sky130_fd_sc_hd__xnor2_1 _6213_ (.A(_1218_),
    .B(_1219_),
    .Y(_1222_));
 sky130_fd_sc_hd__a2bb2o_1 _6214_ (.A1_N(_1213_),
    .A2_N(_1214_),
    .B1(_1215_),
    .B2(_1164_),
    .X(_1223_));
 sky130_fd_sc_hd__or2b_1 _6215_ (.A(_1222_),
    .B_N(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__xnor2_1 _6216_ (.A(_1172_),
    .B(_1187_),
    .Y(_1225_));
 sky130_fd_sc_hd__and3_1 _6217_ (.A(_1221_),
    .B(_1224_),
    .C(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__xor2_1 _6218_ (.A(_1223_),
    .B(_1222_),
    .X(_1227_));
 sky130_fd_sc_hd__or2_1 _6219_ (.A(_0892_),
    .B(_1168_),
    .X(_1228_));
 sky130_fd_sc_hd__nand2_1 _6220_ (.A(_0762_),
    .B(_1128_),
    .Y(_1229_));
 sky130_fd_sc_hd__nor2_1 _6221_ (.A(_0702_),
    .B(_1168_),
    .Y(_1230_));
 sky130_fd_sc_hd__xor2_1 _6222_ (.A(_1229_),
    .B(_1230_),
    .X(_1232_));
 sky130_fd_sc_hd__nand2_1 _6223_ (.A(_1097_),
    .B(_1164_),
    .Y(_1233_));
 sky130_fd_sc_hd__o22ai_1 _6224_ (.A1(_1193_),
    .A2(_1228_),
    .B1(_1232_),
    .B2(_1233_),
    .Y(_1234_));
 sky130_fd_sc_hd__and3_1 _6225_ (.A(_0795_),
    .B(_1164_),
    .C(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__a21oi_1 _6226_ (.A1(_0795_),
    .A2(_1164_),
    .B1(_1234_),
    .Y(_1236_));
 sky130_fd_sc_hd__nor2_1 _6227_ (.A(_1235_),
    .B(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__xnor2_1 _6228_ (.A(_1232_),
    .B(_1233_),
    .Y(_1238_));
 sky130_fd_sc_hd__and2_1 _6229_ (.A(_0706_),
    .B(_1127_),
    .X(_1239_));
 sky130_fd_sc_hd__a2bb2o_1 _6230_ (.A1_N(_0802_),
    .A2_N(_1095_),
    .B1(_1019_),
    .B2(_1102_),
    .X(_1240_));
 sky130_fd_sc_hd__or4b_1 _6231_ (.A(_0802_),
    .B(_1094_),
    .C(_0787_),
    .D_N(_1101_),
    .X(_1241_));
 sky130_fd_sc_hd__a21bo_1 _6232_ (.A1(_1239_),
    .A2(_1240_),
    .B1_N(_1241_),
    .X(_1243_));
 sky130_fd_sc_hd__xnor2_1 _6233_ (.A(_1197_),
    .B(_1201_),
    .Y(_1244_));
 sky130_fd_sc_hd__xor2_1 _6234_ (.A(_1243_),
    .B(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__or2b_1 _6235_ (.A(_1244_),
    .B_N(_1243_),
    .X(_1246_));
 sky130_fd_sc_hd__o21ai_1 _6236_ (.A1(_1238_),
    .A2(_1245_),
    .B1(_1246_),
    .Y(_1247_));
 sky130_fd_sc_hd__xor2_1 _6237_ (.A(_1196_),
    .B(_1206_),
    .X(_1248_));
 sky130_fd_sc_hd__xor2_1 _6238_ (.A(_1247_),
    .B(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__nand2_1 _6239_ (.A(_1247_),
    .B(_1248_),
    .Y(_1250_));
 sky130_fd_sc_hd__a21boi_1 _6240_ (.A1(_1237_),
    .A2(_1249_),
    .B1_N(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__xnor2_1 _6241_ (.A(_1211_),
    .B(_1216_),
    .Y(_1252_));
 sky130_fd_sc_hd__xor2_1 _6242_ (.A(_1251_),
    .B(_1252_),
    .X(_1254_));
 sky130_fd_sc_hd__nor2_1 _6243_ (.A(_1251_),
    .B(_1252_),
    .Y(_1255_));
 sky130_fd_sc_hd__a21oi_1 _6244_ (.A1(_1235_),
    .A2(_1254_),
    .B1(_1255_),
    .Y(_1256_));
 sky130_fd_sc_hd__xnor2_1 _6245_ (.A(_1227_),
    .B(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__xnor2_1 _6246_ (.A(_1237_),
    .B(_1249_),
    .Y(_1258_));
 sky130_fd_sc_hd__nand2_1 _6247_ (.A(_0722_),
    .B(_1164_),
    .Y(_1259_));
 sky130_fd_sc_hd__nor2_1 _6248_ (.A(_1228_),
    .B(_1259_),
    .Y(_1260_));
 sky130_fd_sc_hd__xor2_1 _6249_ (.A(_1238_),
    .B(_1245_),
    .X(_1261_));
 sky130_fd_sc_hd__xor2_1 _6250_ (.A(_1228_),
    .B(_1259_),
    .X(_1262_));
 sky130_fd_sc_hd__nand3_1 _6251_ (.A(_1241_),
    .B(_1239_),
    .C(_1240_),
    .Y(_1263_));
 sky130_fd_sc_hd__a21o_1 _6252_ (.A1(_1241_),
    .A2(_1240_),
    .B1(_1239_),
    .X(_1265_));
 sky130_fd_sc_hd__nor2_1 _6253_ (.A(_0773_),
    .B(_1168_),
    .Y(_1266_));
 sky130_fd_sc_hd__a2bb2o_1 _6254_ (.A1_N(_0787_),
    .A2_N(_1095_),
    .B1(_1128_),
    .B2(_1007_),
    .X(_1267_));
 sky130_fd_sc_hd__or4b_1 _6255_ (.A(_0802_),
    .B(_0787_),
    .C(_1094_),
    .D_N(_1127_),
    .X(_1268_));
 sky130_fd_sc_hd__a21bo_1 _6256_ (.A1(_1266_),
    .A2(_1267_),
    .B1_N(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__a21o_1 _6257_ (.A1(_1263_),
    .A2(_1265_),
    .B1(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__and3_1 _6258_ (.A(_1263_),
    .B(_1265_),
    .C(_1269_),
    .X(_1271_));
 sky130_fd_sc_hd__a21oi_1 _6259_ (.A1(_1262_),
    .A2(_1270_),
    .B1(_1271_),
    .Y(_1272_));
 sky130_fd_sc_hd__xnor2_1 _6260_ (.A(_1261_),
    .B(_1272_),
    .Y(_1273_));
 sky130_fd_sc_hd__and2b_1 _6261_ (.A_N(_1272_),
    .B(_1261_),
    .X(_1274_));
 sky130_fd_sc_hd__a21oi_1 _6262_ (.A1(_1260_),
    .A2(_1273_),
    .B1(_1274_),
    .Y(_1276_));
 sky130_fd_sc_hd__or2_1 _6263_ (.A(_1258_),
    .B(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__xnor2_1 _6264_ (.A(_1258_),
    .B(_1276_),
    .Y(_1278_));
 sky130_fd_sc_hd__and3_1 _6265_ (.A(_1268_),
    .B(_1266_),
    .C(_1267_),
    .X(_1279_));
 sky130_fd_sc_hd__a21oi_1 _6266_ (.A1(_1268_),
    .A2(_1267_),
    .B1(_1266_),
    .Y(_1280_));
 sky130_fd_sc_hd__nor2_1 _6267_ (.A(_1279_),
    .B(_1280_),
    .Y(_1281_));
 sky130_fd_sc_hd__nor2_1 _6268_ (.A(_0802_),
    .B(_1168_),
    .Y(_1282_));
 sky130_fd_sc_hd__a21o_1 _6269_ (.A1(_1019_),
    .A2(_1128_),
    .B1(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__and3_1 _6270_ (.A(_1019_),
    .B(_1128_),
    .C(_1282_),
    .X(_1284_));
 sky130_fd_sc_hd__a31o_1 _6271_ (.A1(_0706_),
    .A2(_1164_),
    .A3(_1283_),
    .B1(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__nand2_1 _6272_ (.A(_1281_),
    .B(_1285_),
    .Y(_1287_));
 sky130_fd_sc_hd__and2_1 _6273_ (.A(_0762_),
    .B(_1164_),
    .X(_1288_));
 sky130_fd_sc_hd__xor2_1 _6274_ (.A(_1281_),
    .B(_1285_),
    .X(_1289_));
 sky130_fd_sc_hd__nand2_1 _6275_ (.A(_1288_),
    .B(_1289_),
    .Y(_1290_));
 sky130_fd_sc_hd__nor2_1 _6276_ (.A(_0706_),
    .B(_1128_),
    .Y(_1291_));
 sky130_fd_sc_hd__o2111a_1 _6277_ (.A1(_1239_),
    .A2(_1291_),
    .B1(_1282_),
    .C1(_1019_),
    .D1(_1164_),
    .X(_1292_));
 sky130_fd_sc_hd__o21ai_1 _6278_ (.A1(_1288_),
    .A2(_1289_),
    .B1(_1292_),
    .Y(_1293_));
 sky130_fd_sc_hd__and2b_1 _6279_ (.A_N(_1271_),
    .B(_1270_),
    .X(_1294_));
 sky130_fd_sc_hd__xnor2_1 _6280_ (.A(_1262_),
    .B(_1294_),
    .Y(_1295_));
 sky130_fd_sc_hd__o21a_1 _6281_ (.A1(_1287_),
    .A2(_1293_),
    .B1(_1295_),
    .X(_1296_));
 sky130_fd_sc_hd__a31o_1 _6282_ (.A1(_1287_),
    .A2(_1290_),
    .A3(_1293_),
    .B1(_1296_),
    .X(_1298_));
 sky130_fd_sc_hd__xnor2_1 _6283_ (.A(_1260_),
    .B(_1273_),
    .Y(_1299_));
 sky130_fd_sc_hd__or3_2 _6284_ (.A(_1278_),
    .B(_1298_),
    .C(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__xnor2_1 _6285_ (.A(_1235_),
    .B(_1254_),
    .Y(_1301_));
 sky130_fd_sc_hd__a21o_1 _6286_ (.A1(_1277_),
    .A2(_1300_),
    .B1(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__a21o_1 _6287_ (.A1(_1221_),
    .A2(_1224_),
    .B1(_1225_),
    .X(_1303_));
 sky130_fd_sc_hd__or2_1 _6288_ (.A(_1227_),
    .B(_1256_),
    .X(_1304_));
 sky130_fd_sc_hd__o211a_1 _6289_ (.A1(_1257_),
    .A2(_1302_),
    .B1(_1303_),
    .C1(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__or4_2 _6290_ (.A(_1157_),
    .B(_1191_),
    .C(_1226_),
    .D(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__inv_2 _6291_ (.A(_1154_),
    .Y(_1307_));
 sky130_fd_sc_hd__or2_1 _6292_ (.A(_1158_),
    .B(_1190_),
    .X(_1309_));
 sky130_fd_sc_hd__a21o_1 _6293_ (.A1(_1307_),
    .A2(_1309_),
    .B1(_1155_),
    .X(_1310_));
 sky130_fd_sc_hd__and2_1 _6294_ (.A(_1000_),
    .B(_1036_),
    .X(_1311_));
 sky130_fd_sc_hd__nor2_1 _6295_ (.A(_1037_),
    .B(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__a21o_1 _6296_ (.A1(_1033_),
    .A2(_1032_),
    .B1(_1027_),
    .X(_1313_));
 sky130_fd_sc_hd__xnor2_1 _6297_ (.A(_1004_),
    .B(_1313_),
    .Y(_1314_));
 sky130_fd_sc_hd__a21oi_1 _6298_ (.A1(_1145_),
    .A2(_1148_),
    .B1(_1314_),
    .Y(_1315_));
 sky130_fd_sc_hd__a21o_1 _6299_ (.A1(_1002_),
    .A2(_1102_),
    .B1(_1001_),
    .X(_1316_));
 sky130_fd_sc_hd__and3_1 _6300_ (.A(_1145_),
    .B(_1148_),
    .C(_1314_),
    .X(_1317_));
 sky130_fd_sc_hd__nor2_1 _6301_ (.A(_1315_),
    .B(_1317_),
    .Y(_1318_));
 sky130_fd_sc_hd__and2_1 _6302_ (.A(_1316_),
    .B(_1318_),
    .X(_1320_));
 sky130_fd_sc_hd__nor3_1 _6303_ (.A(_1312_),
    .B(_1315_),
    .C(_1320_),
    .Y(_1321_));
 sky130_fd_sc_hd__o21ai_1 _6304_ (.A1(_1315_),
    .A2(_1320_),
    .B1(_1312_),
    .Y(_1322_));
 sky130_fd_sc_hd__or2b_1 _6305_ (.A(_1321_),
    .B_N(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__xnor2_1 _6306_ (.A(_1316_),
    .B(_1318_),
    .Y(_1324_));
 sky130_fd_sc_hd__nand2_1 _6307_ (.A(_1150_),
    .B(_1151_),
    .Y(_1325_));
 sky130_fd_sc_hd__a21boi_1 _6308_ (.A1(_1143_),
    .A2(_1152_),
    .B1_N(_1325_),
    .Y(_1326_));
 sky130_fd_sc_hd__nor2_2 _6309_ (.A(_1324_),
    .B(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__and2_1 _6310_ (.A(_1324_),
    .B(_1326_),
    .X(_1328_));
 sky130_fd_sc_hd__or2_1 _6311_ (.A(_1327_),
    .B(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__a211o_1 _6312_ (.A1(_1306_),
    .A2(_1310_),
    .B1(_1323_),
    .C1(_1329_),
    .X(_1331_));
 sky130_fd_sc_hd__inv_2 _6313_ (.A(_1322_),
    .Y(_1332_));
 sky130_fd_sc_hd__o21bai_1 _6314_ (.A1(_1332_),
    .A2(_1327_),
    .B1_N(_1321_),
    .Y(_1333_));
 sky130_fd_sc_hd__or3_1 _6315_ (.A(_1049_),
    .B(_1035_),
    .C(_1037_),
    .X(_1334_));
 sky130_fd_sc_hd__nand2_1 _6316_ (.A(_1050_),
    .B(_1334_),
    .Y(_1335_));
 sky130_fd_sc_hd__a21o_1 _6317_ (.A1(_1331_),
    .A2(_1333_),
    .B1(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__and2b_1 _6318_ (.A_N(_1045_),
    .B(_1042_),
    .X(_1337_));
 sky130_fd_sc_hd__or4b_2 _6319_ (.A(_4210_),
    .B(_0702_),
    .C(_0993_),
    .D_N(_1097_),
    .X(_1338_));
 sky130_fd_sc_hd__a22o_1 _6320_ (.A1(_0762_),
    .A2(_0993_),
    .B1(_0994_),
    .B2(_0722_),
    .X(_1339_));
 sky130_fd_sc_hd__a21o_1 _6321_ (.A1(_1097_),
    .A2(_0994_),
    .B1(_1339_),
    .X(_1340_));
 sky130_fd_sc_hd__nand2_1 _6322_ (.A(_1338_),
    .B(_1340_),
    .Y(_1342_));
 sky130_fd_sc_hd__xor2_1 _6323_ (.A(_1004_),
    .B(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__o21ba_1 _6324_ (.A1(_1004_),
    .A2(_1040_),
    .B1_N(_1039_),
    .X(_1344_));
 sky130_fd_sc_hd__xnor2_1 _6325_ (.A(_1343_),
    .B(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__and2b_1 _6326_ (.A_N(_1000_),
    .B(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__and2b_1 _6327_ (.A_N(_1345_),
    .B(_1000_),
    .X(_1347_));
 sky130_fd_sc_hd__nor2_1 _6328_ (.A(_1346_),
    .B(_1347_),
    .Y(_1348_));
 sky130_fd_sc_hd__o21a_1 _6329_ (.A1(_1337_),
    .A2(_1047_),
    .B1(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__nor3_1 _6330_ (.A(_1348_),
    .B(_1337_),
    .C(_1047_),
    .Y(_1350_));
 sky130_fd_sc_hd__or2_1 _6331_ (.A(_1349_),
    .B(_1350_),
    .X(_1351_));
 sky130_fd_sc_hd__a21o_2 _6332_ (.A1(_1050_),
    .A2(_1336_),
    .B1(_1351_),
    .X(_1353_));
 sky130_fd_sc_hd__nand3_4 _6333_ (.A(_1351_),
    .B(_1050_),
    .C(_1336_),
    .Y(_1354_));
 sky130_fd_sc_hd__inv_2 _6334_ (.A(_4037_),
    .Y(_1355_));
 sky130_fd_sc_hd__and3_1 _6335_ (.A(_1353_),
    .B(_1354_),
    .C(_1355_),
    .X(_1356_));
 sky130_fd_sc_hd__and2b_1 _6336_ (.A_N(_1344_),
    .B(_1343_),
    .X(_1357_));
 sky130_fd_sc_hd__or2_1 _6337_ (.A(_1004_),
    .B(_1342_),
    .X(_1358_));
 sky130_fd_sc_hd__a22o_1 _6338_ (.A1(_0722_),
    .A2(_0993_),
    .B1(_0994_),
    .B2(_1097_),
    .X(_1359_));
 sky130_fd_sc_hd__nand2_1 _6339_ (.A(_0627_),
    .B(_1338_),
    .Y(_1360_));
 sky130_fd_sc_hd__o21ai_1 _6340_ (.A1(_0995_),
    .A2(_1338_),
    .B1(_1360_),
    .Y(_1361_));
 sky130_fd_sc_hd__nand2_1 _6341_ (.A(_0994_),
    .B(_1361_),
    .Y(_1362_));
 sky130_fd_sc_hd__xor2_1 _6342_ (.A(_1359_),
    .B(_1362_),
    .X(_1364_));
 sky130_fd_sc_hd__or2_1 _6343_ (.A(_1358_),
    .B(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__nand2_1 _6344_ (.A(_1358_),
    .B(_1364_),
    .Y(_1366_));
 sky130_fd_sc_hd__nand2_1 _6345_ (.A(_1365_),
    .B(_1366_),
    .Y(_1367_));
 sky130_fd_sc_hd__or2_1 _6346_ (.A(_1000_),
    .B(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__nand2_1 _6347_ (.A(_1000_),
    .B(_1367_),
    .Y(_1369_));
 sky130_fd_sc_hd__and2_1 _6348_ (.A(_1368_),
    .B(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__o21ai_1 _6349_ (.A1(_1357_),
    .A2(_1346_),
    .B1(_1370_),
    .Y(_1371_));
 sky130_fd_sc_hd__or3_1 _6350_ (.A(_1370_),
    .B(_1357_),
    .C(_1346_),
    .X(_1372_));
 sky130_fd_sc_hd__nand2_1 _6351_ (.A(_1371_),
    .B(_1372_),
    .Y(_1373_));
 sky130_fd_sc_hd__inv_2 _6352_ (.A(_1373_),
    .Y(_1375_));
 sky130_fd_sc_hd__or2_1 _6353_ (.A(_1323_),
    .B(_1329_),
    .X(_1376_));
 sky130_fd_sc_hd__or2_1 _6354_ (.A(_1351_),
    .B(_1335_),
    .X(_1377_));
 sky130_fd_sc_hd__a211o_1 _6355_ (.A1(_1306_),
    .A2(_1310_),
    .B1(_1376_),
    .C1(_1377_),
    .X(_1378_));
 sky130_fd_sc_hd__inv_2 _6356_ (.A(_1349_),
    .Y(_1379_));
 sky130_fd_sc_hd__o221a_1 _6357_ (.A1(_1350_),
    .A2(_1050_),
    .B1(_1377_),
    .B2(_1333_),
    .C1(_1379_),
    .X(_1380_));
 sky130_fd_sc_hd__nand2_1 _6358_ (.A(_1378_),
    .B(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__xnor2_1 _6359_ (.A(_1375_),
    .B(_1381_),
    .Y(_1382_));
 sky130_fd_sc_hd__buf_2 _6360_ (.A(_1382_),
    .X(_1383_));
 sky130_fd_sc_hd__buf_4 _6361_ (.A(_3615_),
    .X(_1384_));
 sky130_fd_sc_hd__nor2_2 _6362_ (.A(_1383_),
    .B(_1384_),
    .Y(_1386_));
 sky130_fd_sc_hd__or2b_1 _6363_ (.A(_1362_),
    .B_N(_1359_),
    .X(_1387_));
 sky130_fd_sc_hd__and2_1 _6364_ (.A(_0627_),
    .B(_0994_),
    .X(_1388_));
 sky130_fd_sc_hd__a21o_1 _6365_ (.A1(_1097_),
    .A2(_0993_),
    .B1(_1388_),
    .X(_1389_));
 sky130_fd_sc_hd__inv_2 _6366_ (.A(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__xnor2_1 _6367_ (.A(_1387_),
    .B(_1390_),
    .Y(_1391_));
 sky130_fd_sc_hd__inv_2 _6368_ (.A(_1338_),
    .Y(_1392_));
 sky130_fd_sc_hd__a21o_1 _6369_ (.A1(_0995_),
    .A2(_1391_),
    .B1(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__and3_1 _6370_ (.A(_1365_),
    .B(_1368_),
    .C(_1393_),
    .X(_1394_));
 sky130_fd_sc_hd__a21oi_1 _6371_ (.A1(_1365_),
    .A2(_1368_),
    .B1(_1393_),
    .Y(_1395_));
 sky130_fd_sc_hd__or2_2 _6372_ (.A(_1394_),
    .B(_1395_),
    .X(_1397_));
 sky130_fd_sc_hd__a21bo_1 _6373_ (.A1(_1375_),
    .A2(_1381_),
    .B1_N(_1371_),
    .X(_1398_));
 sky130_fd_sc_hd__xor2_4 _6374_ (.A(_1397_),
    .B(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__clkbuf_4 _6375_ (.A(_1399_),
    .X(_1400_));
 sky130_fd_sc_hd__clkbuf_4 _6376_ (.A(_3817_),
    .X(_1401_));
 sky130_fd_sc_hd__nor2_1 _6377_ (.A(_1400_),
    .B(_1401_),
    .Y(_1402_));
 sky130_fd_sc_hd__xor2_1 _6378_ (.A(_1356_),
    .B(_1386_),
    .X(_1403_));
 sky130_fd_sc_hd__a22o_1 _6379_ (.A1(_1356_),
    .A2(_1386_),
    .B1(_1402_),
    .B2(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__a21oi_2 _6380_ (.A1(_1306_),
    .A2(_1310_),
    .B1(_1329_),
    .Y(_1405_));
 sky130_fd_sc_hd__inv_2 _6381_ (.A(_1323_),
    .Y(_1406_));
 sky130_fd_sc_hd__o21ai_4 _6382_ (.A1(_1327_),
    .A2(_1405_),
    .B1(_1406_),
    .Y(_1408_));
 sky130_fd_sc_hd__or3_4 _6383_ (.A(_1406_),
    .B(_1327_),
    .C(_1405_),
    .X(_1409_));
 sky130_fd_sc_hd__nand2_2 _6384_ (.A(_1408_),
    .B(_1409_),
    .Y(_1410_));
 sky130_fd_sc_hd__or2_1 _6385_ (.A(_4228_),
    .B(_1410_),
    .X(_1411_));
 sky130_fd_sc_hd__and3_1 _6386_ (.A(_1329_),
    .B(_1306_),
    .C(_1310_),
    .X(_1412_));
 sky130_fd_sc_hd__nor2_1 _6387_ (.A(_1405_),
    .B(_1412_),
    .Y(_1413_));
 sky130_fd_sc_hd__clkbuf_4 _6388_ (.A(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__nand2_1 _6389_ (.A(_4217_),
    .B(_1414_),
    .Y(_1415_));
 sky130_fd_sc_hd__nand2_2 _6390_ (.A(_0218_),
    .B(_1414_),
    .Y(_1416_));
 sky130_fd_sc_hd__or2_1 _6391_ (.A(_0303_),
    .B(_1410_),
    .X(_1417_));
 sky130_fd_sc_hd__and2_1 _6392_ (.A(_1416_),
    .B(_1417_),
    .X(_1419_));
 sky130_fd_sc_hd__buf_2 _6393_ (.A(_3840_),
    .X(_1420_));
 sky130_fd_sc_hd__nand2_1 _6394_ (.A(_1331_),
    .B(_1333_),
    .Y(_1421_));
 sky130_fd_sc_hd__xor2_2 _6395_ (.A(_1335_),
    .B(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__clkbuf_4 _6396_ (.A(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__or2_2 _6397_ (.A(_1420_),
    .B(_1423_),
    .X(_1424_));
 sky130_fd_sc_hd__o22a_1 _6398_ (.A1(_1411_),
    .A2(_1415_),
    .B1(_1419_),
    .B2(_1424_),
    .X(_1425_));
 sky130_fd_sc_hd__nor2_1 _6399_ (.A(_1400_),
    .B(_1384_),
    .Y(_1426_));
 sky130_fd_sc_hd__and3_1 _6400_ (.A(_1353_),
    .B(_1354_),
    .C(_4153_),
    .X(_1427_));
 sky130_fd_sc_hd__buf_4 _6401_ (.A(_4037_),
    .X(_1428_));
 sky130_fd_sc_hd__nor2_1 _6402_ (.A(_1383_),
    .B(_1428_),
    .Y(_1430_));
 sky130_fd_sc_hd__xor2_1 _6403_ (.A(_1427_),
    .B(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__xor2_1 _6404_ (.A(_1426_),
    .B(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__xnor2_1 _6405_ (.A(_1425_),
    .B(_1432_),
    .Y(_1433_));
 sky130_fd_sc_hd__and2b_1 _6406_ (.A_N(_1425_),
    .B(_1432_),
    .X(_1434_));
 sky130_fd_sc_hd__a21o_1 _6407_ (.A1(_1404_),
    .A2(_1433_),
    .B1(_1434_),
    .X(_1435_));
 sky130_fd_sc_hd__inv_2 _6408_ (.A(_1395_),
    .Y(_1436_));
 sky130_fd_sc_hd__a21o_1 _6409_ (.A1(_1371_),
    .A2(_1436_),
    .B1(_1394_),
    .X(_1437_));
 sky130_fd_sc_hd__a211o_1 _6410_ (.A1(_1378_),
    .A2(_1380_),
    .B1(_1397_),
    .C1(_1373_),
    .X(_1438_));
 sky130_fd_sc_hd__a21o_1 _6411_ (.A1(_0795_),
    .A2(_0993_),
    .B1(_1388_),
    .X(_1439_));
 sky130_fd_sc_hd__o211a_1 _6412_ (.A1(_1387_),
    .A2(_1390_),
    .B1(_1439_),
    .C1(_1338_),
    .X(_1441_));
 sky130_fd_sc_hd__a21o_1 _6413_ (.A1(_0795_),
    .A2(_1392_),
    .B1(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__and3_1 _6414_ (.A(_1437_),
    .B(_1438_),
    .C(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__a21oi_1 _6415_ (.A1(_1437_),
    .A2(_1438_),
    .B1(_1442_),
    .Y(_1444_));
 sky130_fd_sc_hd__nor2_1 _6416_ (.A(_1443_),
    .B(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__buf_2 _6417_ (.A(_1445_),
    .X(_1446_));
 sky130_fd_sc_hd__or2_1 _6418_ (.A(_1446_),
    .B(_1384_),
    .X(_1447_));
 sky130_fd_sc_hd__nand2_1 _6419_ (.A(_1447_),
    .B(_0105_),
    .Y(_1448_));
 sky130_fd_sc_hd__nor2_1 _6420_ (.A(_1446_),
    .B(_1401_),
    .Y(_1449_));
 sky130_fd_sc_hd__and3_1 _6421_ (.A(_4211_),
    .B(_1449_),
    .C(_0148_),
    .X(_1450_));
 sky130_fd_sc_hd__and3b_1 _6422_ (.A_N(_0148_),
    .B(_1449_),
    .C(_4213_),
    .X(_1452_));
 sky130_fd_sc_hd__nor2_1 _6423_ (.A(_1450_),
    .B(_1452_),
    .Y(_1453_));
 sky130_fd_sc_hd__clkbuf_4 _6424_ (.A(_3795_),
    .X(_1454_));
 sky130_fd_sc_hd__or2_1 _6425_ (.A(_1445_),
    .B(_1454_),
    .X(_1455_));
 sky130_fd_sc_hd__clkbuf_4 _6426_ (.A(_3930_),
    .X(_1456_));
 sky130_fd_sc_hd__or4_2 _6427_ (.A(_4250_),
    .B(_0147_),
    .C(_1455_),
    .D(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__nand2_1 _6428_ (.A(_1448_),
    .B(_1453_),
    .Y(_1458_));
 sky130_fd_sc_hd__xnor2_1 _6429_ (.A(_1435_),
    .B(_1458_),
    .Y(_1459_));
 sky130_fd_sc_hd__and2b_1 _6430_ (.A_N(_1457_),
    .B(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__a31o_1 _6431_ (.A1(_1435_),
    .A2(_1448_),
    .A3(_1453_),
    .B1(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__nor2_1 _6432_ (.A(_0082_),
    .B(_1423_),
    .Y(_1463_));
 sky130_fd_sc_hd__or2_1 _6433_ (.A(_1420_),
    .B(_1399_),
    .X(_1464_));
 sky130_fd_sc_hd__nand3_1 _6434_ (.A(_0218_),
    .B(_1353_),
    .C(_1354_),
    .Y(_1465_));
 sky130_fd_sc_hd__nor2_1 _6435_ (.A(_1383_),
    .B(_0303_),
    .Y(_1466_));
 sky130_fd_sc_hd__xnor2_1 _6436_ (.A(_1465_),
    .B(_1466_),
    .Y(_1467_));
 sky130_fd_sc_hd__xnor2_1 _6437_ (.A(_1464_),
    .B(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__or2_1 _6438_ (.A(_4232_),
    .B(_1410_),
    .X(_1469_));
 sky130_fd_sc_hd__nor2_1 _6439_ (.A(_0080_),
    .B(_1423_),
    .Y(_1470_));
 sky130_fd_sc_hd__and2b_1 _6440_ (.A_N(_1469_),
    .B(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__xnor2_1 _6441_ (.A(_1468_),
    .B(_1471_),
    .Y(_1472_));
 sky130_fd_sc_hd__nor2_1 _6442_ (.A(_1399_),
    .B(_1428_),
    .Y(_1474_));
 sky130_fd_sc_hd__and3_1 _6443_ (.A(_4217_),
    .B(_1353_),
    .C(_1354_),
    .X(_1475_));
 sky130_fd_sc_hd__or2_1 _6444_ (.A(_1383_),
    .B(_3840_),
    .X(_1476_));
 sky130_fd_sc_hd__xnor2_1 _6445_ (.A(_1475_),
    .B(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__a22oi_2 _6446_ (.A1(_1466_),
    .A2(_1427_),
    .B1(_1474_),
    .B2(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__xor2_1 _6447_ (.A(_1472_),
    .B(_1478_),
    .X(_1479_));
 sky130_fd_sc_hd__xnor2_1 _6448_ (.A(_1463_),
    .B(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__a22o_1 _6449_ (.A1(_1427_),
    .A2(_1430_),
    .B1(_1426_),
    .B2(_1431_),
    .X(_1481_));
 sky130_fd_sc_hd__inv_2 _6450_ (.A(_1423_),
    .Y(_1482_));
 sky130_fd_sc_hd__a32o_1 _6451_ (.A1(_0218_),
    .A2(_1408_),
    .A3(_1409_),
    .B1(_1414_),
    .B2(_0121_),
    .X(_1483_));
 sky130_fd_sc_hd__o21a_1 _6452_ (.A1(_1469_),
    .A2(_1416_),
    .B1(_1483_),
    .X(_1485_));
 sky130_fd_sc_hd__nor2_1 _6453_ (.A(_1469_),
    .B(_1416_),
    .Y(_1486_));
 sky130_fd_sc_hd__a31o_1 _6454_ (.A1(_4217_),
    .A2(_1482_),
    .A3(_1485_),
    .B1(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__xor2_1 _6455_ (.A(_1474_),
    .B(_1477_),
    .X(_1488_));
 sky130_fd_sc_hd__xor2_1 _6456_ (.A(_1487_),
    .B(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__xor2_1 _6457_ (.A(_1481_),
    .B(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__xnor2_1 _6458_ (.A(_1469_),
    .B(_1470_),
    .Y(_1491_));
 sky130_fd_sc_hd__and2_1 _6459_ (.A(_1490_),
    .B(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__xnor2_1 _6460_ (.A(_1480_),
    .B(_1492_),
    .Y(_1493_));
 sky130_fd_sc_hd__nand2_1 _6461_ (.A(_1487_),
    .B(_1488_),
    .Y(_1494_));
 sky130_fd_sc_hd__a21boi_1 _6462_ (.A1(_1481_),
    .A2(_1489_),
    .B1_N(_1494_),
    .Y(_1496_));
 sky130_fd_sc_hd__or2_1 _6463_ (.A(_1446_),
    .B(_1428_),
    .X(_1497_));
 sky130_fd_sc_hd__nor2_1 _6464_ (.A(_4250_),
    .B(_1428_),
    .Y(_1498_));
 sky130_fd_sc_hd__or3_1 _6465_ (.A(_1498_),
    .B(_1447_),
    .C(_0105_),
    .X(_1499_));
 sky130_fd_sc_hd__or3_1 _6466_ (.A(_1497_),
    .B(_4211_),
    .C(_1449_),
    .X(_1500_));
 sky130_fd_sc_hd__nand2_1 _6467_ (.A(_1499_),
    .B(_1500_),
    .Y(_1501_));
 sky130_fd_sc_hd__a21o_1 _6468_ (.A1(_1497_),
    .A2(_4211_),
    .B1(_1501_),
    .X(_1502_));
 sky130_fd_sc_hd__xor2_1 _6469_ (.A(_1496_),
    .B(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__xor2_1 _6470_ (.A(_1503_),
    .B(_1450_),
    .X(_1504_));
 sky130_fd_sc_hd__xnor2_1 _6471_ (.A(_1493_),
    .B(_1504_),
    .Y(_1505_));
 sky130_fd_sc_hd__xnor2_1 _6472_ (.A(_1490_),
    .B(_1491_),
    .Y(_1507_));
 sky130_fd_sc_hd__o31a_1 _6473_ (.A1(_1191_),
    .A2(_1226_),
    .A3(_1305_),
    .B1(_1309_),
    .X(_1508_));
 sky130_fd_sc_hd__xnor2_2 _6474_ (.A(_1157_),
    .B(_1508_),
    .Y(_1509_));
 sky130_fd_sc_hd__buf_4 _6475_ (.A(_1509_),
    .X(_1510_));
 sky130_fd_sc_hd__nor2_4 _6476_ (.A(_4232_),
    .B(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__xor2_2 _6477_ (.A(_1416_),
    .B(_1417_),
    .X(_1512_));
 sky130_fd_sc_hd__xnor2_4 _6478_ (.A(_1512_),
    .B(_1424_),
    .Y(_1513_));
 sky130_fd_sc_hd__or2_1 _6479_ (.A(_0303_),
    .B(_1423_),
    .X(_1514_));
 sky130_fd_sc_hd__xnor2_1 _6480_ (.A(_1514_),
    .B(_1485_),
    .Y(_1515_));
 sky130_fd_sc_hd__and3_1 _6481_ (.A(_1511_),
    .B(_1513_),
    .C(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__a21oi_1 _6482_ (.A1(_1511_),
    .A2(_1513_),
    .B1(_1515_),
    .Y(_1518_));
 sky130_fd_sc_hd__nor2_1 _6483_ (.A(_1516_),
    .B(_1518_),
    .Y(_1519_));
 sky130_fd_sc_hd__xor2_1 _6484_ (.A(_1404_),
    .B(_1433_),
    .X(_1520_));
 sky130_fd_sc_hd__a21o_1 _6485_ (.A1(_1519_),
    .A2(_1520_),
    .B1(_1516_),
    .X(_1521_));
 sky130_fd_sc_hd__xnor2_1 _6486_ (.A(_1507_),
    .B(_1521_),
    .Y(_1522_));
 sky130_fd_sc_hd__xnor2_1 _6487_ (.A(_1457_),
    .B(_1459_),
    .Y(_1523_));
 sky130_fd_sc_hd__and2b_1 _6488_ (.A_N(_1507_),
    .B(_1521_),
    .X(_1524_));
 sky130_fd_sc_hd__a21oi_1 _6489_ (.A1(_1522_),
    .A2(_1523_),
    .B1(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__nor2_1 _6490_ (.A(_1505_),
    .B(_1525_),
    .Y(_1526_));
 sky130_fd_sc_hd__nand2_1 _6491_ (.A(_1505_),
    .B(_1525_),
    .Y(_1527_));
 sky130_fd_sc_hd__and2b_1 _6492_ (.A_N(_1526_),
    .B(_1527_),
    .X(_1529_));
 sky130_fd_sc_hd__xnor2_1 _6493_ (.A(_1461_),
    .B(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hd__buf_4 _6494_ (.A(_3907_),
    .X(_1531_));
 sky130_fd_sc_hd__o21a_1 _6495_ (.A1(_1443_),
    .A2(_1444_),
    .B1(_1531_),
    .X(_1532_));
 sky130_fd_sc_hd__nor2_1 _6496_ (.A(_1446_),
    .B(_1456_),
    .Y(_1533_));
 sky130_fd_sc_hd__nor2_1 _6497_ (.A(_4157_),
    .B(_1533_),
    .Y(_1534_));
 sky130_fd_sc_hd__or3_1 _6498_ (.A(_1191_),
    .B(_1226_),
    .C(_1305_),
    .X(_1535_));
 sky130_fd_sc_hd__o21ai_1 _6499_ (.A1(_1226_),
    .A2(_1305_),
    .B1(_1191_),
    .Y(_1536_));
 sky130_fd_sc_hd__nand2_4 _6500_ (.A(_1535_),
    .B(_1536_),
    .Y(_1537_));
 sky130_fd_sc_hd__clkbuf_4 _6501_ (.A(_1537_),
    .X(_1538_));
 sky130_fd_sc_hd__or2_1 _6502_ (.A(_0082_),
    .B(_1538_),
    .X(_1540_));
 sky130_fd_sc_hd__o2bb2a_1 _6503_ (.A1_N(_1532_),
    .A2_N(_0184_),
    .B1(_1534_),
    .B2(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__xor2_2 _6504_ (.A(_1455_),
    .B(_0184_),
    .X(_1542_));
 sky130_fd_sc_hd__nor2_1 _6505_ (.A(_1541_),
    .B(_1542_),
    .Y(_1543_));
 sky130_fd_sc_hd__and3_1 _6506_ (.A(_1353_),
    .B(_1354_),
    .C(_0147_),
    .X(_1544_));
 sky130_fd_sc_hd__or2_1 _6507_ (.A(_1383_),
    .B(_1401_),
    .X(_1545_));
 sky130_fd_sc_hd__and3_1 _6508_ (.A(_1353_),
    .B(_1354_),
    .C(_3986_),
    .X(_1546_));
 sky130_fd_sc_hd__xnor2_2 _6509_ (.A(_1545_),
    .B(_1546_),
    .Y(_1547_));
 sky130_fd_sc_hd__nor2_1 _6510_ (.A(_1400_),
    .B(_1454_),
    .Y(_1548_));
 sky130_fd_sc_hd__a22oi_4 _6511_ (.A1(_1544_),
    .A2(_1386_),
    .B1(_1547_),
    .B2(_1548_),
    .Y(_1549_));
 sky130_fd_sc_hd__nand2_1 _6512_ (.A(_4153_),
    .B(_1414_),
    .Y(_1551_));
 sky130_fd_sc_hd__o21ai_1 _6513_ (.A1(_1420_),
    .A2(_1410_),
    .B1(_1415_),
    .Y(_1552_));
 sky130_fd_sc_hd__o21a_2 _6514_ (.A1(_1551_),
    .A2(_1417_),
    .B1(_1552_),
    .X(_1553_));
 sky130_fd_sc_hd__nor2_2 _6515_ (.A(_1428_),
    .B(_1423_),
    .Y(_1554_));
 sky130_fd_sc_hd__a2bb2o_1 _6516_ (.A1_N(_1551_),
    .A2_N(_1417_),
    .B1(_1553_),
    .B2(_1554_),
    .X(_1555_));
 sky130_fd_sc_hd__xor2_1 _6517_ (.A(_1402_),
    .B(_1403_),
    .X(_1556_));
 sky130_fd_sc_hd__xnor2_1 _6518_ (.A(_1555_),
    .B(_1556_),
    .Y(_1557_));
 sky130_fd_sc_hd__nand2_1 _6519_ (.A(_1555_),
    .B(_1556_),
    .Y(_1558_));
 sky130_fd_sc_hd__o21a_1 _6520_ (.A1(_1549_),
    .A2(_1557_),
    .B1(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__or3_1 _6521_ (.A(_0105_),
    .B(_1455_),
    .C(_0184_),
    .X(_1560_));
 sky130_fd_sc_hd__o211a_1 _6522_ (.A1(_1449_),
    .A2(_0148_),
    .B1(_1457_),
    .C1(_1560_),
    .X(_1562_));
 sky130_fd_sc_hd__xnor2_1 _6523_ (.A(_1559_),
    .B(_1562_),
    .Y(_1563_));
 sky130_fd_sc_hd__or2b_1 _6524_ (.A(_1559_),
    .B_N(_1562_),
    .X(_1564_));
 sky130_fd_sc_hd__a21bo_1 _6525_ (.A1(_1543_),
    .A2(_1563_),
    .B1_N(_1564_),
    .X(_1565_));
 sky130_fd_sc_hd__xor2_4 _6526_ (.A(_1553_),
    .B(_1554_),
    .X(_1566_));
 sky130_fd_sc_hd__nor2_2 _6527_ (.A(_0080_),
    .B(_1510_),
    .Y(_1567_));
 sky130_fd_sc_hd__xor2_4 _6528_ (.A(_1511_),
    .B(_1513_),
    .X(_1568_));
 sky130_fd_sc_hd__nand2_1 _6529_ (.A(_1566_),
    .B(_1567_),
    .Y(_1569_));
 sky130_fd_sc_hd__xnor2_2 _6530_ (.A(_1569_),
    .B(_1568_),
    .Y(_1570_));
 sky130_fd_sc_hd__xor2_2 _6531_ (.A(_1549_),
    .B(_1557_),
    .X(_1571_));
 sky130_fd_sc_hd__a32oi_4 _6532_ (.A1(_1566_),
    .A2(_1567_),
    .A3(_1568_),
    .B1(_1570_),
    .B2(_1571_),
    .Y(_1573_));
 sky130_fd_sc_hd__xnor2_1 _6533_ (.A(_1519_),
    .B(_1520_),
    .Y(_1574_));
 sky130_fd_sc_hd__xor2_1 _6534_ (.A(_1573_),
    .B(_1574_),
    .X(_1575_));
 sky130_fd_sc_hd__xor2_1 _6535_ (.A(_1543_),
    .B(_1563_),
    .X(_1576_));
 sky130_fd_sc_hd__nor2_1 _6536_ (.A(_1573_),
    .B(_1574_),
    .Y(_1577_));
 sky130_fd_sc_hd__a21o_1 _6537_ (.A1(_1575_),
    .A2(_1576_),
    .B1(_1577_),
    .X(_1578_));
 sky130_fd_sc_hd__xnor2_1 _6538_ (.A(_1522_),
    .B(_1523_),
    .Y(_1579_));
 sky130_fd_sc_hd__xnor2_1 _6539_ (.A(_1578_),
    .B(_1579_),
    .Y(_1580_));
 sky130_fd_sc_hd__and2b_1 _6540_ (.A_N(_1579_),
    .B(_1578_),
    .X(_1581_));
 sky130_fd_sc_hd__a21oi_1 _6541_ (.A1(_1565_),
    .A2(_1580_),
    .B1(_1581_),
    .Y(_1582_));
 sky130_fd_sc_hd__nor2_1 _6542_ (.A(_1530_),
    .B(_1582_),
    .Y(_1584_));
 sky130_fd_sc_hd__a2bb2o_1 _6543_ (.A1_N(_1496_),
    .A2_N(_1502_),
    .B1(_1503_),
    .B2(_1450_),
    .X(_1585_));
 sky130_fd_sc_hd__nand2_1 _6544_ (.A(_1468_),
    .B(_1471_),
    .Y(_1586_));
 sky130_fd_sc_hd__o21ai_1 _6545_ (.A1(_1472_),
    .A2(_1478_),
    .B1(_1586_),
    .Y(_1587_));
 sky130_fd_sc_hd__nor2_1 _6546_ (.A(_1420_),
    .B(_1446_),
    .Y(_1588_));
 sky130_fd_sc_hd__a21o_1 _6547_ (.A1(_1498_),
    .A2(_1447_),
    .B1(_1588_),
    .X(_1589_));
 sky130_fd_sc_hd__o31a_1 _6548_ (.A1(_4219_),
    .A2(_1497_),
    .A3(_4213_),
    .B1(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__xor2_1 _6549_ (.A(_1587_),
    .B(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__xnor2_1 _6550_ (.A(_1499_),
    .B(_1591_),
    .Y(_1592_));
 sky130_fd_sc_hd__or2_1 _6551_ (.A(_4228_),
    .B(_1383_),
    .X(_1593_));
 sky130_fd_sc_hd__and2b_1 _6552_ (.A_N(_1593_),
    .B(_1475_),
    .X(_1595_));
 sky130_fd_sc_hd__inv_2 _6553_ (.A(_1400_),
    .Y(_1596_));
 sky130_fd_sc_hd__and3_1 _6554_ (.A(_4153_),
    .B(_1596_),
    .C(_1467_),
    .X(_1597_));
 sky130_fd_sc_hd__or2_1 _6555_ (.A(_0303_),
    .B(_1400_),
    .X(_1598_));
 sky130_fd_sc_hd__nand2_1 _6556_ (.A(_1353_),
    .B(_1354_),
    .Y(_1599_));
 sky130_fd_sc_hd__or2_1 _6557_ (.A(_1599_),
    .B(_4232_),
    .X(_1600_));
 sky130_fd_sc_hd__xnor2_1 _6558_ (.A(_1593_),
    .B(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__xor2_1 _6559_ (.A(_1598_),
    .B(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__o21ai_1 _6560_ (.A1(_1595_),
    .A2(_1597_),
    .B1(_1602_),
    .Y(_1603_));
 sky130_fd_sc_hd__or3_1 _6561_ (.A(_1595_),
    .B(_1597_),
    .C(_1602_),
    .X(_1604_));
 sky130_fd_sc_hd__nand2_1 _6562_ (.A(_1603_),
    .B(_1604_),
    .Y(_1606_));
 sky130_fd_sc_hd__nand2_1 _6563_ (.A(_1463_),
    .B(_1479_),
    .Y(_1607_));
 sky130_fd_sc_hd__xor2_1 _6564_ (.A(_1606_),
    .B(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__xnor2_1 _6565_ (.A(_1592_),
    .B(_1608_),
    .Y(_1609_));
 sky130_fd_sc_hd__and2b_1 _6566_ (.A_N(_1480_),
    .B(_1492_),
    .X(_1610_));
 sky130_fd_sc_hd__a21oi_1 _6567_ (.A1(_1493_),
    .A2(_1504_),
    .B1(_1610_),
    .Y(_1611_));
 sky130_fd_sc_hd__nor2_1 _6568_ (.A(_1609_),
    .B(_1611_),
    .Y(_1612_));
 sky130_fd_sc_hd__nand2_1 _6569_ (.A(_1609_),
    .B(_1611_),
    .Y(_1613_));
 sky130_fd_sc_hd__and2b_1 _6570_ (.A_N(_1612_),
    .B(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__xnor2_1 _6571_ (.A(_1585_),
    .B(_1614_),
    .Y(_1615_));
 sky130_fd_sc_hd__a21oi_1 _6572_ (.A1(_1461_),
    .A2(_1527_),
    .B1(_1526_),
    .Y(_1617_));
 sky130_fd_sc_hd__xor2_1 _6573_ (.A(_1615_),
    .B(_1617_),
    .X(_1618_));
 sky130_fd_sc_hd__xnor2_1 _6574_ (.A(_1584_),
    .B(_1618_),
    .Y(_1619_));
 sky130_fd_sc_hd__or2_1 _6575_ (.A(_1615_),
    .B(_1617_),
    .X(_1620_));
 sky130_fd_sc_hd__and2b_1 _6576_ (.A_N(_1499_),
    .B(_1591_),
    .X(_1621_));
 sky130_fd_sc_hd__a21o_1 _6577_ (.A1(_1587_),
    .A2(_1590_),
    .B1(_1621_),
    .X(_1622_));
 sky130_fd_sc_hd__and3b_1 _6578_ (.A_N(_1497_),
    .B(_4213_),
    .C(_4219_),
    .X(_1623_));
 sky130_fd_sc_hd__or2_1 _6579_ (.A(_1420_),
    .B(_1446_),
    .X(_1624_));
 sky130_fd_sc_hd__nor2_1 _6580_ (.A(_0303_),
    .B(_1446_),
    .Y(_1625_));
 sky130_fd_sc_hd__a21o_1 _6581_ (.A1(_4235_),
    .A2(_1497_),
    .B1(_1625_),
    .X(_1626_));
 sky130_fd_sc_hd__o31a_1 _6582_ (.A1(_1624_),
    .A2(_4251_),
    .A3(_1498_),
    .B1(_1626_),
    .X(_1628_));
 sky130_fd_sc_hd__xnor2_1 _6583_ (.A(_1603_),
    .B(_1628_),
    .Y(_1629_));
 sky130_fd_sc_hd__xor2_1 _6584_ (.A(_1623_),
    .B(_1629_),
    .X(_1630_));
 sky130_fd_sc_hd__or2_1 _6585_ (.A(_1383_),
    .B(_0082_),
    .X(_1631_));
 sky130_fd_sc_hd__or2_1 _6586_ (.A(_1465_),
    .B(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__or2_1 _6587_ (.A(_1598_),
    .B(_1601_),
    .X(_1633_));
 sky130_fd_sc_hd__or3_1 _6588_ (.A(_0080_),
    .B(_1400_),
    .C(_1631_),
    .X(_1634_));
 sky130_fd_sc_hd__o21ai_1 _6589_ (.A1(_0080_),
    .A2(_1400_),
    .B1(_1631_),
    .Y(_1635_));
 sky130_fd_sc_hd__and2_1 _6590_ (.A(_1634_),
    .B(_1635_),
    .X(_1636_));
 sky130_fd_sc_hd__a21bo_1 _6591_ (.A1(_1632_),
    .A2(_1633_),
    .B1_N(_1636_),
    .X(_1637_));
 sky130_fd_sc_hd__nand2_1 _6592_ (.A(_1632_),
    .B(_1633_),
    .Y(_1639_));
 sky130_fd_sc_hd__or2_1 _6593_ (.A(_1639_),
    .B(_1636_),
    .X(_1640_));
 sky130_fd_sc_hd__and2_1 _6594_ (.A(_1637_),
    .B(_1640_),
    .X(_1641_));
 sky130_fd_sc_hd__nand2_1 _6595_ (.A(_1630_),
    .B(_1641_),
    .Y(_1642_));
 sky130_fd_sc_hd__or2_1 _6596_ (.A(_1630_),
    .B(_1641_),
    .X(_1643_));
 sky130_fd_sc_hd__nand2_1 _6597_ (.A(_1642_),
    .B(_1643_),
    .Y(_1644_));
 sky130_fd_sc_hd__nand2_1 _6598_ (.A(_1592_),
    .B(_1608_),
    .Y(_1645_));
 sky130_fd_sc_hd__o21a_1 _6599_ (.A1(_1606_),
    .A2(_1607_),
    .B1(_1645_),
    .X(_1646_));
 sky130_fd_sc_hd__xor2_1 _6600_ (.A(_1644_),
    .B(_1646_),
    .X(_1647_));
 sky130_fd_sc_hd__xnor2_1 _6601_ (.A(_1622_),
    .B(_1647_),
    .Y(_1648_));
 sky130_fd_sc_hd__a21oi_1 _6602_ (.A1(_1585_),
    .A2(_1613_),
    .B1(_1612_),
    .Y(_1650_));
 sky130_fd_sc_hd__xnor2_1 _6603_ (.A(_1648_),
    .B(_1650_),
    .Y(_1651_));
 sky130_fd_sc_hd__xnor2_1 _6604_ (.A(_1620_),
    .B(_1651_),
    .Y(_1652_));
 sky130_fd_sc_hd__or2_1 _6605_ (.A(_1619_),
    .B(_1652_),
    .X(_1653_));
 sky130_fd_sc_hd__nor2_2 _6606_ (.A(_0303_),
    .B(_1510_),
    .Y(_1654_));
 sky130_fd_sc_hd__or2_2 _6607_ (.A(_1428_),
    .B(_1410_),
    .X(_1655_));
 sky130_fd_sc_hd__xor2_2 _6608_ (.A(_1655_),
    .B(_1551_),
    .X(_1656_));
 sky130_fd_sc_hd__nor2_1 _6609_ (.A(_1384_),
    .B(_1423_),
    .Y(_1657_));
 sky130_fd_sc_hd__xor2_2 _6610_ (.A(_1656_),
    .B(_1657_),
    .X(_1658_));
 sky130_fd_sc_hd__xnor2_1 _6611_ (.A(_1654_),
    .B(_1658_),
    .Y(_1659_));
 sky130_fd_sc_hd__nor2_1 _6612_ (.A(_1420_),
    .B(_1510_),
    .Y(_1661_));
 sky130_fd_sc_hd__and2_1 _6613_ (.A(_1301_),
    .B(_1300_),
    .X(_1662_));
 sky130_fd_sc_hd__a21bo_1 _6614_ (.A1(_1277_),
    .A2(_1662_),
    .B1_N(_1302_),
    .X(_1663_));
 sky130_fd_sc_hd__buf_2 _6615_ (.A(_1663_),
    .X(_1664_));
 sky130_fd_sc_hd__nor2_2 _6616_ (.A(_4037_),
    .B(_1664_),
    .Y(_1665_));
 sky130_fd_sc_hd__nand2_1 _6617_ (.A(_1665_),
    .B(_1511_),
    .Y(_1666_));
 sky130_fd_sc_hd__mux2_1 _6618_ (.A0(_1420_),
    .A1(_1661_),
    .S(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__nand2_2 _6619_ (.A(_3986_),
    .B(_1414_),
    .Y(_1668_));
 sky130_fd_sc_hd__o2bb2a_1 _6620_ (.A1_N(_1355_),
    .A2_N(_1414_),
    .B1(_1410_),
    .B2(_1384_),
    .X(_1669_));
 sky130_fd_sc_hd__o21ba_1 _6621_ (.A1(_1655_),
    .A2(_1668_),
    .B1_N(_1669_),
    .X(_1670_));
 sky130_fd_sc_hd__or2_1 _6622_ (.A(_1423_),
    .B(_1401_),
    .X(_1672_));
 sky130_fd_sc_hd__xnor2_1 _6623_ (.A(_1670_),
    .B(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__o2bb2a_1 _6624_ (.A1_N(_1667_),
    .A2_N(_1673_),
    .B1(_1420_),
    .B2(_1666_),
    .X(_1674_));
 sky130_fd_sc_hd__xor2_1 _6625_ (.A(_1659_),
    .B(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__buf_4 _6626_ (.A(_3703_),
    .X(_1676_));
 sky130_fd_sc_hd__or2_1 _6627_ (.A(_1382_),
    .B(_1456_),
    .X(_1677_));
 sky130_fd_sc_hd__nand3_1 _6628_ (.A(_1353_),
    .B(_1354_),
    .C(_4089_),
    .Y(_1678_));
 sky130_fd_sc_hd__xnor2_1 _6629_ (.A(_1677_),
    .B(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__or2_1 _6630_ (.A(_1677_),
    .B(_1678_),
    .X(_1680_));
 sky130_fd_sc_hd__o31a_1 _6631_ (.A1(_1400_),
    .A2(_1676_),
    .A3(_1679_),
    .B1(_1680_),
    .X(_1681_));
 sky130_fd_sc_hd__o22ai_2 _6632_ (.A1(_1655_),
    .A2(_1668_),
    .B1(_1672_),
    .B2(_1669_),
    .Y(_1683_));
 sky130_fd_sc_hd__or2_1 _6633_ (.A(_1383_),
    .B(_1454_),
    .X(_1684_));
 sky130_fd_sc_hd__xnor2_1 _6634_ (.A(_1684_),
    .B(_1544_),
    .Y(_1685_));
 sky130_fd_sc_hd__nor2_1 _6635_ (.A(_1400_),
    .B(_1456_),
    .Y(_1686_));
 sky130_fd_sc_hd__xor2_2 _6636_ (.A(_1685_),
    .B(_1686_),
    .X(_1687_));
 sky130_fd_sc_hd__xor2_1 _6637_ (.A(_1683_),
    .B(_1687_),
    .X(_1688_));
 sky130_fd_sc_hd__xnor2_1 _6638_ (.A(_1681_),
    .B(_1688_),
    .Y(_1689_));
 sky130_fd_sc_hd__nor2_1 _6639_ (.A(_1659_),
    .B(_1674_),
    .Y(_1690_));
 sky130_fd_sc_hd__a21oi_1 _6640_ (.A1(_1675_),
    .A2(_1689_),
    .B1(_1690_),
    .Y(_1691_));
 sky130_fd_sc_hd__nand2_1 _6641_ (.A(_1654_),
    .B(_1658_),
    .Y(_1692_));
 sky130_fd_sc_hd__xor2_2 _6642_ (.A(_1566_),
    .B(_1567_),
    .X(_1694_));
 sky130_fd_sc_hd__xnor2_2 _6643_ (.A(_1692_),
    .B(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__a2bb2o_1 _6644_ (.A1_N(_1678_),
    .A2_N(_1545_),
    .B1(_1685_),
    .B2(_1686_),
    .X(_1696_));
 sky130_fd_sc_hd__a2bb2oi_1 _6645_ (.A1_N(_1655_),
    .A2_N(_1551_),
    .B1(_1656_),
    .B2(_1657_),
    .Y(_1697_));
 sky130_fd_sc_hd__xor2_1 _6646_ (.A(_1548_),
    .B(_1547_),
    .X(_1698_));
 sky130_fd_sc_hd__xnor2_1 _6647_ (.A(_1697_),
    .B(_1698_),
    .Y(_1699_));
 sky130_fd_sc_hd__xor2_2 _6648_ (.A(_1696_),
    .B(_1699_),
    .X(_1700_));
 sky130_fd_sc_hd__xnor2_1 _6649_ (.A(_1695_),
    .B(_1700_),
    .Y(_1701_));
 sky130_fd_sc_hd__xor2_1 _6650_ (.A(_1691_),
    .B(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__or2_1 _6651_ (.A(_0548_),
    .B(_1537_),
    .X(_1703_));
 sky130_fd_sc_hd__inv_2 _6652_ (.A(_1703_),
    .Y(_1705_));
 sky130_fd_sc_hd__nand2_1 _6653_ (.A(_1625_),
    .B(_1705_),
    .Y(_1706_));
 sky130_fd_sc_hd__xor2_1 _6654_ (.A(_4018_),
    .B(_1532_),
    .X(_1707_));
 sky130_fd_sc_hd__nor2_1 _6655_ (.A(_0080_),
    .B(_1538_),
    .Y(_1708_));
 sky130_fd_sc_hd__xnor2_1 _6656_ (.A(_1707_),
    .B(_1708_),
    .Y(_1709_));
 sky130_fd_sc_hd__xor2_1 _6657_ (.A(_1706_),
    .B(_1709_),
    .X(_1710_));
 sky130_fd_sc_hd__or2_2 _6658_ (.A(_1257_),
    .B(_1302_),
    .X(_1711_));
 sky130_fd_sc_hd__a21oi_1 _6659_ (.A1(_1221_),
    .A2(_1224_),
    .B1(_1225_),
    .Y(_1712_));
 sky130_fd_sc_hd__or2_1 _6660_ (.A(_1712_),
    .B(_1226_),
    .X(_1713_));
 sky130_fd_sc_hd__a21oi_1 _6661_ (.A1(_1304_),
    .A2(_1711_),
    .B1(_1713_),
    .Y(_1714_));
 sky130_fd_sc_hd__and3_1 _6662_ (.A(_1304_),
    .B(_1711_),
    .C(_1713_),
    .X(_1716_));
 sky130_fd_sc_hd__or2_1 _6663_ (.A(_1714_),
    .B(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__buf_2 _6664_ (.A(_1717_),
    .X(_1718_));
 sky130_fd_sc_hd__nor2_1 _6665_ (.A(_0082_),
    .B(_1718_),
    .Y(_1719_));
 sky130_fd_sc_hd__nor2_1 _6666_ (.A(_1706_),
    .B(_1709_),
    .Y(_1720_));
 sky130_fd_sc_hd__a21o_1 _6667_ (.A1(_1710_),
    .A2(_1719_),
    .B1(_1720_),
    .X(_1721_));
 sky130_fd_sc_hd__nor2_1 _6668_ (.A(_1683_),
    .B(_1687_),
    .Y(_1722_));
 sky130_fd_sc_hd__nand2_1 _6669_ (.A(_1683_),
    .B(_1687_),
    .Y(_1723_));
 sky130_fd_sc_hd__o21a_1 _6670_ (.A1(_1681_),
    .A2(_1722_),
    .B1(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__nor2_1 _6671_ (.A(_1446_),
    .B(_0548_),
    .Y(_1725_));
 sky130_fd_sc_hd__a22o_1 _6672_ (.A1(_1725_),
    .A2(_4157_),
    .B1(_1707_),
    .B2(_1708_),
    .X(_1727_));
 sky130_fd_sc_hd__xor2_1 _6673_ (.A(_4157_),
    .B(_1533_),
    .X(_1728_));
 sky130_fd_sc_hd__xnor2_1 _6674_ (.A(_1540_),
    .B(_1728_),
    .Y(_1729_));
 sky130_fd_sc_hd__xnor2_1 _6675_ (.A(_1727_),
    .B(_1729_),
    .Y(_1730_));
 sky130_fd_sc_hd__xnor2_1 _6676_ (.A(_1724_),
    .B(_1730_),
    .Y(_1731_));
 sky130_fd_sc_hd__xnor2_1 _6677_ (.A(_1721_),
    .B(_1731_),
    .Y(_1732_));
 sky130_fd_sc_hd__nor2_1 _6678_ (.A(_1691_),
    .B(_1701_),
    .Y(_1733_));
 sky130_fd_sc_hd__a21oi_1 _6679_ (.A1(_1702_),
    .A2(_1732_),
    .B1(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__a32oi_4 _6680_ (.A1(_1654_),
    .A2(_1658_),
    .A3(_1694_),
    .B1(_1695_),
    .B2(_1700_),
    .Y(_1735_));
 sky130_fd_sc_hd__xnor2_1 _6681_ (.A(_1570_),
    .B(_1571_),
    .Y(_1736_));
 sky130_fd_sc_hd__xor2_1 _6682_ (.A(_1735_),
    .B(_1736_),
    .X(_1738_));
 sky130_fd_sc_hd__nand2_1 _6683_ (.A(_1727_),
    .B(_1729_),
    .Y(_1739_));
 sky130_fd_sc_hd__or2b_1 _6684_ (.A(_1697_),
    .B_N(_1698_),
    .X(_1740_));
 sky130_fd_sc_hd__a21bo_1 _6685_ (.A1(_1696_),
    .A2(_1699_),
    .B1_N(_1740_),
    .X(_1741_));
 sky130_fd_sc_hd__xnor2_1 _6686_ (.A(_1541_),
    .B(_1542_),
    .Y(_1742_));
 sky130_fd_sc_hd__xor2_1 _6687_ (.A(_1741_),
    .B(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__xor2_1 _6688_ (.A(_1739_),
    .B(_1743_),
    .X(_1744_));
 sky130_fd_sc_hd__xnor2_1 _6689_ (.A(_1738_),
    .B(_1744_),
    .Y(_1745_));
 sky130_fd_sc_hd__or2_1 _6690_ (.A(_1734_),
    .B(_1745_),
    .X(_1746_));
 sky130_fd_sc_hd__nand2_1 _6691_ (.A(_1724_),
    .B(_1730_),
    .Y(_1747_));
 sky130_fd_sc_hd__nor2_1 _6692_ (.A(_1724_),
    .B(_1730_),
    .Y(_1749_));
 sky130_fd_sc_hd__a21o_1 _6693_ (.A1(_1721_),
    .A2(_1747_),
    .B1(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__xor2_1 _6694_ (.A(_1734_),
    .B(_1745_),
    .X(_1751_));
 sky130_fd_sc_hd__nand2_1 _6695_ (.A(_1750_),
    .B(_1751_),
    .Y(_1752_));
 sky130_fd_sc_hd__or2b_1 _6696_ (.A(_1742_),
    .B_N(_1741_),
    .X(_1753_));
 sky130_fd_sc_hd__o21ai_1 _6697_ (.A1(_1739_),
    .A2(_1743_),
    .B1(_1753_),
    .Y(_1754_));
 sky130_fd_sc_hd__nor2_1 _6698_ (.A(_1735_),
    .B(_1736_),
    .Y(_1755_));
 sky130_fd_sc_hd__a21o_1 _6699_ (.A1(_1738_),
    .A2(_1744_),
    .B1(_1755_),
    .X(_1756_));
 sky130_fd_sc_hd__xor2_1 _6700_ (.A(_1575_),
    .B(_1576_),
    .X(_1757_));
 sky130_fd_sc_hd__xnor2_1 _6701_ (.A(_1756_),
    .B(_1757_),
    .Y(_1758_));
 sky130_fd_sc_hd__xor2_1 _6702_ (.A(_1754_),
    .B(_1758_),
    .X(_1760_));
 sky130_fd_sc_hd__a21o_1 _6703_ (.A1(_1746_),
    .A2(_1752_),
    .B1(_1760_),
    .X(_1761_));
 sky130_fd_sc_hd__nand2_1 _6704_ (.A(_1756_),
    .B(_1757_),
    .Y(_1762_));
 sky130_fd_sc_hd__or2b_1 _6705_ (.A(_1758_),
    .B_N(_1754_),
    .X(_1763_));
 sky130_fd_sc_hd__xnor2_1 _6706_ (.A(_1565_),
    .B(_1580_),
    .Y(_1764_));
 sky130_fd_sc_hd__a21o_1 _6707_ (.A1(_1762_),
    .A2(_1763_),
    .B1(_1764_),
    .X(_1765_));
 sky130_fd_sc_hd__nand3_1 _6708_ (.A(_1762_),
    .B(_1763_),
    .C(_1764_),
    .Y(_1766_));
 sky130_fd_sc_hd__and2_1 _6709_ (.A(_1765_),
    .B(_1766_),
    .X(_1767_));
 sky130_fd_sc_hd__xor2_1 _6710_ (.A(_1761_),
    .B(_1767_),
    .X(_1768_));
 sky130_fd_sc_hd__xor2_1 _6711_ (.A(_1530_),
    .B(_1582_),
    .X(_1769_));
 sky130_fd_sc_hd__xnor2_1 _6712_ (.A(_1765_),
    .B(_1769_),
    .Y(_1771_));
 sky130_fd_sc_hd__or2b_1 _6713_ (.A(_1768_),
    .B_N(_1771_),
    .X(_1772_));
 sky130_fd_sc_hd__or2_1 _6714_ (.A(_1653_),
    .B(_1772_),
    .X(_1773_));
 sky130_fd_sc_hd__xnor2_1 _6715_ (.A(_1702_),
    .B(_1732_),
    .Y(_1774_));
 sky130_fd_sc_hd__or2_1 _6716_ (.A(_0080_),
    .B(_1718_),
    .X(_1775_));
 sky130_fd_sc_hd__or2_1 _6717_ (.A(_0303_),
    .B(_1537_),
    .X(_1776_));
 sky130_fd_sc_hd__xnor2_1 _6718_ (.A(_1776_),
    .B(_1725_),
    .Y(_1777_));
 sky130_fd_sc_hd__or2b_1 _6719_ (.A(_1775_),
    .B_N(_1777_),
    .X(_1778_));
 sky130_fd_sc_hd__or2_1 _6720_ (.A(_1599_),
    .B(_1676_),
    .X(_1779_));
 sky130_fd_sc_hd__nor2_1 _6721_ (.A(_1400_),
    .B(_0548_),
    .Y(_1780_));
 sky130_fd_sc_hd__clkbuf_4 _6722_ (.A(_3868_),
    .X(_1782_));
 sky130_fd_sc_hd__and3_1 _6723_ (.A(_1353_),
    .B(_1354_),
    .C(_1782_),
    .X(_1783_));
 sky130_fd_sc_hd__or2_1 _6724_ (.A(_1383_),
    .B(_3703_),
    .X(_1784_));
 sky130_fd_sc_hd__xnor2_2 _6725_ (.A(_1783_),
    .B(_1784_),
    .Y(_1785_));
 sky130_fd_sc_hd__a2bb2oi_2 _6726_ (.A1_N(_1677_),
    .A2_N(_1779_),
    .B1(_1780_),
    .B2(_1785_),
    .Y(_1786_));
 sky130_fd_sc_hd__or2_1 _6727_ (.A(_1410_),
    .B(_1401_),
    .X(_1787_));
 sky130_fd_sc_hd__and3_1 _6728_ (.A(_1408_),
    .B(_1409_),
    .C(_0147_),
    .X(_1788_));
 sky130_fd_sc_hd__xnor2_1 _6729_ (.A(_1668_),
    .B(_1788_),
    .Y(_1789_));
 sky130_fd_sc_hd__nor2_1 _6730_ (.A(_1423_),
    .B(_1454_),
    .Y(_1790_));
 sky130_fd_sc_hd__nand2_1 _6731_ (.A(_1789_),
    .B(_1790_),
    .Y(_1791_));
 sky130_fd_sc_hd__o21ai_1 _6732_ (.A1(_1668_),
    .A2(_1787_),
    .B1(_1791_),
    .Y(_1793_));
 sky130_fd_sc_hd__nor2_1 _6733_ (.A(_1399_),
    .B(_1676_),
    .Y(_1794_));
 sky130_fd_sc_hd__xnor2_1 _6734_ (.A(_1794_),
    .B(_1679_),
    .Y(_1795_));
 sky130_fd_sc_hd__nor2_1 _6735_ (.A(_1793_),
    .B(_1795_),
    .Y(_1796_));
 sky130_fd_sc_hd__nand2_1 _6736_ (.A(_1793_),
    .B(_1795_),
    .Y(_1797_));
 sky130_fd_sc_hd__o21ai_2 _6737_ (.A1(_1786_),
    .A2(_1796_),
    .B1(_1797_),
    .Y(_1798_));
 sky130_fd_sc_hd__xor2_1 _6738_ (.A(_1710_),
    .B(_1719_),
    .X(_1799_));
 sky130_fd_sc_hd__xnor2_1 _6739_ (.A(_1798_),
    .B(_1799_),
    .Y(_1800_));
 sky130_fd_sc_hd__xor2_1 _6740_ (.A(_1778_),
    .B(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__xnor2_1 _6741_ (.A(_1675_),
    .B(_1689_),
    .Y(_1802_));
 sky130_fd_sc_hd__xnor2_1 _6742_ (.A(_1667_),
    .B(_1673_),
    .Y(_1804_));
 sky130_fd_sc_hd__xor2_1 _6743_ (.A(_1789_),
    .B(_1790_),
    .X(_1805_));
 sky130_fd_sc_hd__nor2_1 _6744_ (.A(_4232_),
    .B(_1664_),
    .Y(_1806_));
 sky130_fd_sc_hd__o21ba_1 _6745_ (.A1(_1428_),
    .A2(_1510_),
    .B1_N(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__a21o_1 _6746_ (.A1(_1665_),
    .A2(_1511_),
    .B1(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__o21ai_2 _6747_ (.A1(_1298_),
    .A2(_1299_),
    .B1(_1278_),
    .Y(_1809_));
 sky130_fd_sc_hd__and3_1 _6748_ (.A(_0218_),
    .B(_1300_),
    .C(_1809_),
    .X(_1810_));
 sky130_fd_sc_hd__nor2_1 _6749_ (.A(_1384_),
    .B(_1510_),
    .Y(_1811_));
 sky130_fd_sc_hd__and2_1 _6750_ (.A(_1300_),
    .B(_1809_),
    .X(_1812_));
 sky130_fd_sc_hd__clkbuf_2 _6751_ (.A(_1812_),
    .X(_1813_));
 sky130_fd_sc_hd__o2bb2a_1 _6752_ (.A1_N(_1813_),
    .A2_N(_0121_),
    .B1(_4228_),
    .B2(_1664_),
    .X(_1815_));
 sky130_fd_sc_hd__a21oi_1 _6753_ (.A1(_1806_),
    .A2(_1810_),
    .B1(_1815_),
    .Y(_1816_));
 sky130_fd_sc_hd__a22oi_2 _6754_ (.A1(_1806_),
    .A2(_1810_),
    .B1(_1811_),
    .B2(_1816_),
    .Y(_1817_));
 sky130_fd_sc_hd__nor2_1 _6755_ (.A(_1808_),
    .B(_1817_),
    .Y(_1818_));
 sky130_fd_sc_hd__and2_1 _6756_ (.A(_1808_),
    .B(_1817_),
    .X(_1819_));
 sky130_fd_sc_hd__nor2_1 _6757_ (.A(_1818_),
    .B(_1819_),
    .Y(_1820_));
 sky130_fd_sc_hd__a21oi_1 _6758_ (.A1(_1805_),
    .A2(_1820_),
    .B1(_1818_),
    .Y(_1821_));
 sky130_fd_sc_hd__xor2_1 _6759_ (.A(_1804_),
    .B(_1821_),
    .X(_1822_));
 sky130_fd_sc_hd__xor2_1 _6760_ (.A(_1793_),
    .B(_1795_),
    .X(_1823_));
 sky130_fd_sc_hd__xnor2_1 _6761_ (.A(_1786_),
    .B(_1823_),
    .Y(_1824_));
 sky130_fd_sc_hd__nor2_1 _6762_ (.A(_1804_),
    .B(_1821_),
    .Y(_1826_));
 sky130_fd_sc_hd__a21oi_1 _6763_ (.A1(_1822_),
    .A2(_1824_),
    .B1(_1826_),
    .Y(_1827_));
 sky130_fd_sc_hd__xor2_1 _6764_ (.A(_1802_),
    .B(_1827_),
    .X(_1828_));
 sky130_fd_sc_hd__nor2_1 _6765_ (.A(_1802_),
    .B(_1827_),
    .Y(_1829_));
 sky130_fd_sc_hd__a21o_1 _6766_ (.A1(_1801_),
    .A2(_1828_),
    .B1(_1829_),
    .X(_1830_));
 sky130_fd_sc_hd__or2b_1 _6767_ (.A(_1774_),
    .B_N(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__nand2_1 _6768_ (.A(_1798_),
    .B(_1799_),
    .Y(_1832_));
 sky130_fd_sc_hd__o21ai_1 _6769_ (.A1(_1778_),
    .A2(_1800_),
    .B1(_1832_),
    .Y(_1833_));
 sky130_fd_sc_hd__xnor2_1 _6770_ (.A(_1830_),
    .B(_1774_),
    .Y(_1834_));
 sky130_fd_sc_hd__nand2_1 _6771_ (.A(_1833_),
    .B(_1834_),
    .Y(_1835_));
 sky130_fd_sc_hd__xnor2_1 _6772_ (.A(_1750_),
    .B(_1751_),
    .Y(_1837_));
 sky130_fd_sc_hd__a21o_1 _6773_ (.A1(_1831_),
    .A2(_1835_),
    .B1(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__nand3_1 _6774_ (.A(_1831_),
    .B(_1835_),
    .C(_1837_),
    .Y(_1839_));
 sky130_fd_sc_hd__and2_1 _6775_ (.A(_1838_),
    .B(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__xnor2_1 _6776_ (.A(_1801_),
    .B(_1828_),
    .Y(_1841_));
 sky130_fd_sc_hd__or2_1 _6777_ (.A(_1420_),
    .B(_1718_),
    .X(_1842_));
 sky130_fd_sc_hd__or2_1 _6778_ (.A(_1776_),
    .B(_1842_),
    .X(_1843_));
 sky130_fd_sc_hd__or2_1 _6779_ (.A(_1383_),
    .B(_4126_),
    .X(_1844_));
 sky130_fd_sc_hd__or2_1 _6780_ (.A(_1779_),
    .B(_1844_),
    .X(_1845_));
 sky130_fd_sc_hd__nand2_1 _6781_ (.A(_0147_),
    .B(_1413_),
    .Y(_1846_));
 sky130_fd_sc_hd__and3_1 _6782_ (.A(_1408_),
    .B(_1409_),
    .C(_4089_),
    .X(_1848_));
 sky130_fd_sc_hd__xnor2_1 _6783_ (.A(_1846_),
    .B(_1848_),
    .Y(_1849_));
 sky130_fd_sc_hd__nand2_1 _6784_ (.A(_1413_),
    .B(_4089_),
    .Y(_1850_));
 sky130_fd_sc_hd__nor2_1 _6785_ (.A(_1787_),
    .B(_1850_),
    .Y(_1851_));
 sky130_fd_sc_hd__a31o_1 _6786_ (.A1(_1482_),
    .A2(_1782_),
    .A3(_1849_),
    .B1(_1851_),
    .X(_1852_));
 sky130_fd_sc_hd__or2_1 _6787_ (.A(_1399_),
    .B(_4126_),
    .X(_1853_));
 sky130_fd_sc_hd__xnor2_2 _6788_ (.A(_1853_),
    .B(_1785_),
    .Y(_1854_));
 sky130_fd_sc_hd__nor2_1 _6789_ (.A(_1852_),
    .B(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__nand2_1 _6790_ (.A(_1852_),
    .B(_1854_),
    .Y(_1856_));
 sky130_fd_sc_hd__o21ai_1 _6791_ (.A1(_1845_),
    .A2(_1855_),
    .B1(_1856_),
    .Y(_1857_));
 sky130_fd_sc_hd__xnor2_1 _6792_ (.A(_1775_),
    .B(_1777_),
    .Y(_1859_));
 sky130_fd_sc_hd__xor2_1 _6793_ (.A(_1857_),
    .B(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__xnor2_1 _6794_ (.A(_1843_),
    .B(_1860_),
    .Y(_1861_));
 sky130_fd_sc_hd__xnor2_1 _6795_ (.A(_1822_),
    .B(_1824_),
    .Y(_1862_));
 sky130_fd_sc_hd__xnor2_1 _6796_ (.A(_1805_),
    .B(_1820_),
    .Y(_1863_));
 sky130_fd_sc_hd__xnor2_1 _6797_ (.A(_1811_),
    .B(_1816_),
    .Y(_1864_));
 sky130_fd_sc_hd__nor2_1 _6798_ (.A(_3988_),
    .B(_1664_),
    .Y(_1865_));
 sky130_fd_sc_hd__nor2_1 _6799_ (.A(_1401_),
    .B(_1510_),
    .Y(_1866_));
 sky130_fd_sc_hd__xor2_1 _6800_ (.A(_1810_),
    .B(_1865_),
    .X(_1867_));
 sky130_fd_sc_hd__a22o_1 _6801_ (.A1(_1810_),
    .A2(_1865_),
    .B1(_1866_),
    .B2(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__and2b_1 _6802_ (.A_N(_1864_),
    .B(_1868_),
    .X(_1870_));
 sky130_fd_sc_hd__and2b_1 _6803_ (.A_N(_1868_),
    .B(_1864_),
    .X(_1871_));
 sky130_fd_sc_hd__nor2_1 _6804_ (.A(_1870_),
    .B(_1871_),
    .Y(_1872_));
 sky130_fd_sc_hd__or2_1 _6805_ (.A(_1422_),
    .B(_1456_),
    .X(_1873_));
 sky130_fd_sc_hd__xnor2_1 _6806_ (.A(_1873_),
    .B(_1849_),
    .Y(_1874_));
 sky130_fd_sc_hd__a21oi_1 _6807_ (.A1(_1872_),
    .A2(_1874_),
    .B1(_1870_),
    .Y(_1875_));
 sky130_fd_sc_hd__nor2_1 _6808_ (.A(_1863_),
    .B(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__and2_1 _6809_ (.A(_1863_),
    .B(_1875_),
    .X(_1877_));
 sky130_fd_sc_hd__nor2_1 _6810_ (.A(_1876_),
    .B(_1877_),
    .Y(_1878_));
 sky130_fd_sc_hd__xor2_1 _6811_ (.A(_1852_),
    .B(_1854_),
    .X(_1879_));
 sky130_fd_sc_hd__xnor2_1 _6812_ (.A(_1845_),
    .B(_1879_),
    .Y(_1881_));
 sky130_fd_sc_hd__a21o_1 _6813_ (.A1(_1878_),
    .A2(_1881_),
    .B1(_1876_),
    .X(_1882_));
 sky130_fd_sc_hd__xnor2_1 _6814_ (.A(_1862_),
    .B(_1882_),
    .Y(_1883_));
 sky130_fd_sc_hd__or2b_1 _6815_ (.A(_1862_),
    .B_N(_1882_),
    .X(_1884_));
 sky130_fd_sc_hd__a21boi_1 _6816_ (.A1(_1861_),
    .A2(_1883_),
    .B1_N(_1884_),
    .Y(_1885_));
 sky130_fd_sc_hd__or2_1 _6817_ (.A(_1841_),
    .B(_1885_),
    .X(_1886_));
 sky130_fd_sc_hd__nand2_1 _6818_ (.A(_1841_),
    .B(_1885_),
    .Y(_1887_));
 sky130_fd_sc_hd__nand2_1 _6819_ (.A(_1886_),
    .B(_1887_),
    .Y(_1888_));
 sky130_fd_sc_hd__or2b_1 _6820_ (.A(_1843_),
    .B_N(_1860_),
    .X(_1889_));
 sky130_fd_sc_hd__a21bo_1 _6821_ (.A1(_1857_),
    .A2(_1859_),
    .B1_N(_1889_),
    .X(_1890_));
 sky130_fd_sc_hd__or2b_1 _6822_ (.A(_1888_),
    .B_N(_1890_),
    .X(_1892_));
 sky130_fd_sc_hd__or2_1 _6823_ (.A(_1833_),
    .B(_1834_),
    .X(_1893_));
 sky130_fd_sc_hd__nand2_1 _6824_ (.A(_1835_),
    .B(_1893_),
    .Y(_1894_));
 sky130_fd_sc_hd__a21oi_2 _6825_ (.A1(_1886_),
    .A2(_1892_),
    .B1(_1894_),
    .Y(_1895_));
 sky130_fd_sc_hd__xnor2_1 _6826_ (.A(_1840_),
    .B(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__nand3_1 _6827_ (.A(_1746_),
    .B(_1752_),
    .C(_1760_),
    .Y(_1897_));
 sky130_fd_sc_hd__nand2_1 _6828_ (.A(_1761_),
    .B(_1897_),
    .Y(_1898_));
 sky130_fd_sc_hd__xnor2_1 _6829_ (.A(_1838_),
    .B(_1898_),
    .Y(_1899_));
 sky130_fd_sc_hd__nor2_1 _6830_ (.A(_1896_),
    .B(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__xor2_1 _6831_ (.A(_1890_),
    .B(_1888_),
    .X(_1901_));
 sky130_fd_sc_hd__xnor2_1 _6832_ (.A(_1861_),
    .B(_1883_),
    .Y(_1903_));
 sky130_fd_sc_hd__xnor2_1 _6833_ (.A(_1866_),
    .B(_1867_),
    .Y(_1904_));
 sky130_fd_sc_hd__and3_1 _6834_ (.A(_1300_),
    .B(_4153_),
    .C(_1809_),
    .X(_1905_));
 sky130_fd_sc_hd__nor2_1 _6835_ (.A(_1454_),
    .B(_1510_),
    .Y(_1906_));
 sky130_fd_sc_hd__nor2_1 _6836_ (.A(_3840_),
    .B(_1664_),
    .Y(_1907_));
 sky130_fd_sc_hd__a21oi_1 _6837_ (.A1(_4217_),
    .A2(_1813_),
    .B1(_1907_),
    .Y(_1908_));
 sky130_fd_sc_hd__a21oi_1 _6838_ (.A1(_1865_),
    .A2(_1905_),
    .B1(_1908_),
    .Y(_1909_));
 sky130_fd_sc_hd__a22o_1 _6839_ (.A1(_1865_),
    .A2(_1905_),
    .B1(_1906_),
    .B2(_1909_),
    .X(_1910_));
 sky130_fd_sc_hd__xnor2_1 _6840_ (.A(_1904_),
    .B(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__or2_1 _6841_ (.A(_1422_),
    .B(_3703_),
    .X(_1912_));
 sky130_fd_sc_hd__and3_1 _6842_ (.A(_1408_),
    .B(_1409_),
    .C(_1782_),
    .X(_1914_));
 sky130_fd_sc_hd__xnor2_1 _6843_ (.A(_1850_),
    .B(_1914_),
    .Y(_1915_));
 sky130_fd_sc_hd__xnor2_1 _6844_ (.A(_1912_),
    .B(_1915_),
    .Y(_1916_));
 sky130_fd_sc_hd__and2b_1 _6845_ (.A_N(_1904_),
    .B(_1910_),
    .X(_1917_));
 sky130_fd_sc_hd__a21o_1 _6846_ (.A1(_1911_),
    .A2(_1916_),
    .B1(_1917_),
    .X(_1918_));
 sky130_fd_sc_hd__xor2_1 _6847_ (.A(_1872_),
    .B(_1874_),
    .X(_1919_));
 sky130_fd_sc_hd__xor2_1 _6848_ (.A(_1918_),
    .B(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__and3_1 _6849_ (.A(_1414_),
    .B(_1782_),
    .C(_1848_),
    .X(_1921_));
 sky130_fd_sc_hd__a31oi_2 _6850_ (.A1(_1482_),
    .A2(_1531_),
    .A3(_1915_),
    .B1(_1921_),
    .Y(_1922_));
 sky130_fd_sc_hd__xnor2_1 _6851_ (.A(_1779_),
    .B(_1844_),
    .Y(_1923_));
 sky130_fd_sc_hd__xor2_1 _6852_ (.A(_1922_),
    .B(_1923_),
    .X(_1925_));
 sky130_fd_sc_hd__nand2_1 _6853_ (.A(_1918_),
    .B(_1919_),
    .Y(_1926_));
 sky130_fd_sc_hd__a21bo_1 _6854_ (.A1(_1920_),
    .A2(_1925_),
    .B1_N(_1926_),
    .X(_1927_));
 sky130_fd_sc_hd__xnor2_1 _6855_ (.A(_1878_),
    .B(_1881_),
    .Y(_1928_));
 sky130_fd_sc_hd__xnor2_1 _6856_ (.A(_1927_),
    .B(_1928_),
    .Y(_1929_));
 sky130_fd_sc_hd__or2_1 _6857_ (.A(_1420_),
    .B(_1538_),
    .X(_1930_));
 sky130_fd_sc_hd__or2_1 _6858_ (.A(_1428_),
    .B(_1718_),
    .X(_1931_));
 sky130_fd_sc_hd__or2_1 _6859_ (.A(_1930_),
    .B(_1931_),
    .X(_1932_));
 sky130_fd_sc_hd__or2_1 _6860_ (.A(_1922_),
    .B(_1923_),
    .X(_1933_));
 sky130_fd_sc_hd__o21ai_1 _6861_ (.A1(_0303_),
    .A2(_1718_),
    .B1(_1930_),
    .Y(_1934_));
 sky130_fd_sc_hd__and2_1 _6862_ (.A(_1843_),
    .B(_1934_),
    .X(_1936_));
 sky130_fd_sc_hd__xnor2_1 _6863_ (.A(_1933_),
    .B(_1936_),
    .Y(_1937_));
 sky130_fd_sc_hd__xnor2_1 _6864_ (.A(_1932_),
    .B(_1937_),
    .Y(_1938_));
 sky130_fd_sc_hd__and2b_1 _6865_ (.A_N(_1928_),
    .B(_1927_),
    .X(_1939_));
 sky130_fd_sc_hd__a21oi_1 _6866_ (.A1(_1929_),
    .A2(_1938_),
    .B1(_1939_),
    .Y(_1940_));
 sky130_fd_sc_hd__xnor2_1 _6867_ (.A(_1903_),
    .B(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hd__inv_2 _6868_ (.A(_1936_),
    .Y(_1942_));
 sky130_fd_sc_hd__or2b_1 _6869_ (.A(_1932_),
    .B_N(_1937_),
    .X(_1943_));
 sky130_fd_sc_hd__o21ai_1 _6870_ (.A1(_1933_),
    .A2(_1942_),
    .B1(_1943_),
    .Y(_1944_));
 sky130_fd_sc_hd__or2b_1 _6871_ (.A(_1941_),
    .B_N(_1944_),
    .X(_1945_));
 sky130_fd_sc_hd__o21ai_2 _6872_ (.A1(_1903_),
    .A2(_1940_),
    .B1(_1945_),
    .Y(_1947_));
 sky130_fd_sc_hd__and2b_1 _6873_ (.A_N(_1901_),
    .B(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__xor2_1 _6874_ (.A(_1947_),
    .B(_1901_),
    .X(_1949_));
 sky130_fd_sc_hd__nand2_2 _6875_ (.A(_1257_),
    .B(_1302_),
    .Y(_1950_));
 sky130_fd_sc_hd__and3_1 _6876_ (.A(_1711_),
    .B(_0121_),
    .C(_1950_),
    .X(_1951_));
 sky130_fd_sc_hd__xor2_1 _6877_ (.A(_1944_),
    .B(_1941_),
    .X(_1952_));
 sky130_fd_sc_hd__nor2_1 _6878_ (.A(_1428_),
    .B(_1538_),
    .Y(_1953_));
 sky130_fd_sc_hd__nor2_1 _6879_ (.A(_1384_),
    .B(_1718_),
    .Y(_1954_));
 sky130_fd_sc_hd__nand2_1 _6880_ (.A(_1413_),
    .B(_1782_),
    .Y(_1955_));
 sky130_fd_sc_hd__nand3_1 _6881_ (.A(_1408_),
    .B(_1409_),
    .C(_1531_),
    .Y(_1956_));
 sky130_fd_sc_hd__xnor2_1 _6882_ (.A(_1955_),
    .B(_1956_),
    .Y(_1958_));
 sky130_fd_sc_hd__or2_1 _6883_ (.A(_1955_),
    .B(_1956_),
    .X(_1959_));
 sky130_fd_sc_hd__o31a_1 _6884_ (.A1(_1423_),
    .A2(_0548_),
    .A3(_1958_),
    .B1(_1959_),
    .X(_1960_));
 sky130_fd_sc_hd__or3_1 _6885_ (.A(_1599_),
    .B(_0548_),
    .C(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__xnor2_1 _6886_ (.A(_1842_),
    .B(_1953_),
    .Y(_1962_));
 sky130_fd_sc_hd__xnor2_1 _6887_ (.A(_1961_),
    .B(_1962_),
    .Y(_1963_));
 sky130_fd_sc_hd__and2b_1 _6888_ (.A_N(_1961_),
    .B(_1962_),
    .X(_1964_));
 sky130_fd_sc_hd__a31o_1 _6889_ (.A1(_1953_),
    .A2(_1954_),
    .A3(_1963_),
    .B1(_1964_),
    .X(_1965_));
 sky130_fd_sc_hd__xnor2_1 _6890_ (.A(_1906_),
    .B(_1909_),
    .Y(_1966_));
 sky130_fd_sc_hd__or2_1 _6891_ (.A(_1509_),
    .B(_3930_),
    .X(_1967_));
 sky130_fd_sc_hd__and3_1 _6892_ (.A(_1300_),
    .B(_1355_),
    .C(_1809_),
    .X(_1969_));
 sky130_fd_sc_hd__nor2_1 _6893_ (.A(_1665_),
    .B(_1905_),
    .Y(_1970_));
 sky130_fd_sc_hd__a21o_1 _6894_ (.A1(_1907_),
    .A2(_1969_),
    .B1(_1970_),
    .X(_1971_));
 sky130_fd_sc_hd__o2bb2ai_1 _6895_ (.A1_N(_1665_),
    .A2_N(_1905_),
    .B1(_1967_),
    .B2(_1971_),
    .Y(_1972_));
 sky130_fd_sc_hd__and2b_1 _6896_ (.A_N(_1966_),
    .B(_1972_),
    .X(_1973_));
 sky130_fd_sc_hd__and2b_1 _6897_ (.A_N(_1972_),
    .B(_1966_),
    .X(_1974_));
 sky130_fd_sc_hd__nor2_1 _6898_ (.A(_1973_),
    .B(_1974_),
    .Y(_1975_));
 sky130_fd_sc_hd__nor2_1 _6899_ (.A(_1422_),
    .B(_4126_),
    .Y(_1976_));
 sky130_fd_sc_hd__xnor2_1 _6900_ (.A(_1976_),
    .B(_1958_),
    .Y(_1977_));
 sky130_fd_sc_hd__a21oi_1 _6901_ (.A1(_1975_),
    .A2(_1977_),
    .B1(_1973_),
    .Y(_1978_));
 sky130_fd_sc_hd__xnor2_1 _6902_ (.A(_1911_),
    .B(_1916_),
    .Y(_1980_));
 sky130_fd_sc_hd__xor2_1 _6903_ (.A(_1978_),
    .B(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__nor2_1 _6904_ (.A(_1599_),
    .B(_0548_),
    .Y(_1982_));
 sky130_fd_sc_hd__xnor2_1 _6905_ (.A(_1982_),
    .B(_1960_),
    .Y(_1983_));
 sky130_fd_sc_hd__nor2_1 _6906_ (.A(_1978_),
    .B(_1980_),
    .Y(_1984_));
 sky130_fd_sc_hd__a21o_1 _6907_ (.A1(_1981_),
    .A2(_1983_),
    .B1(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__xor2_1 _6908_ (.A(_1920_),
    .B(_1925_),
    .X(_1986_));
 sky130_fd_sc_hd__xor2_1 _6909_ (.A(_1985_),
    .B(_1986_),
    .X(_1987_));
 sky130_fd_sc_hd__nand2_1 _6910_ (.A(_1953_),
    .B(_1954_),
    .Y(_1988_));
 sky130_fd_sc_hd__xnor2_1 _6911_ (.A(_1988_),
    .B(_1963_),
    .Y(_1989_));
 sky130_fd_sc_hd__nand2_1 _6912_ (.A(_1985_),
    .B(_1986_),
    .Y(_1991_));
 sky130_fd_sc_hd__a21bo_1 _6913_ (.A1(_1987_),
    .A2(_1989_),
    .B1_N(_1991_),
    .X(_1992_));
 sky130_fd_sc_hd__xnor2_1 _6914_ (.A(_1929_),
    .B(_1938_),
    .Y(_1993_));
 sky130_fd_sc_hd__xnor2_1 _6915_ (.A(_1992_),
    .B(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__or2b_1 _6916_ (.A(_1993_),
    .B_N(_1992_),
    .X(_1995_));
 sky130_fd_sc_hd__a21boi_1 _6917_ (.A1(_1965_),
    .A2(_1994_),
    .B1_N(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__xor2_1 _6918_ (.A(_1952_),
    .B(_1996_),
    .X(_1997_));
 sky130_fd_sc_hd__nor2_1 _6919_ (.A(_1952_),
    .B(_1996_),
    .Y(_1998_));
 sky130_fd_sc_hd__a21o_1 _6920_ (.A1(_1951_),
    .A2(_1997_),
    .B1(_1998_),
    .X(_1999_));
 sky130_fd_sc_hd__and2b_1 _6921_ (.A_N(_1949_),
    .B(_1999_),
    .X(_2000_));
 sky130_fd_sc_hd__and3_1 _6922_ (.A(_1886_),
    .B(_1892_),
    .C(_1894_),
    .X(_2002_));
 sky130_fd_sc_hd__nor2_2 _6923_ (.A(_1895_),
    .B(_2002_),
    .Y(_2003_));
 sky130_fd_sc_hd__o21a_1 _6924_ (.A1(_1948_),
    .A2(_2000_),
    .B1(_2003_),
    .X(_2004_));
 sky130_fd_sc_hd__nand2_1 _6925_ (.A(_1840_),
    .B(_1895_),
    .Y(_2005_));
 sky130_fd_sc_hd__a21oi_1 _6926_ (.A1(_1838_),
    .A2(_2005_),
    .B1(_1898_),
    .Y(_2006_));
 sky130_fd_sc_hd__a21o_1 _6927_ (.A1(_1900_),
    .A2(_2004_),
    .B1(_2006_),
    .X(_2007_));
 sky130_fd_sc_hd__or2b_1 _6928_ (.A(_1773_),
    .B_N(_2007_),
    .X(_2008_));
 sky130_fd_sc_hd__and3_1 _6929_ (.A(_0218_),
    .B(_1711_),
    .C(_1950_),
    .X(_2009_));
 sky130_fd_sc_hd__and3_1 _6930_ (.A(_1408_),
    .B(_1409_),
    .C(_3804_),
    .X(_2010_));
 sky130_fd_sc_hd__and3_1 _6931_ (.A(_1414_),
    .B(_1531_),
    .C(_2010_),
    .X(_2011_));
 sky130_fd_sc_hd__xnor2_1 _6932_ (.A(_1967_),
    .B(_1971_),
    .Y(_2013_));
 sky130_fd_sc_hd__and3_1 _6933_ (.A(_1300_),
    .B(_3986_),
    .C(_1809_),
    .X(_2014_));
 sky130_fd_sc_hd__or2_1 _6934_ (.A(_3615_),
    .B(_1663_),
    .X(_2015_));
 sky130_fd_sc_hd__xnor2_1 _6935_ (.A(_1969_),
    .B(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__or3b_1 _6936_ (.A(_1509_),
    .B(_3703_),
    .C_N(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__a21bo_1 _6937_ (.A1(_1665_),
    .A2(_2014_),
    .B1_N(_2017_),
    .X(_2018_));
 sky130_fd_sc_hd__xnor2_1 _6938_ (.A(_2013_),
    .B(_2018_),
    .Y(_2019_));
 sky130_fd_sc_hd__nand2_1 _6939_ (.A(_1414_),
    .B(_1531_),
    .Y(_2020_));
 sky130_fd_sc_hd__xnor2_1 _6940_ (.A(_2020_),
    .B(_2010_),
    .Y(_2021_));
 sky130_fd_sc_hd__and2b_1 _6941_ (.A_N(_2013_),
    .B(_2018_),
    .X(_2022_));
 sky130_fd_sc_hd__a21o_1 _6942_ (.A1(_2019_),
    .A2(_2021_),
    .B1(_2022_),
    .X(_2024_));
 sky130_fd_sc_hd__xor2_1 _6943_ (.A(_1975_),
    .B(_1977_),
    .X(_2025_));
 sky130_fd_sc_hd__xor2_1 _6944_ (.A(_2024_),
    .B(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__and2_1 _6945_ (.A(_2024_),
    .B(_2025_),
    .X(_2027_));
 sky130_fd_sc_hd__a21oi_1 _6946_ (.A1(_2011_),
    .A2(_2026_),
    .B1(_2027_),
    .Y(_2028_));
 sky130_fd_sc_hd__xnor2_1 _6947_ (.A(_1981_),
    .B(_1983_),
    .Y(_2029_));
 sky130_fd_sc_hd__xor2_1 _6948_ (.A(_2028_),
    .B(_2029_),
    .X(_2030_));
 sky130_fd_sc_hd__nor2_1 _6949_ (.A(_1384_),
    .B(_1538_),
    .Y(_2031_));
 sky130_fd_sc_hd__nor2_1 _6950_ (.A(_1401_),
    .B(_1718_),
    .Y(_2032_));
 sky130_fd_sc_hd__and3_1 _6951_ (.A(_1931_),
    .B(_2031_),
    .C(_2032_),
    .X(_2033_));
 sky130_fd_sc_hd__o21ai_1 _6952_ (.A1(_1384_),
    .A2(_1538_),
    .B1(_1931_),
    .Y(_2035_));
 sky130_fd_sc_hd__nand2_1 _6953_ (.A(_2031_),
    .B(_2032_),
    .Y(_2036_));
 sky130_fd_sc_hd__a21boi_1 _6954_ (.A1(_1988_),
    .A2(_2035_),
    .B1_N(_2036_),
    .Y(_2037_));
 sky130_fd_sc_hd__nor2_1 _6955_ (.A(_2033_),
    .B(_2037_),
    .Y(_2038_));
 sky130_fd_sc_hd__nor2_1 _6956_ (.A(_2028_),
    .B(_2029_),
    .Y(_2039_));
 sky130_fd_sc_hd__a21o_1 _6957_ (.A1(_2030_),
    .A2(_2038_),
    .B1(_2039_),
    .X(_2040_));
 sky130_fd_sc_hd__xor2_1 _6958_ (.A(_1987_),
    .B(_1989_),
    .X(_2041_));
 sky130_fd_sc_hd__xor2_1 _6959_ (.A(_2040_),
    .B(_2041_),
    .X(_2042_));
 sky130_fd_sc_hd__a22o_1 _6960_ (.A1(_2040_),
    .A2(_2041_),
    .B1(_2042_),
    .B2(_2033_),
    .X(_2043_));
 sky130_fd_sc_hd__xnor2_1 _6961_ (.A(_1965_),
    .B(_1994_),
    .Y(_2044_));
 sky130_fd_sc_hd__xnor2_1 _6962_ (.A(_2043_),
    .B(_2044_),
    .Y(_2046_));
 sky130_fd_sc_hd__xnor2_1 _6963_ (.A(_2009_),
    .B(_2046_),
    .Y(_2047_));
 sky130_fd_sc_hd__xnor2_1 _6964_ (.A(_2019_),
    .B(_2021_),
    .Y(_2048_));
 sky130_fd_sc_hd__o21bai_1 _6965_ (.A1(_1510_),
    .A2(_3703_),
    .B1_N(_2016_),
    .Y(_2049_));
 sky130_fd_sc_hd__o21ba_1 _6966_ (.A1(_3817_),
    .A2(_1663_),
    .B1_N(_2014_),
    .X(_2050_));
 sky130_fd_sc_hd__nand2_1 _6967_ (.A(_0147_),
    .B(_1813_),
    .Y(_2051_));
 sky130_fd_sc_hd__or2_1 _6968_ (.A(_2015_),
    .B(_2051_),
    .X(_2052_));
 sky130_fd_sc_hd__o31ai_1 _6969_ (.A1(_1510_),
    .A2(_4126_),
    .A3(_2050_),
    .B1(_2052_),
    .Y(_2053_));
 sky130_fd_sc_hd__nand3_1 _6970_ (.A(_2017_),
    .B(_2049_),
    .C(_2053_),
    .Y(_2054_));
 sky130_fd_sc_hd__and2_1 _6971_ (.A(_1414_),
    .B(_3804_),
    .X(_2055_));
 sky130_fd_sc_hd__a21o_1 _6972_ (.A1(_2017_),
    .A2(_2049_),
    .B1(_2053_),
    .X(_2057_));
 sky130_fd_sc_hd__nand3_1 _6973_ (.A(_2055_),
    .B(_2054_),
    .C(_2057_),
    .Y(_2058_));
 sky130_fd_sc_hd__nand2_1 _6974_ (.A(_2054_),
    .B(_2058_),
    .Y(_2059_));
 sky130_fd_sc_hd__or2b_1 _6975_ (.A(_2048_),
    .B_N(_2059_),
    .X(_2060_));
 sky130_fd_sc_hd__xor2_1 _6976_ (.A(_2011_),
    .B(_2026_),
    .X(_2061_));
 sky130_fd_sc_hd__xor2_1 _6977_ (.A(_2060_),
    .B(_2061_),
    .X(_2062_));
 sky130_fd_sc_hd__or2_1 _6978_ (.A(_1454_),
    .B(_1718_),
    .X(_2063_));
 sky130_fd_sc_hd__or3_1 _6979_ (.A(_1401_),
    .B(_1537_),
    .C(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__nor2_1 _6980_ (.A(_1401_),
    .B(_1538_),
    .Y(_2065_));
 sky130_fd_sc_hd__o21ai_1 _6981_ (.A1(_1954_),
    .A2(_2065_),
    .B1(_2036_),
    .Y(_2066_));
 sky130_fd_sc_hd__and2b_1 _6982_ (.A_N(_2064_),
    .B(_2036_),
    .X(_2068_));
 sky130_fd_sc_hd__a21oi_1 _6983_ (.A1(_2064_),
    .A2(_2066_),
    .B1(_2068_),
    .Y(_2069_));
 sky130_fd_sc_hd__inv_2 _6984_ (.A(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__or2b_1 _6985_ (.A(_2060_),
    .B_N(_2061_),
    .X(_2071_));
 sky130_fd_sc_hd__o21a_1 _6986_ (.A1(_2062_),
    .A2(_2070_),
    .B1(_2071_),
    .X(_2072_));
 sky130_fd_sc_hd__xnor2_1 _6987_ (.A(_2030_),
    .B(_2038_),
    .Y(_2073_));
 sky130_fd_sc_hd__xor2_1 _6988_ (.A(_2072_),
    .B(_2073_),
    .X(_2074_));
 sky130_fd_sc_hd__a2bb2o_1 _6989_ (.A1_N(_2072_),
    .A2_N(_2073_),
    .B1(_2074_),
    .B2(_2068_),
    .X(_2075_));
 sky130_fd_sc_hd__xor2_1 _6990_ (.A(_2033_),
    .B(_2042_),
    .X(_2076_));
 sky130_fd_sc_hd__and2_1 _6991_ (.A(_1711_),
    .B(_1950_),
    .X(_2077_));
 sky130_fd_sc_hd__buf_2 _6992_ (.A(_2077_),
    .X(_2079_));
 sky130_fd_sc_hd__xor2_1 _6993_ (.A(_2075_),
    .B(_2076_),
    .X(_2080_));
 sky130_fd_sc_hd__and3_1 _6994_ (.A(_4217_),
    .B(_2079_),
    .C(_2080_),
    .X(_2081_));
 sky130_fd_sc_hd__a21oi_1 _6995_ (.A1(_2075_),
    .A2(_2076_),
    .B1(_2081_),
    .Y(_2082_));
 sky130_fd_sc_hd__nor2_1 _6996_ (.A(_2047_),
    .B(_2082_),
    .Y(_2083_));
 sky130_fd_sc_hd__and2_1 _6997_ (.A(_2047_),
    .B(_2082_),
    .X(_2084_));
 sky130_fd_sc_hd__nor2_2 _6998_ (.A(_2083_),
    .B(_2084_),
    .Y(_2085_));
 sky130_fd_sc_hd__or2_1 _6999_ (.A(_1456_),
    .B(_1717_),
    .X(_2086_));
 sky130_fd_sc_hd__nor2_1 _7000_ (.A(_1454_),
    .B(_1537_),
    .Y(_2087_));
 sky130_fd_sc_hd__and3b_1 _7001_ (.A_N(_2086_),
    .B(_2064_),
    .C(_2087_),
    .X(_2088_));
 sky130_fd_sc_hd__xor2_1 _7002_ (.A(_2059_),
    .B(_2048_),
    .X(_2090_));
 sky130_fd_sc_hd__a21o_1 _7003_ (.A1(_2054_),
    .A2(_2057_),
    .B1(_2055_),
    .X(_2091_));
 sky130_fd_sc_hd__or2_1 _7004_ (.A(_1509_),
    .B(_4126_),
    .X(_2092_));
 sky130_fd_sc_hd__o21ba_1 _7005_ (.A1(_2015_),
    .A2(_2051_),
    .B1_N(_2050_),
    .X(_2093_));
 sky130_fd_sc_hd__xnor2_1 _7006_ (.A(_2092_),
    .B(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hd__or2_1 _7007_ (.A(_1454_),
    .B(_1664_),
    .X(_2095_));
 sky130_fd_sc_hd__nor2_1 _7008_ (.A(_2051_),
    .B(_2095_),
    .Y(_2096_));
 sky130_fd_sc_hd__and2_1 _7009_ (.A(_2094_),
    .B(_2096_),
    .X(_2097_));
 sky130_fd_sc_hd__nand3_2 _7010_ (.A(_2058_),
    .B(_2091_),
    .C(_2097_),
    .Y(_2098_));
 sky130_fd_sc_hd__xor2_1 _7011_ (.A(_2090_),
    .B(_2098_),
    .X(_2099_));
 sky130_fd_sc_hd__inv_2 _7012_ (.A(_2088_),
    .Y(_2101_));
 sky130_fd_sc_hd__or4_1 _7013_ (.A(_1401_),
    .B(_1782_),
    .C(_1538_),
    .D(_2063_),
    .X(_2102_));
 sky130_fd_sc_hd__o211a_1 _7014_ (.A1(_2032_),
    .A2(_2087_),
    .B1(_2101_),
    .C1(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__nand2_1 _7015_ (.A(_2099_),
    .B(_2103_),
    .Y(_2104_));
 sky130_fd_sc_hd__o21ai_1 _7016_ (.A1(_2090_),
    .A2(_2098_),
    .B1(_2104_),
    .Y(_2105_));
 sky130_fd_sc_hd__xnor2_1 _7017_ (.A(_2062_),
    .B(_2070_),
    .Y(_2106_));
 sky130_fd_sc_hd__xnor2_1 _7018_ (.A(_2105_),
    .B(_2106_),
    .Y(_2107_));
 sky130_fd_sc_hd__or2b_1 _7019_ (.A(_2106_),
    .B_N(_2105_),
    .X(_2108_));
 sky130_fd_sc_hd__a21boi_1 _7020_ (.A1(_2088_),
    .A2(_2107_),
    .B1_N(_2108_),
    .Y(_2109_));
 sky130_fd_sc_hd__xnor2_1 _7021_ (.A(_2068_),
    .B(_2074_),
    .Y(_2110_));
 sky130_fd_sc_hd__or2_1 _7022_ (.A(_2109_),
    .B(_2110_),
    .X(_2112_));
 sky130_fd_sc_hd__nand2_1 _7023_ (.A(_4153_),
    .B(_2079_),
    .Y(_2113_));
 sky130_fd_sc_hd__xor2_1 _7024_ (.A(_2109_),
    .B(_2110_),
    .X(_2114_));
 sky130_fd_sc_hd__or2b_1 _7025_ (.A(_2113_),
    .B_N(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__nand2_1 _7026_ (.A(_4217_),
    .B(_2079_),
    .Y(_2116_));
 sky130_fd_sc_hd__xor2_1 _7027_ (.A(_2116_),
    .B(_2080_),
    .X(_2117_));
 sky130_fd_sc_hd__a21o_1 _7028_ (.A1(_2112_),
    .A2(_2115_),
    .B1(_2117_),
    .X(_2118_));
 sky130_fd_sc_hd__and3_1 _7029_ (.A(_2112_),
    .B(_2115_),
    .C(_2117_),
    .X(_2119_));
 sky130_fd_sc_hd__inv_2 _7030_ (.A(_2119_),
    .Y(_2120_));
 sky130_fd_sc_hd__xor2_1 _7031_ (.A(_2113_),
    .B(_2114_),
    .X(_2121_));
 sky130_fd_sc_hd__and3_1 _7032_ (.A(_1711_),
    .B(_1355_),
    .C(_1950_),
    .X(_2123_));
 sky130_fd_sc_hd__a21o_1 _7033_ (.A1(_2058_),
    .A2(_2091_),
    .B1(_2097_),
    .X(_2124_));
 sky130_fd_sc_hd__nand2_1 _7034_ (.A(_1782_),
    .B(_1813_),
    .Y(_2125_));
 sky130_fd_sc_hd__or2_1 _7035_ (.A(_2095_),
    .B(_2125_),
    .X(_2126_));
 sky130_fd_sc_hd__and2_1 _7036_ (.A(_2051_),
    .B(_2095_),
    .X(_2127_));
 sky130_fd_sc_hd__or2_1 _7037_ (.A(_2096_),
    .B(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__xnor2_1 _7038_ (.A(_2094_),
    .B(_2096_),
    .Y(_2129_));
 sky130_fd_sc_hd__nor3_1 _7039_ (.A(_2126_),
    .B(_2128_),
    .C(_2129_),
    .Y(_2130_));
 sky130_fd_sc_hd__nand3_1 _7040_ (.A(_2098_),
    .B(_2124_),
    .C(_2130_),
    .Y(_2131_));
 sky130_fd_sc_hd__a21o_1 _7041_ (.A1(_2098_),
    .A2(_2124_),
    .B1(_2130_),
    .X(_2132_));
 sky130_fd_sc_hd__or4_1 _7042_ (.A(_4089_),
    .B(_1676_),
    .C(_1537_),
    .D(_2086_),
    .X(_2134_));
 sky130_fd_sc_hd__o21ai_1 _7043_ (.A1(_1456_),
    .A2(_1537_),
    .B1(_2063_),
    .Y(_2135_));
 sky130_fd_sc_hd__or4_1 _7044_ (.A(_1454_),
    .B(_1531_),
    .C(_1537_),
    .D(_2086_),
    .X(_2136_));
 sky130_fd_sc_hd__and3_1 _7045_ (.A(_2134_),
    .B(_2135_),
    .C(_2136_),
    .X(_2137_));
 sky130_fd_sc_hd__and3_1 _7046_ (.A(_2131_),
    .B(_2132_),
    .C(_2137_),
    .X(_2138_));
 sky130_fd_sc_hd__a31o_1 _7047_ (.A1(_2098_),
    .A2(_2124_),
    .A3(_2130_),
    .B1(_2138_),
    .X(_2139_));
 sky130_fd_sc_hd__or2_1 _7048_ (.A(_2099_),
    .B(_2103_),
    .X(_2140_));
 sky130_fd_sc_hd__nand2_1 _7049_ (.A(_2104_),
    .B(_2140_),
    .Y(_2141_));
 sky130_fd_sc_hd__xnor2_1 _7050_ (.A(_2139_),
    .B(_2141_),
    .Y(_2142_));
 sky130_fd_sc_hd__nor4_1 _7051_ (.A(_4089_),
    .B(_1676_),
    .C(_1538_),
    .D(_2086_),
    .Y(_2143_));
 sky130_fd_sc_hd__a32o_1 _7052_ (.A1(_2104_),
    .A2(_2139_),
    .A3(_2140_),
    .B1(_2142_),
    .B2(_2143_),
    .X(_2145_));
 sky130_fd_sc_hd__xnor2_1 _7053_ (.A(_2088_),
    .B(_2107_),
    .Y(_2146_));
 sky130_fd_sc_hd__xnor2_1 _7054_ (.A(_2145_),
    .B(_2146_),
    .Y(_2147_));
 sky130_fd_sc_hd__and2b_1 _7055_ (.A_N(_2146_),
    .B(_2145_),
    .X(_2148_));
 sky130_fd_sc_hd__a21oi_1 _7056_ (.A1(_2123_),
    .A2(_2147_),
    .B1(_2148_),
    .Y(_2149_));
 sky130_fd_sc_hd__xnor2_1 _7057_ (.A(_2121_),
    .B(_2149_),
    .Y(_2150_));
 sky130_fd_sc_hd__inv_2 _7058_ (.A(_2150_),
    .Y(_2151_));
 sky130_fd_sc_hd__xnor2_1 _7059_ (.A(_2123_),
    .B(_2147_),
    .Y(_2152_));
 sky130_fd_sc_hd__xor2_1 _7060_ (.A(_2134_),
    .B(_2142_),
    .X(_2153_));
 sky130_fd_sc_hd__a21oi_1 _7061_ (.A1(_2131_),
    .A2(_2132_),
    .B1(_2137_),
    .Y(_2154_));
 sky130_fd_sc_hd__or2_1 _7062_ (.A(_1664_),
    .B(_1456_),
    .X(_2156_));
 sky130_fd_sc_hd__nand2_1 _7063_ (.A(_1531_),
    .B(_1813_),
    .Y(_2157_));
 sky130_fd_sc_hd__nor2_1 _7064_ (.A(_2156_),
    .B(_2157_),
    .Y(_2158_));
 sky130_fd_sc_hd__nand2_1 _7065_ (.A(_1454_),
    .B(_2158_),
    .Y(_2159_));
 sky130_fd_sc_hd__nor2_1 _7066_ (.A(_4126_),
    .B(_1718_),
    .Y(_2160_));
 sky130_fd_sc_hd__or4_1 _7067_ (.A(_1676_),
    .B(_1537_),
    .C(_2086_),
    .D(_2160_),
    .X(_2161_));
 sky130_fd_sc_hd__o31ai_1 _7068_ (.A1(_1676_),
    .A2(_1537_),
    .A3(_2160_),
    .B1(_2086_),
    .Y(_2162_));
 sky130_fd_sc_hd__nand2_1 _7069_ (.A(_2161_),
    .B(_2162_),
    .Y(_2163_));
 sky130_fd_sc_hd__o21a_1 _7070_ (.A1(_2156_),
    .A2(_2157_),
    .B1(_2126_),
    .X(_2164_));
 sky130_fd_sc_hd__nor2_1 _7071_ (.A(_2128_),
    .B(_2164_),
    .Y(_2165_));
 sky130_fd_sc_hd__xnor2_1 _7072_ (.A(_2129_),
    .B(_2165_),
    .Y(_2167_));
 sky130_fd_sc_hd__or2b_1 _7073_ (.A(_2163_),
    .B_N(_2167_),
    .X(_2168_));
 sky130_fd_sc_hd__o31a_1 _7074_ (.A1(_2128_),
    .A2(_2129_),
    .A3(_2159_),
    .B1(_2168_),
    .X(_2169_));
 sky130_fd_sc_hd__or3_1 _7075_ (.A(_2138_),
    .B(_2154_),
    .C(_2169_),
    .X(_2170_));
 sky130_fd_sc_hd__nor2_1 _7076_ (.A(_1676_),
    .B(_1718_),
    .Y(_2171_));
 sky130_fd_sc_hd__o211a_1 _7077_ (.A1(_1456_),
    .A2(_1538_),
    .B1(_1705_),
    .C1(_2171_),
    .X(_2172_));
 sky130_fd_sc_hd__o21ai_1 _7078_ (.A1(_2138_),
    .A2(_2154_),
    .B1(_2169_),
    .Y(_2173_));
 sky130_fd_sc_hd__nand3_1 _7079_ (.A(_2172_),
    .B(_2170_),
    .C(_2173_),
    .Y(_2174_));
 sky130_fd_sc_hd__and2_1 _7080_ (.A(_2170_),
    .B(_2174_),
    .X(_2175_));
 sky130_fd_sc_hd__nand2_1 _7081_ (.A(_3986_),
    .B(_2079_),
    .Y(_2176_));
 sky130_fd_sc_hd__xor2_1 _7082_ (.A(_2153_),
    .B(_2175_),
    .X(_2178_));
 sky130_fd_sc_hd__or2b_1 _7083_ (.A(_2176_),
    .B_N(_2178_),
    .X(_2179_));
 sky130_fd_sc_hd__o21a_1 _7084_ (.A1(_2153_),
    .A2(_2175_),
    .B1(_2179_),
    .X(_2180_));
 sky130_fd_sc_hd__nand2_1 _7085_ (.A(_2152_),
    .B(_2180_),
    .Y(_2181_));
 sky130_fd_sc_hd__xor2_1 _7086_ (.A(_2176_),
    .B(_2178_),
    .X(_2182_));
 sky130_fd_sc_hd__a21o_1 _7087_ (.A1(_2170_),
    .A2(_2173_),
    .B1(_2172_),
    .X(_2183_));
 sky130_fd_sc_hd__xor2_1 _7088_ (.A(_2163_),
    .B(_2167_),
    .X(_2184_));
 sky130_fd_sc_hd__or4_1 _7089_ (.A(_1664_),
    .B(_1782_),
    .C(_4126_),
    .D(_2157_),
    .X(_2185_));
 sky130_fd_sc_hd__a21boi_1 _7090_ (.A1(_4089_),
    .A2(_1813_),
    .B1_N(_2156_),
    .Y(_2186_));
 sky130_fd_sc_hd__a21oi_1 _7091_ (.A1(_4089_),
    .A2(_2158_),
    .B1(_2164_),
    .Y(_2187_));
 sky130_fd_sc_hd__or3_1 _7092_ (.A(_2185_),
    .B(_2186_),
    .C(_2187_),
    .X(_2189_));
 sky130_fd_sc_hd__and2_1 _7093_ (.A(_2128_),
    .B(_2164_),
    .X(_2190_));
 sky130_fd_sc_hd__or2_1 _7094_ (.A(_2165_),
    .B(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__xor2_1 _7095_ (.A(_2189_),
    .B(_2191_),
    .X(_2192_));
 sky130_fd_sc_hd__xnor2_1 _7096_ (.A(_1703_),
    .B(_2171_),
    .Y(_2193_));
 sky130_fd_sc_hd__nor2_1 _7097_ (.A(_2189_),
    .B(_2191_),
    .Y(_2194_));
 sky130_fd_sc_hd__a21oi_1 _7098_ (.A1(_2192_),
    .A2(_2193_),
    .B1(_2194_),
    .Y(_2195_));
 sky130_fd_sc_hd__nor2_1 _7099_ (.A(_2184_),
    .B(_2195_),
    .Y(_2196_));
 sky130_fd_sc_hd__nand3_1 _7100_ (.A(_2174_),
    .B(_2183_),
    .C(_2196_),
    .Y(_2197_));
 sky130_fd_sc_hd__and3_1 _7101_ (.A(_2174_),
    .B(_2183_),
    .C(_2196_),
    .X(_2198_));
 sky130_fd_sc_hd__nand2_1 _7102_ (.A(_0147_),
    .B(_2079_),
    .Y(_2200_));
 sky130_fd_sc_hd__a21oi_1 _7103_ (.A1(_2174_),
    .A2(_2183_),
    .B1(_2196_),
    .Y(_2201_));
 sky130_fd_sc_hd__or3_1 _7104_ (.A(_2198_),
    .B(_2200_),
    .C(_2201_),
    .X(_2202_));
 sky130_fd_sc_hd__nand3_1 _7105_ (.A(_2182_),
    .B(_2197_),
    .C(_2202_),
    .Y(_2203_));
 sky130_fd_sc_hd__o21ai_1 _7106_ (.A1(_2198_),
    .A2(_2201_),
    .B1(_2200_),
    .Y(_2204_));
 sky130_fd_sc_hd__and2_1 _7107_ (.A(_2184_),
    .B(_2195_),
    .X(_2205_));
 sky130_fd_sc_hd__or2_1 _7108_ (.A(_2196_),
    .B(_2205_),
    .X(_2206_));
 sky130_fd_sc_hd__xor2_1 _7109_ (.A(_2192_),
    .B(_2193_),
    .X(_2207_));
 sky130_fd_sc_hd__o21ai_1 _7110_ (.A1(_2186_),
    .A2(_2187_),
    .B1(_2185_),
    .Y(_2208_));
 sky130_fd_sc_hd__and2_1 _7111_ (.A(_2189_),
    .B(_2208_),
    .X(_2209_));
 sky130_fd_sc_hd__and2_1 _7112_ (.A(_2160_),
    .B(_2209_),
    .X(_2211_));
 sky130_fd_sc_hd__nand2_1 _7113_ (.A(_2207_),
    .B(_2211_),
    .Y(_2212_));
 sky130_fd_sc_hd__and3_1 _7114_ (.A(_1711_),
    .B(_4089_),
    .C(_1950_),
    .X(_2213_));
 sky130_fd_sc_hd__and2_1 _7115_ (.A(_2207_),
    .B(_2211_),
    .X(_2214_));
 sky130_fd_sc_hd__xnor2_1 _7116_ (.A(_2206_),
    .B(_2214_),
    .Y(_2215_));
 sky130_fd_sc_hd__nand2_1 _7117_ (.A(_2213_),
    .B(_2215_),
    .Y(_2216_));
 sky130_fd_sc_hd__o21ai_1 _7118_ (.A1(_2206_),
    .A2(_2212_),
    .B1(_2216_),
    .Y(_2217_));
 sky130_fd_sc_hd__and3_1 _7119_ (.A(_2202_),
    .B(_2204_),
    .C(_2217_),
    .X(_2218_));
 sky130_fd_sc_hd__a21oi_1 _7120_ (.A1(_2202_),
    .A2(_2204_),
    .B1(_2217_),
    .Y(_2219_));
 sky130_fd_sc_hd__nor2_1 _7121_ (.A(_2218_),
    .B(_2219_),
    .Y(_2220_));
 sky130_fd_sc_hd__or2_1 _7122_ (.A(_2213_),
    .B(_2215_),
    .X(_2222_));
 sky130_fd_sc_hd__nand2_1 _7123_ (.A(_2216_),
    .B(_2222_),
    .Y(_2223_));
 sky130_fd_sc_hd__nor2_1 _7124_ (.A(_2207_),
    .B(_2211_),
    .Y(_2224_));
 sky130_fd_sc_hd__nor2_1 _7125_ (.A(_2214_),
    .B(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__a21oi_1 _7126_ (.A1(_1782_),
    .A2(_2079_),
    .B1(_2225_),
    .Y(_2226_));
 sky130_fd_sc_hd__nor2_1 _7127_ (.A(_2160_),
    .B(_2209_),
    .Y(_2227_));
 sky130_fd_sc_hd__or2_1 _7128_ (.A(_2211_),
    .B(_2227_),
    .X(_2228_));
 sky130_fd_sc_hd__nand2_1 _7129_ (.A(_1531_),
    .B(_2079_),
    .Y(_2229_));
 sky130_fd_sc_hd__xor2_1 _7130_ (.A(_2228_),
    .B(_2229_),
    .X(_2230_));
 sky130_fd_sc_hd__o21ai_1 _7131_ (.A1(_1664_),
    .A2(_1676_),
    .B1(_2125_),
    .Y(_2231_));
 sky130_fd_sc_hd__and4_1 _7132_ (.A(_3804_),
    .B(_2079_),
    .C(_2185_),
    .D(_2231_),
    .X(_2233_));
 sky130_fd_sc_hd__and2_1 _7133_ (.A(_2230_),
    .B(_2233_),
    .X(_2234_));
 sky130_fd_sc_hd__o21ba_1 _7134_ (.A1(_2228_),
    .A2(_2229_),
    .B1_N(_2234_),
    .X(_2235_));
 sky130_fd_sc_hd__and3_1 _7135_ (.A(_1782_),
    .B(_2079_),
    .C(_2225_),
    .X(_2236_));
 sky130_fd_sc_hd__o21ba_1 _7136_ (.A1(_2226_),
    .A2(_2235_),
    .B1_N(_2236_),
    .X(_2237_));
 sky130_fd_sc_hd__nor2_1 _7137_ (.A(_2223_),
    .B(_2237_),
    .Y(_2238_));
 sky130_fd_sc_hd__a21o_1 _7138_ (.A1(_2220_),
    .A2(_2238_),
    .B1(_2218_),
    .X(_2239_));
 sky130_fd_sc_hd__a21o_1 _7139_ (.A1(_2197_),
    .A2(_2202_),
    .B1(_2182_),
    .X(_2240_));
 sky130_fd_sc_hd__a21bo_1 _7140_ (.A1(_2203_),
    .A2(_2239_),
    .B1_N(_2240_),
    .X(_2241_));
 sky130_fd_sc_hd__nor2_1 _7141_ (.A(_2152_),
    .B(_2180_),
    .Y(_2242_));
 sky130_fd_sc_hd__a21o_1 _7142_ (.A1(_2181_),
    .A2(_2241_),
    .B1(_2242_),
    .X(_2244_));
 sky130_fd_sc_hd__or2_1 _7143_ (.A(_2121_),
    .B(_2149_),
    .X(_2245_));
 sky130_fd_sc_hd__a21oi_1 _7144_ (.A1(_2118_),
    .A2(_2245_),
    .B1(_2119_),
    .Y(_2246_));
 sky130_fd_sc_hd__a41o_2 _7145_ (.A1(_2118_),
    .A2(_2120_),
    .A3(_2151_),
    .A4(_2244_),
    .B1(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__and2b_1 _7146_ (.A_N(_2044_),
    .B(_2043_),
    .X(_2248_));
 sky130_fd_sc_hd__and2_1 _7147_ (.A(_2009_),
    .B(_2046_),
    .X(_2249_));
 sky130_fd_sc_hd__xor2_1 _7148_ (.A(_1951_),
    .B(_1997_),
    .X(_2250_));
 sky130_fd_sc_hd__o21a_1 _7149_ (.A1(_2248_),
    .A2(_2249_),
    .B1(_2250_),
    .X(_2251_));
 sky130_fd_sc_hd__or3_1 _7150_ (.A(_2248_),
    .B(_2249_),
    .C(_2250_),
    .X(_2252_));
 sky130_fd_sc_hd__and2b_2 _7151_ (.A_N(_2251_),
    .B(_2252_),
    .X(_2253_));
 sky130_fd_sc_hd__o21a_1 _7152_ (.A1(_2251_),
    .A2(_2083_),
    .B1(_2252_),
    .X(_2255_));
 sky130_fd_sc_hd__a31oi_4 _7153_ (.A1(_2085_),
    .A2(_2247_),
    .A3(_2253_),
    .B1(_2255_),
    .Y(_2256_));
 sky130_fd_sc_hd__and2b_1 _7154_ (.A_N(_1999_),
    .B(_1949_),
    .X(_2257_));
 sky130_fd_sc_hd__or2_2 _7155_ (.A(_2000_),
    .B(_2257_),
    .X(_2258_));
 sky130_fd_sc_hd__xnor2_4 _7156_ (.A(_2003_),
    .B(_1948_),
    .Y(_2259_));
 sky130_fd_sc_hd__nor2_1 _7157_ (.A(_2258_),
    .B(_2259_),
    .Y(_2260_));
 sky130_fd_sc_hd__or4bb_1 _7158_ (.A(_1773_),
    .B(_2256_),
    .C_N(_2260_),
    .D_N(_1900_),
    .X(_2261_));
 sky130_fd_sc_hd__inv_2 _7159_ (.A(_1765_),
    .Y(_2262_));
 sky130_fd_sc_hd__and2b_1 _7160_ (.A_N(_1761_),
    .B(_1767_),
    .X(_2263_));
 sky130_fd_sc_hd__o21ai_1 _7161_ (.A1(_2262_),
    .A2(_2263_),
    .B1(_1769_),
    .Y(_2264_));
 sky130_fd_sc_hd__nand2_1 _7162_ (.A(_1584_),
    .B(_1618_),
    .Y(_2266_));
 sky130_fd_sc_hd__a21o_1 _7163_ (.A1(_1620_),
    .A2(_2266_),
    .B1(_1651_),
    .X(_2267_));
 sky130_fd_sc_hd__o21a_1 _7164_ (.A1(_1653_),
    .A2(_2264_),
    .B1(_2267_),
    .X(_2268_));
 sky130_fd_sc_hd__nor2_1 _7165_ (.A(_1648_),
    .B(_1650_),
    .Y(_2269_));
 sky130_fd_sc_hd__o21a_1 _7166_ (.A1(_1595_),
    .A2(_1597_),
    .B1(_1602_),
    .X(_2270_));
 sky130_fd_sc_hd__a22o_1 _7167_ (.A1(_2270_),
    .A2(_1628_),
    .B1(_1623_),
    .B2(_1629_),
    .X(_2271_));
 sky130_fd_sc_hd__and3_1 _7168_ (.A(_1588_),
    .B(_4251_),
    .C(_1498_),
    .X(_2272_));
 sky130_fd_sc_hd__or2_1 _7169_ (.A(_0080_),
    .B(_1446_),
    .X(_2273_));
 sky130_fd_sc_hd__nor2_1 _7170_ (.A(_4250_),
    .B(_0303_),
    .Y(_2274_));
 sky130_fd_sc_hd__and3b_1 _7171_ (.A_N(_2273_),
    .B(_1624_),
    .C(_2274_),
    .X(_2275_));
 sky130_fd_sc_hd__and3_1 _7172_ (.A(_0080_),
    .B(_1588_),
    .C(_2274_),
    .X(_2277_));
 sky130_fd_sc_hd__a211o_1 _7173_ (.A1(_4251_),
    .A2(_2273_),
    .B1(_2275_),
    .C1(_2277_),
    .X(_2278_));
 sky130_fd_sc_hd__nor2_1 _7174_ (.A(_1637_),
    .B(_2278_),
    .Y(_2279_));
 sky130_fd_sc_hd__and2_1 _7175_ (.A(_1637_),
    .B(_2278_),
    .X(_2280_));
 sky130_fd_sc_hd__nor2_1 _7176_ (.A(_2279_),
    .B(_2280_),
    .Y(_2281_));
 sky130_fd_sc_hd__and2_1 _7177_ (.A(_2272_),
    .B(_2281_),
    .X(_2282_));
 sky130_fd_sc_hd__nor2_1 _7178_ (.A(_2272_),
    .B(_2281_),
    .Y(_2283_));
 sky130_fd_sc_hd__or2_1 _7179_ (.A(_2282_),
    .B(_2283_),
    .X(_2284_));
 sky130_fd_sc_hd__and3_1 _7180_ (.A(_1593_),
    .B(_1596_),
    .C(_0121_),
    .X(_2285_));
 sky130_fd_sc_hd__xnor2_1 _7181_ (.A(_2284_),
    .B(_2285_),
    .Y(_2286_));
 sky130_fd_sc_hd__xnor2_1 _7182_ (.A(_1642_),
    .B(_2286_),
    .Y(_2288_));
 sky130_fd_sc_hd__xnor2_1 _7183_ (.A(_2271_),
    .B(_2288_),
    .Y(_2289_));
 sky130_fd_sc_hd__nor2_1 _7184_ (.A(_1644_),
    .B(_1646_),
    .Y(_2290_));
 sky130_fd_sc_hd__a21oi_1 _7185_ (.A1(_1622_),
    .A2(_1647_),
    .B1(_2290_),
    .Y(_2291_));
 sky130_fd_sc_hd__or2_1 _7186_ (.A(_2289_),
    .B(_2291_),
    .X(_2292_));
 sky130_fd_sc_hd__nand2_1 _7187_ (.A(_2289_),
    .B(_2291_),
    .Y(_2293_));
 sky130_fd_sc_hd__and2_1 _7188_ (.A(_2292_),
    .B(_2293_),
    .X(_2294_));
 sky130_fd_sc_hd__nand2_1 _7189_ (.A(_2269_),
    .B(_2294_),
    .Y(_2295_));
 sky130_fd_sc_hd__or2_1 _7190_ (.A(_2269_),
    .B(_2294_),
    .X(_2296_));
 sky130_fd_sc_hd__nand2_1 _7191_ (.A(_2295_),
    .B(_2296_),
    .Y(_2297_));
 sky130_fd_sc_hd__or3b_1 _7192_ (.A(_2282_),
    .B(_2283_),
    .C_N(_2285_),
    .X(_2299_));
 sky130_fd_sc_hd__o21ai_1 _7193_ (.A1(_0082_),
    .A2(_1446_),
    .B1(_0083_),
    .Y(_2300_));
 sky130_fd_sc_hd__o21ai_1 _7194_ (.A1(_2274_),
    .A2(_2273_),
    .B1(_2300_),
    .Y(_2301_));
 sky130_fd_sc_hd__o21bai_2 _7195_ (.A1(_1634_),
    .A2(_2301_),
    .B1_N(_2277_),
    .Y(_2302_));
 sky130_fd_sc_hd__and2_1 _7196_ (.A(_1634_),
    .B(_2301_),
    .X(_2303_));
 sky130_fd_sc_hd__nor2_1 _7197_ (.A(_2302_),
    .B(_2303_),
    .Y(_2304_));
 sky130_fd_sc_hd__xnor2_1 _7198_ (.A(_2299_),
    .B(_2304_),
    .Y(_2305_));
 sky130_fd_sc_hd__o21ai_1 _7199_ (.A1(_2279_),
    .A2(_2282_),
    .B1(_2305_),
    .Y(_2306_));
 sky130_fd_sc_hd__or3_1 _7200_ (.A(_2279_),
    .B(_2282_),
    .C(_2305_),
    .X(_2307_));
 sky130_fd_sc_hd__nand2_1 _7201_ (.A(_2306_),
    .B(_2307_),
    .Y(_2308_));
 sky130_fd_sc_hd__and3_1 _7202_ (.A(_1630_),
    .B(_1641_),
    .C(_2286_),
    .X(_2310_));
 sky130_fd_sc_hd__a21oi_1 _7203_ (.A1(_2271_),
    .A2(_2288_),
    .B1(_2310_),
    .Y(_2311_));
 sky130_fd_sc_hd__or2_1 _7204_ (.A(_2308_),
    .B(_2311_),
    .X(_2312_));
 sky130_fd_sc_hd__nand2_1 _7205_ (.A(_2308_),
    .B(_2311_),
    .Y(_2313_));
 sky130_fd_sc_hd__and2_1 _7206_ (.A(_2312_),
    .B(_2313_),
    .X(_2314_));
 sky130_fd_sc_hd__xor2_1 _7207_ (.A(_2292_),
    .B(_2314_),
    .X(_2315_));
 sky130_fd_sc_hd__a311o_1 _7208_ (.A1(_2008_),
    .A2(_2261_),
    .A3(_2268_),
    .B1(_2297_),
    .C1(_2315_),
    .X(_2316_));
 sky130_fd_sc_hd__a21bo_1 _7209_ (.A1(_2292_),
    .A2(_2295_),
    .B1_N(_2314_),
    .X(_2317_));
 sky130_fd_sc_hd__or3_1 _7210_ (.A(_2299_),
    .B(_2302_),
    .C(_2303_),
    .X(_2318_));
 sky130_fd_sc_hd__nor2_4 _7211_ (.A(_4250_),
    .B(_3989_),
    .Y(_2319_));
 sky130_fd_sc_hd__nand2_1 _7212_ (.A(_2273_),
    .B(_2319_),
    .Y(_2321_));
 sky130_fd_sc_hd__xor2_1 _7213_ (.A(_2302_),
    .B(_2321_),
    .X(_2322_));
 sky130_fd_sc_hd__a21o_1 _7214_ (.A1(_2318_),
    .A2(_2306_),
    .B1(_2322_),
    .X(_2323_));
 sky130_fd_sc_hd__nand3_1 _7215_ (.A(_2318_),
    .B(_2306_),
    .C(_2322_),
    .Y(_2324_));
 sky130_fd_sc_hd__nand2_1 _7216_ (.A(_2323_),
    .B(_2324_),
    .Y(_2325_));
 sky130_fd_sc_hd__xnor2_1 _7217_ (.A(_2312_),
    .B(_2325_),
    .Y(_2326_));
 sky130_fd_sc_hd__a21o_1 _7218_ (.A1(_2316_),
    .A2(_2317_),
    .B1(_2326_),
    .X(_2327_));
 sky130_fd_sc_hd__inv_2 _7219_ (.A(_2302_),
    .Y(_2328_));
 sky130_fd_sc_hd__o211a_1 _7220_ (.A1(_2328_),
    .A2(_0092_),
    .B1(_2323_),
    .C1(_2273_),
    .X(_2329_));
 sky130_fd_sc_hd__o21a_1 _7221_ (.A1(_2312_),
    .A2(_2325_),
    .B1(_2329_),
    .X(_2330_));
 sky130_fd_sc_hd__and4_1 _7222_ (.A(_3925_),
    .B(_3828_),
    .C(_3771_),
    .D(_3845_),
    .X(_2332_));
 sky130_fd_sc_hd__nand3b_2 _7223_ (.A_N(_0698_),
    .B(_0687_),
    .C(_2332_),
    .Y(_2333_));
 sky130_fd_sc_hd__and3_1 _7224_ (.A(_2327_),
    .B(_2330_),
    .C(_2333_),
    .X(_2334_));
 sky130_fd_sc_hd__clkbuf_4 _7225_ (.A(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__xnor2_1 _7226_ (.A(_0385_),
    .B(_2335_),
    .Y(_2336_));
 sky130_fd_sc_hd__nor2_1 _7227_ (.A(_0387_),
    .B(_2335_),
    .Y(_2337_));
 sky130_fd_sc_hd__a21oi_1 _7228_ (.A1(_0388_),
    .A2(_2336_),
    .B1(_2337_),
    .Y(_2338_));
 sky130_fd_sc_hd__nand2_1 _7229_ (.A(_3722_),
    .B(_0373_),
    .Y(_2339_));
 sky130_fd_sc_hd__o21a_1 _7230_ (.A1(_3722_),
    .A2(_3788_),
    .B1(_2339_),
    .X(_2340_));
 sky130_fd_sc_hd__xnor2_1 _7231_ (.A(_0369_),
    .B(_2338_),
    .Y(_2341_));
 sky130_fd_sc_hd__a2bb2o_2 _7232_ (.A1_N(_0370_),
    .A2_N(_2338_),
    .B1(_2340_),
    .B2(_2341_),
    .X(_2343_));
 sky130_fd_sc_hd__and2_1 _7233_ (.A(_0356_),
    .B(_0363_),
    .X(_2344_));
 sky130_fd_sc_hd__a21oi_1 _7234_ (.A1(_0603_),
    .A2(_2343_),
    .B1(_2344_),
    .Y(_2345_));
 sky130_fd_sc_hd__nor2_2 _7235_ (.A(_0346_),
    .B(_0350_),
    .Y(_2346_));
 sky130_fd_sc_hd__a211o_4 _7236_ (.A1(_0603_),
    .A2(_2343_),
    .B1(_2346_),
    .C1(_2344_),
    .X(_2347_));
 sky130_fd_sc_hd__o21a_1 _7237_ (.A1(_0351_),
    .A2(_2345_),
    .B1(_2347_),
    .X(_2348_));
 sky130_fd_sc_hd__or3_4 _7238_ (.A(_2980_),
    .B(_0082_),
    .C(_0400_),
    .X(_2349_));
 sky130_fd_sc_hd__inv_2 _7239_ (.A(_2349_),
    .Y(_2350_));
 sky130_fd_sc_hd__nand2_1 _7240_ (.A(_0349_),
    .B(_0433_),
    .Y(_2351_));
 sky130_fd_sc_hd__a21o_1 _7241_ (.A1(_0342_),
    .A2(_0349_),
    .B1(_0433_),
    .X(_2352_));
 sky130_fd_sc_hd__o21a_2 _7242_ (.A1(_0348_),
    .A2(_2351_),
    .B1(_2352_),
    .X(_2354_));
 sky130_fd_sc_hd__nand2_1 _7243_ (.A(_0430_),
    .B(_0425_),
    .Y(_2355_));
 sky130_fd_sc_hd__inv_2 _7244_ (.A(_2355_),
    .Y(_2356_));
 sky130_fd_sc_hd__nor2_1 _7245_ (.A(_0430_),
    .B(_0425_),
    .Y(_2357_));
 sky130_fd_sc_hd__nor2_2 _7246_ (.A(_2356_),
    .B(_2357_),
    .Y(_2358_));
 sky130_fd_sc_hd__and2_1 _7247_ (.A(_2354_),
    .B(_2358_),
    .X(_2359_));
 sky130_fd_sc_hd__and2b_1 _7248_ (.A_N(_0422_),
    .B(_0417_),
    .X(_2360_));
 sky130_fd_sc_hd__nor2_1 _7249_ (.A(_2360_),
    .B(_0415_),
    .Y(_2361_));
 sky130_fd_sc_hd__and2_1 _7250_ (.A(_2360_),
    .B(_0415_),
    .X(_2362_));
 sky130_fd_sc_hd__or2_1 _7251_ (.A(_2361_),
    .B(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__clkbuf_2 _7252_ (.A(_2363_),
    .X(_2365_));
 sky130_fd_sc_hd__and2b_1 _7253_ (.A_N(_0405_),
    .B(_0412_),
    .X(_2366_));
 sky130_fd_sc_hd__or2_1 _7254_ (.A(_2366_),
    .B(_0462_),
    .X(_2367_));
 sky130_fd_sc_hd__nand2_1 _7255_ (.A(_2366_),
    .B(_0462_),
    .Y(_2368_));
 sky130_fd_sc_hd__nand2_2 _7256_ (.A(_2367_),
    .B(_2368_),
    .Y(_2369_));
 sky130_fd_sc_hd__nor2_1 _7257_ (.A(_2365_),
    .B(_2369_),
    .Y(_2370_));
 sky130_fd_sc_hd__a21oi_1 _7258_ (.A1(_2352_),
    .A2(_2355_),
    .B1(_2357_),
    .Y(_2371_));
 sky130_fd_sc_hd__inv_2 _7259_ (.A(_2371_),
    .Y(_2372_));
 sky130_fd_sc_hd__o21ai_1 _7260_ (.A1(_2362_),
    .A2(_2372_),
    .B1(_2367_),
    .Y(_2373_));
 sky130_fd_sc_hd__o21a_1 _7261_ (.A1(_2361_),
    .A2(_2373_),
    .B1(_2368_),
    .X(_2374_));
 sky130_fd_sc_hd__a31oi_4 _7262_ (.A1(_2347_),
    .A2(_2359_),
    .A3(_2370_),
    .B1(_2374_),
    .Y(_2376_));
 sky130_fd_sc_hd__or3_1 _7263_ (.A(_2348_),
    .B(_2350_),
    .C(_2376_),
    .X(_2377_));
 sky130_fd_sc_hd__o21ai_2 _7264_ (.A1(_2350_),
    .A2(_2376_),
    .B1(_2348_),
    .Y(_2378_));
 sky130_fd_sc_hd__and2_1 _7265_ (.A(_2377_),
    .B(_2378_),
    .X(_2379_));
 sky130_fd_sc_hd__xnor2_1 _7266_ (.A(_2343_),
    .B(_0442_),
    .Y(_2380_));
 sky130_fd_sc_hd__xor2_2 _7267_ (.A(_0388_),
    .B(_2336_),
    .X(_2381_));
 sky130_fd_sc_hd__xnor2_2 _7268_ (.A(_0374_),
    .B(_2341_),
    .Y(_2382_));
 sky130_fd_sc_hd__nor2_1 _7269_ (.A(_2381_),
    .B(_2382_),
    .Y(_2383_));
 sky130_fd_sc_hd__o2111a_1 _7270_ (.A1(_0351_),
    .A2(_2345_),
    .B1(_2380_),
    .C1(_2383_),
    .D1(_2347_),
    .X(_2384_));
 sky130_fd_sc_hd__nand2_1 _7271_ (.A(_2384_),
    .B(_2354_),
    .Y(_2385_));
 sky130_fd_sc_hd__a21boi_2 _7272_ (.A1(_2347_),
    .A2(_2354_),
    .B1_N(_2352_),
    .Y(_2387_));
 sky130_fd_sc_hd__xnor2_4 _7273_ (.A(_2358_),
    .B(_2387_),
    .Y(_2388_));
 sky130_fd_sc_hd__a21oi_2 _7274_ (.A1(_2347_),
    .A2(_2359_),
    .B1(_2371_),
    .Y(_2389_));
 sky130_fd_sc_hd__xor2_1 _7275_ (.A(_2365_),
    .B(_2389_),
    .X(_2390_));
 sky130_fd_sc_hd__a31o_1 _7276_ (.A1(_2347_),
    .A2(_2359_),
    .A3(_2370_),
    .B1(_2374_),
    .X(_2391_));
 sky130_fd_sc_hd__nand2_2 _7277_ (.A(_2349_),
    .B(_2391_),
    .Y(_2392_));
 sky130_fd_sc_hd__o31a_2 _7278_ (.A1(_2385_),
    .A2(_2388_),
    .A3(_2390_),
    .B1(_2392_),
    .X(_2393_));
 sky130_fd_sc_hd__o21ba_1 _7279_ (.A1(_2362_),
    .A2(_2389_),
    .B1_N(_2361_),
    .X(_2394_));
 sky130_fd_sc_hd__xnor2_4 _7280_ (.A(_2369_),
    .B(_2394_),
    .Y(_2395_));
 sky130_fd_sc_hd__xnor2_1 _7281_ (.A(_2393_),
    .B(_2395_),
    .Y(_2396_));
 sky130_fd_sc_hd__xnor2_2 _7282_ (.A(_2365_),
    .B(_2389_),
    .Y(_2398_));
 sky130_fd_sc_hd__o211ai_4 _7283_ (.A1(_2385_),
    .A2(_2388_),
    .B1(_2398_),
    .C1(_2392_),
    .Y(_2399_));
 sky130_fd_sc_hd__o2bb2a_1 _7284_ (.A1_N(_2384_),
    .A2_N(_2354_),
    .B1(_2376_),
    .B2(_2350_),
    .X(_2400_));
 sky130_fd_sc_hd__a211o_1 _7285_ (.A1(_2392_),
    .A2(_2388_),
    .B1(_2398_),
    .C1(_2400_),
    .X(_2401_));
 sky130_fd_sc_hd__a21o_1 _7286_ (.A1(_2377_),
    .A2(_2378_),
    .B1(_2384_),
    .X(_2402_));
 sky130_fd_sc_hd__a21oi_2 _7287_ (.A1(_2349_),
    .A2(_2391_),
    .B1(_2384_),
    .Y(_2403_));
 sky130_fd_sc_hd__xor2_2 _7288_ (.A(_2347_),
    .B(_2354_),
    .X(_2404_));
 sky130_fd_sc_hd__xnor2_2 _7289_ (.A(_2403_),
    .B(_2404_),
    .Y(_2405_));
 sky130_fd_sc_hd__xnor2_2 _7290_ (.A(_2400_),
    .B(_2388_),
    .Y(_2406_));
 sky130_fd_sc_hd__a2111oi_2 _7291_ (.A1(_2399_),
    .A2(_2401_),
    .B1(_2402_),
    .C1(_2405_),
    .D1(_2406_),
    .Y(_2407_));
 sky130_fd_sc_hd__or3_1 _7292_ (.A(_2379_),
    .B(_2396_),
    .C(_2407_),
    .X(_2409_));
 sky130_fd_sc_hd__buf_2 _7293_ (.A(_2409_),
    .X(_2410_));
 sky130_fd_sc_hd__and3b_1 _7294_ (.A_N(_0698_),
    .B(_0687_),
    .C(_2332_),
    .X(_2411_));
 sky130_fd_sc_hd__buf_4 _7295_ (.A(_2411_),
    .X(_2412_));
 sky130_fd_sc_hd__o21bai_2 _7296_ (.A1(_2256_),
    .A2(_2258_),
    .B1_N(_2000_),
    .Y(_2413_));
 sky130_fd_sc_hd__xor2_4 _7297_ (.A(_2259_),
    .B(_2413_),
    .X(_2414_));
 sky130_fd_sc_hd__and2_1 _7298_ (.A(_2327_),
    .B(_2330_),
    .X(_2415_));
 sky130_fd_sc_hd__clkbuf_4 _7299_ (.A(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__a31o_1 _7300_ (.A1(_2085_),
    .A2(_2247_),
    .A3(_2253_),
    .B1(_2255_),
    .X(_2417_));
 sky130_fd_sc_hd__a21oi_1 _7301_ (.A1(_2417_),
    .A2(_2260_),
    .B1(_2004_),
    .Y(_2418_));
 sky130_fd_sc_hd__or2_1 _7302_ (.A(_1896_),
    .B(_2418_),
    .X(_2420_));
 sky130_fd_sc_hd__nand2_1 _7303_ (.A(_1896_),
    .B(_2418_),
    .Y(_2421_));
 sky130_fd_sc_hd__a21oi_1 _7304_ (.A1(_2420_),
    .A2(_2421_),
    .B1(_2412_),
    .Y(_2422_));
 sky130_fd_sc_hd__and2b_1 _7305_ (.A_N(_2416_),
    .B(_2422_),
    .X(_2423_));
 sky130_fd_sc_hd__a221oi_4 _7306_ (.A1(_1676_),
    .A2(_2412_),
    .B1(_2335_),
    .B2(_2414_),
    .C1(_2423_),
    .Y(_2424_));
 sky130_fd_sc_hd__nand2_2 _7307_ (.A(_2377_),
    .B(_2378_),
    .Y(_2425_));
 sky130_fd_sc_hd__xor2_4 _7308_ (.A(_2393_),
    .B(_2395_),
    .X(_2426_));
 sky130_fd_sc_hd__a2111o_4 _7309_ (.A1(_2399_),
    .A2(_2401_),
    .B1(_2402_),
    .C1(_2405_),
    .D1(_2406_),
    .X(_2427_));
 sky130_fd_sc_hd__o21ai_1 _7310_ (.A1(_1896_),
    .A2(_2418_),
    .B1(_2005_),
    .Y(_2428_));
 sky130_fd_sc_hd__nand2_1 _7311_ (.A(_1899_),
    .B(_2428_),
    .Y(_2429_));
 sky130_fd_sc_hd__buf_2 _7312_ (.A(_2333_),
    .X(_2431_));
 sky130_fd_sc_hd__o211a_1 _7313_ (.A1(_1899_),
    .A2(_2428_),
    .B1(_2429_),
    .C1(_2431_),
    .X(_2432_));
 sky130_fd_sc_hd__mux2_1 _7314_ (.A0(_2432_),
    .A1(_2422_),
    .S(_2416_),
    .X(_2433_));
 sky130_fd_sc_hd__a21oi_1 _7315_ (.A1(_1456_),
    .A2(_2412_),
    .B1(_2433_),
    .Y(_2434_));
 sky130_fd_sc_hd__a31o_1 _7316_ (.A1(_2425_),
    .A2(_2426_),
    .A3(_2427_),
    .B1(_2434_),
    .X(_2435_));
 sky130_fd_sc_hd__o21a_1 _7317_ (.A1(_2410_),
    .A2(_2424_),
    .B1(_2435_),
    .X(_2436_));
 sky130_fd_sc_hd__or2_2 _7318_ (.A(_2416_),
    .B(_2412_),
    .X(_2437_));
 sky130_fd_sc_hd__xnor2_2 _7319_ (.A(_2256_),
    .B(_2258_),
    .Y(_2438_));
 sky130_fd_sc_hd__a21oi_1 _7320_ (.A1(_2085_),
    .A2(_2247_),
    .B1(_2083_),
    .Y(_2439_));
 sky130_fd_sc_hd__xor2_2 _7321_ (.A(_2253_),
    .B(_2439_),
    .X(_2440_));
 sky130_fd_sc_hd__nand2_1 _7322_ (.A(_2416_),
    .B(_2431_),
    .Y(_2442_));
 sky130_fd_sc_hd__o22ai_2 _7323_ (.A1(_2437_),
    .A2(_2438_),
    .B1(_2440_),
    .B2(_2442_),
    .Y(_2443_));
 sky130_fd_sc_hd__clkinv_2 _7324_ (.A(_2437_),
    .Y(_2444_));
 sky130_fd_sc_hd__nor2_1 _7325_ (.A(_3804_),
    .B(_2431_),
    .Y(_2445_));
 sky130_fd_sc_hd__a221oi_2 _7326_ (.A1(_2414_),
    .A2(_2444_),
    .B1(_2438_),
    .B2(_2335_),
    .C1(_2445_),
    .Y(_2446_));
 sky130_fd_sc_hd__mux2_1 _7327_ (.A0(_2443_),
    .A1(_2446_),
    .S(_2410_),
    .X(_2447_));
 sky130_fd_sc_hd__xor2_1 _7328_ (.A(_2403_),
    .B(_2404_),
    .X(_2448_));
 sky130_fd_sc_hd__xnor2_1 _7329_ (.A(_2402_),
    .B(_2448_),
    .Y(_2449_));
 sky130_fd_sc_hd__and3b_1 _7330_ (.A_N(_2449_),
    .B(_2426_),
    .C(_2427_),
    .X(_2450_));
 sky130_fd_sc_hd__buf_2 _7331_ (.A(_2450_),
    .X(_2451_));
 sky130_fd_sc_hd__mux2_1 _7332_ (.A0(_2436_),
    .A1(_2447_),
    .S(_2451_),
    .X(_2453_));
 sky130_fd_sc_hd__buf_2 _7333_ (.A(_2409_),
    .X(_2454_));
 sky130_fd_sc_hd__a31oi_1 _7334_ (.A1(_1900_),
    .A2(_2417_),
    .A3(_2260_),
    .B1(_2007_),
    .Y(_2455_));
 sky130_fd_sc_hd__nor2_1 _7335_ (.A(_1768_),
    .B(_2455_),
    .Y(_2456_));
 sky130_fd_sc_hd__and2_1 _7336_ (.A(_1768_),
    .B(_2455_),
    .X(_2457_));
 sky130_fd_sc_hd__nor2_1 _7337_ (.A(_2456_),
    .B(_2457_),
    .Y(_2458_));
 sky130_fd_sc_hd__nand2_1 _7338_ (.A(_2416_),
    .B(_2432_),
    .Y(_2459_));
 sky130_fd_sc_hd__o221a_1 _7339_ (.A1(_4089_),
    .A2(_2431_),
    .B1(_2437_),
    .B2(_2458_),
    .C1(_2459_),
    .X(_2460_));
 sky130_fd_sc_hd__nor2_1 _7340_ (.A(_2263_),
    .B(_2456_),
    .Y(_2461_));
 sky130_fd_sc_hd__xnor2_1 _7341_ (.A(_1771_),
    .B(_2461_),
    .Y(_2462_));
 sky130_fd_sc_hd__or2_1 _7342_ (.A(_2442_),
    .B(_2458_),
    .X(_2464_));
 sky130_fd_sc_hd__o221a_1 _7343_ (.A1(_0147_),
    .A2(_2431_),
    .B1(_2437_),
    .B2(_2462_),
    .C1(_2464_),
    .X(_2465_));
 sky130_fd_sc_hd__a31o_1 _7344_ (.A1(_2425_),
    .A2(_2426_),
    .A3(_2427_),
    .B1(_2465_),
    .X(_2466_));
 sky130_fd_sc_hd__o21ai_1 _7345_ (.A1(_2454_),
    .A2(_2460_),
    .B1(_2466_),
    .Y(_2467_));
 sky130_fd_sc_hd__a21boi_1 _7346_ (.A1(_1771_),
    .A2(_2456_),
    .B1_N(_2264_),
    .Y(_2468_));
 sky130_fd_sc_hd__o21a_1 _7347_ (.A1(_1619_),
    .A2(_2468_),
    .B1(_2266_),
    .X(_2469_));
 sky130_fd_sc_hd__xnor2_2 _7348_ (.A(_1652_),
    .B(_2469_),
    .Y(_2470_));
 sky130_fd_sc_hd__xnor2_1 _7349_ (.A(_1619_),
    .B(_2468_),
    .Y(_2471_));
 sky130_fd_sc_hd__and2_1 _7350_ (.A(_2335_),
    .B(_2471_),
    .X(_2472_));
 sky130_fd_sc_hd__a221oi_4 _7351_ (.A1(_1428_),
    .A2(_2412_),
    .B1(_2444_),
    .B2(_2470_),
    .C1(_2472_),
    .Y(_2473_));
 sky130_fd_sc_hd__a31o_1 _7352_ (.A1(_2425_),
    .A2(_2426_),
    .A3(_2427_),
    .B1(_2473_),
    .X(_2475_));
 sky130_fd_sc_hd__nand2_1 _7353_ (.A(_2444_),
    .B(_2471_),
    .Y(_2476_));
 sky130_fd_sc_hd__o221a_1 _7354_ (.A1(_3986_),
    .A2(_2431_),
    .B1(_2442_),
    .B2(_2462_),
    .C1(_2476_),
    .X(_2477_));
 sky130_fd_sc_hd__or4_1 _7355_ (.A(_2379_),
    .B(_2396_),
    .C(_2407_),
    .D(_2477_),
    .X(_2478_));
 sky130_fd_sc_hd__a21oi_1 _7356_ (.A1(_2475_),
    .A2(_2478_),
    .B1(_2451_),
    .Y(_2479_));
 sky130_fd_sc_hd__a21oi_1 _7357_ (.A1(_2451_),
    .A2(_2467_),
    .B1(_2479_),
    .Y(_2480_));
 sky130_fd_sc_hd__nand2_1 _7358_ (.A(_2426_),
    .B(_2427_),
    .Y(_2481_));
 sky130_fd_sc_hd__nor2_1 _7359_ (.A(_2402_),
    .B(_2405_),
    .Y(_2482_));
 sky130_fd_sc_hd__xnor2_1 _7360_ (.A(_2482_),
    .B(_2406_),
    .Y(_2483_));
 sky130_fd_sc_hd__or2_1 _7361_ (.A(_2481_),
    .B(_2483_),
    .X(_2484_));
 sky130_fd_sc_hd__clkbuf_4 _7362_ (.A(_2484_),
    .X(_2486_));
 sky130_fd_sc_hd__mux2_1 _7363_ (.A0(_2453_),
    .A1(_2480_),
    .S(_2486_),
    .X(_2487_));
 sky130_fd_sc_hd__xor2_2 _7364_ (.A(_2343_),
    .B(_0442_),
    .X(_2488_));
 sky130_fd_sc_hd__a31o_1 _7365_ (.A1(_2425_),
    .A2(_2426_),
    .A3(_2427_),
    .B1(_2488_),
    .X(_2489_));
 sky130_fd_sc_hd__o21a_1 _7366_ (.A1(_2382_),
    .A2(_2410_),
    .B1(_2489_),
    .X(_2490_));
 sky130_fd_sc_hd__nor2_1 _7367_ (.A(_2350_),
    .B(_2376_),
    .Y(_2491_));
 sky130_fd_sc_hd__a2bb2o_1 _7368_ (.A1_N(_2378_),
    .A2_N(_2481_),
    .B1(_2410_),
    .B2(_2491_),
    .X(_2492_));
 sky130_fd_sc_hd__or3_1 _7369_ (.A(_2396_),
    .B(_2407_),
    .C(_2449_),
    .X(_2493_));
 sky130_fd_sc_hd__buf_2 _7370_ (.A(_2493_),
    .X(_2494_));
 sky130_fd_sc_hd__mux2_1 _7371_ (.A0(_2490_),
    .A1(_2492_),
    .S(_2494_),
    .X(_2495_));
 sky130_fd_sc_hd__and3_1 _7372_ (.A(_2008_),
    .B(_2261_),
    .C(_2268_),
    .X(_2497_));
 sky130_fd_sc_hd__xor2_1 _7373_ (.A(_2297_),
    .B(_2497_),
    .X(_2498_));
 sky130_fd_sc_hd__or2_1 _7374_ (.A(_2412_),
    .B(_2498_),
    .X(_2499_));
 sky130_fd_sc_hd__nand2_1 _7375_ (.A(_2335_),
    .B(_2470_),
    .Y(_2500_));
 sky130_fd_sc_hd__o221a_1 _7376_ (.A1(_4153_),
    .A2(_2431_),
    .B1(_2499_),
    .B2(_2416_),
    .C1(_2500_),
    .X(_2501_));
 sky130_fd_sc_hd__o21a_1 _7377_ (.A1(_2297_),
    .A2(_2497_),
    .B1(_2295_),
    .X(_2502_));
 sky130_fd_sc_hd__xor2_1 _7378_ (.A(_2315_),
    .B(_2502_),
    .X(_2503_));
 sky130_fd_sc_hd__a21oi_1 _7379_ (.A1(_2316_),
    .A2(_2317_),
    .B1(_2326_),
    .Y(_2504_));
 sky130_fd_sc_hd__or3b_1 _7380_ (.A(_2499_),
    .B(_2504_),
    .C_N(_2330_),
    .X(_2505_));
 sky130_fd_sc_hd__o221a_1 _7381_ (.A1(_4217_),
    .A2(_2431_),
    .B1(_2437_),
    .B2(_2503_),
    .C1(_2505_),
    .X(_2506_));
 sky130_fd_sc_hd__mux2_1 _7382_ (.A0(_2501_),
    .A1(_2506_),
    .S(_2410_),
    .X(_2508_));
 sky130_fd_sc_hd__and3_1 _7383_ (.A(_2316_),
    .B(_2317_),
    .C(_2326_),
    .X(_2509_));
 sky130_fd_sc_hd__o21ai_1 _7384_ (.A1(_2504_),
    .A2(_2509_),
    .B1(_2444_),
    .Y(_2510_));
 sky130_fd_sc_hd__o221a_1 _7385_ (.A1(_0218_),
    .A2(_2431_),
    .B1(_2442_),
    .B2(_2503_),
    .C1(_2510_),
    .X(_2511_));
 sky130_fd_sc_hd__mux2_1 _7386_ (.A0(_2511_),
    .A1(_2381_),
    .S(_2409_),
    .X(_2512_));
 sky130_fd_sc_hd__mux2_1 _7387_ (.A0(_2508_),
    .A1(_2512_),
    .S(_2494_),
    .X(_2513_));
 sky130_fd_sc_hd__nor2_4 _7388_ (.A(_2481_),
    .B(_2483_),
    .Y(_2514_));
 sky130_fd_sc_hd__mux2_1 _7389_ (.A0(_2495_),
    .A1(_2513_),
    .S(_2514_),
    .X(_2515_));
 sky130_fd_sc_hd__nand2_1 _7390_ (.A(_2399_),
    .B(_2401_),
    .Y(_2516_));
 sky130_fd_sc_hd__or3_1 _7391_ (.A(_2402_),
    .B(_2405_),
    .C(_2406_),
    .X(_2517_));
 sky130_fd_sc_hd__or3b_1 _7392_ (.A(_2516_),
    .B(_2396_),
    .C_N(_2517_),
    .X(_2519_));
 sky130_fd_sc_hd__buf_2 _7393_ (.A(_2519_),
    .X(_2520_));
 sky130_fd_sc_hd__mux2_2 _7394_ (.A0(_2487_),
    .A1(_2515_),
    .S(_2520_),
    .X(_2521_));
 sky130_fd_sc_hd__buf_2 _7395_ (.A(_2494_),
    .X(_2522_));
 sky130_fd_sc_hd__mux2_1 _7396_ (.A0(_2446_),
    .A1(_2424_),
    .S(_2410_),
    .X(_2523_));
 sky130_fd_sc_hd__xor2_2 _7397_ (.A(_2085_),
    .B(_2247_),
    .X(_2524_));
 sky130_fd_sc_hd__a2bb2o_1 _7398_ (.A1_N(_2437_),
    .A2_N(_2440_),
    .B1(_2524_),
    .B2(_2335_),
    .X(_2525_));
 sky130_fd_sc_hd__a31o_1 _7399_ (.A1(_2425_),
    .A2(_2426_),
    .A3(_2427_),
    .B1(_2443_),
    .X(_2526_));
 sky130_fd_sc_hd__o211a_1 _7400_ (.A1(_2454_),
    .A2(_2525_),
    .B1(_2526_),
    .C1(_2451_),
    .X(_2527_));
 sky130_fd_sc_hd__a21o_1 _7401_ (.A1(_2522_),
    .A2(_2523_),
    .B1(_2527_),
    .X(_2528_));
 sky130_fd_sc_hd__nand2_1 _7402_ (.A(_2118_),
    .B(_2120_),
    .Y(_2530_));
 sky130_fd_sc_hd__nand2_1 _7403_ (.A(_2151_),
    .B(_2244_),
    .Y(_2531_));
 sky130_fd_sc_hd__and2_1 _7404_ (.A(_2245_),
    .B(_2531_),
    .X(_2532_));
 sky130_fd_sc_hd__a21oi_1 _7405_ (.A1(_2530_),
    .A2(_2532_),
    .B1(_2412_),
    .Y(_2533_));
 sky130_fd_sc_hd__o21a_1 _7406_ (.A1(_2530_),
    .A2(_2532_),
    .B1(_2533_),
    .X(_2534_));
 sky130_fd_sc_hd__a22o_1 _7407_ (.A1(_2444_),
    .A2(_2524_),
    .B1(_2534_),
    .B2(_2416_),
    .X(_2535_));
 sky130_fd_sc_hd__xnor2_2 _7408_ (.A(_2151_),
    .B(_2244_),
    .Y(_2536_));
 sky130_fd_sc_hd__inv_2 _7409_ (.A(_2534_),
    .Y(_2537_));
 sky130_fd_sc_hd__o22ai_1 _7410_ (.A1(_2442_),
    .A2(_2536_),
    .B1(_2537_),
    .B2(_2416_),
    .Y(_2538_));
 sky130_fd_sc_hd__mux2_1 _7411_ (.A0(_2538_),
    .A1(_2525_),
    .S(_2454_),
    .X(_2539_));
 sky130_fd_sc_hd__or2_1 _7412_ (.A(_2535_),
    .B(_2539_),
    .X(_2541_));
 sky130_fd_sc_hd__and2b_1 _7413_ (.A_N(_2239_),
    .B(_2240_),
    .X(_2542_));
 sky130_fd_sc_hd__nand2_1 _7414_ (.A(_0548_),
    .B(_2158_),
    .Y(_2543_));
 sky130_fd_sc_hd__a32o_1 _7415_ (.A1(_2185_),
    .A2(_2543_),
    .A3(_2231_),
    .B1(_2079_),
    .B2(_3804_),
    .X(_2544_));
 sky130_fd_sc_hd__o21ba_1 _7416_ (.A1(_2230_),
    .A2(_2544_),
    .B1_N(_2234_),
    .X(_2545_));
 sky130_fd_sc_hd__nor2_1 _7417_ (.A(_1664_),
    .B(_0548_),
    .Y(_2546_));
 sky130_fd_sc_hd__o22a_1 _7418_ (.A1(_1531_),
    .A2(_3804_),
    .B1(_1813_),
    .B2(_2546_),
    .X(_2547_));
 sky130_fd_sc_hd__and2_1 _7419_ (.A(_2223_),
    .B(_2226_),
    .X(_2548_));
 sky130_fd_sc_hd__mux2_1 _7420_ (.A0(_2548_),
    .A1(_2238_),
    .S(_2220_),
    .X(_2549_));
 sky130_fd_sc_hd__or3b_1 _7421_ (.A(_2545_),
    .B(_2547_),
    .C_N(_2549_),
    .X(_2550_));
 sky130_fd_sc_hd__or2b_1 _7422_ (.A(_2242_),
    .B_N(_2181_),
    .X(_2552_));
 sky130_fd_sc_hd__xnor2_1 _7423_ (.A(_2552_),
    .B(_2542_),
    .Y(_2553_));
 sky130_fd_sc_hd__nand2_1 _7424_ (.A(_2536_),
    .B(_2553_),
    .Y(_2554_));
 sky130_fd_sc_hd__xnor2_1 _7425_ (.A(_2552_),
    .B(_2241_),
    .Y(_2555_));
 sky130_fd_sc_hd__mux2_1 _7426_ (.A0(_2554_),
    .A1(_2555_),
    .S(_2416_),
    .X(_2556_));
 sky130_fd_sc_hd__a211o_1 _7427_ (.A1(_2203_),
    .A2(_2542_),
    .B1(_2550_),
    .C1(_2556_),
    .X(_2557_));
 sky130_fd_sc_hd__a22o_1 _7428_ (.A1(_2454_),
    .A2(_2538_),
    .B1(_2557_),
    .B2(_2431_),
    .X(_2558_));
 sky130_fd_sc_hd__or3_1 _7429_ (.A(_2522_),
    .B(_2447_),
    .C(_2558_),
    .X(_2559_));
 sky130_fd_sc_hd__o41a_1 _7430_ (.A1(_2451_),
    .A2(_2436_),
    .A3(_2514_),
    .A4(_2541_),
    .B1(_2559_),
    .X(_2560_));
 sky130_fd_sc_hd__a31o_1 _7431_ (.A1(_2425_),
    .A2(_2426_),
    .A3(_2427_),
    .B1(_2460_),
    .X(_2561_));
 sky130_fd_sc_hd__or4_1 _7432_ (.A(_2379_),
    .B(_2396_),
    .C(_2407_),
    .D(_2434_),
    .X(_2563_));
 sky130_fd_sc_hd__and3_1 _7433_ (.A(_2494_),
    .B(_2561_),
    .C(_2563_),
    .X(_2564_));
 sky130_fd_sc_hd__a21oi_1 _7434_ (.A1(_2451_),
    .A2(_2523_),
    .B1(_2564_),
    .Y(_2565_));
 sky130_fd_sc_hd__o21ai_1 _7435_ (.A1(_2454_),
    .A2(_2424_),
    .B1(_2435_),
    .Y(_2566_));
 sky130_fd_sc_hd__mux2_1 _7436_ (.A0(_2566_),
    .A1(_2467_),
    .S(_2494_),
    .X(_2567_));
 sky130_fd_sc_hd__nand2_1 _7437_ (.A(_2565_),
    .B(_2567_),
    .Y(_2568_));
 sky130_fd_sc_hd__buf_2 _7438_ (.A(_2486_),
    .X(_2569_));
 sky130_fd_sc_hd__a211o_1 _7439_ (.A1(_2449_),
    .A2(_2541_),
    .B1(_2558_),
    .C1(_2569_),
    .X(_2570_));
 sky130_fd_sc_hd__o31a_1 _7440_ (.A1(_2528_),
    .A2(_2560_),
    .A3(_2568_),
    .B1(_2570_),
    .X(_2571_));
 sky130_fd_sc_hd__o21a_1 _7441_ (.A1(_2454_),
    .A2(_2525_),
    .B1(_2526_),
    .X(_2572_));
 sky130_fd_sc_hd__a211o_1 _7442_ (.A1(_2569_),
    .A2(_2558_),
    .B1(_2572_),
    .C1(_2447_),
    .X(_2574_));
 sky130_fd_sc_hd__mux2_1 _7443_ (.A0(_2541_),
    .A1(_2574_),
    .S(_2522_),
    .X(_2575_));
 sky130_fd_sc_hd__mux2_1 _7444_ (.A0(_2480_),
    .A1(_2513_),
    .S(_2569_),
    .X(_2576_));
 sky130_fd_sc_hd__mux2_1 _7445_ (.A0(_2473_),
    .A1(_2501_),
    .S(_2410_),
    .X(_2577_));
 sky130_fd_sc_hd__mux2_1 _7446_ (.A0(_2506_),
    .A1(_2511_),
    .S(_2410_),
    .X(_2578_));
 sky130_fd_sc_hd__mux2_1 _7447_ (.A0(_2577_),
    .A1(_2578_),
    .S(_2494_),
    .X(_2579_));
 sky130_fd_sc_hd__a31o_1 _7448_ (.A1(_2425_),
    .A2(_2426_),
    .A3(_2427_),
    .B1(_2477_),
    .X(_2580_));
 sky130_fd_sc_hd__o21a_1 _7449_ (.A1(_2454_),
    .A2(_2465_),
    .B1(_2580_),
    .X(_2581_));
 sky130_fd_sc_hd__and3_1 _7450_ (.A(_2450_),
    .B(_2561_),
    .C(_2563_),
    .X(_2582_));
 sky130_fd_sc_hd__a211o_1 _7451_ (.A1(_2522_),
    .A2(_2581_),
    .B1(_2582_),
    .C1(_2569_),
    .X(_2583_));
 sky130_fd_sc_hd__o21ai_1 _7452_ (.A1(_2514_),
    .A2(_2579_),
    .B1(_2583_),
    .Y(_2585_));
 sky130_fd_sc_hd__o211a_1 _7453_ (.A1(_2454_),
    .A2(_2465_),
    .B1(_2580_),
    .C1(_2451_),
    .X(_2586_));
 sky130_fd_sc_hd__a21oi_1 _7454_ (.A1(_2522_),
    .A2(_2577_),
    .B1(_2586_),
    .Y(_2587_));
 sky130_fd_sc_hd__mux2_1 _7455_ (.A0(_2565_),
    .A1(_2587_),
    .S(_2486_),
    .X(_2588_));
 sky130_fd_sc_hd__a31o_1 _7456_ (.A1(_2425_),
    .A2(_2426_),
    .A3(_2427_),
    .B1(_2382_),
    .X(_2589_));
 sky130_fd_sc_hd__o211a_1 _7457_ (.A1(_2381_),
    .A2(_2454_),
    .B1(_2589_),
    .C1(_2493_),
    .X(_2590_));
 sky130_fd_sc_hd__a21oi_1 _7458_ (.A1(_2451_),
    .A2(_2578_),
    .B1(_2590_),
    .Y(_2591_));
 sky130_fd_sc_hd__mux2_1 _7459_ (.A0(_2587_),
    .A1(_2591_),
    .S(_2569_),
    .X(_2592_));
 sky130_fd_sc_hd__and3_1 _7460_ (.A(_2450_),
    .B(_2475_),
    .C(_2478_),
    .X(_2593_));
 sky130_fd_sc_hd__a21oi_1 _7461_ (.A1(_2522_),
    .A2(_2508_),
    .B1(_2593_),
    .Y(_2594_));
 sky130_fd_sc_hd__o211a_1 _7462_ (.A1(_2382_),
    .A2(_2454_),
    .B1(_2489_),
    .C1(_2494_),
    .X(_2596_));
 sky130_fd_sc_hd__a21oi_1 _7463_ (.A1(_2451_),
    .A2(_2512_),
    .B1(_2596_),
    .Y(_2597_));
 sky130_fd_sc_hd__mux2_1 _7464_ (.A0(_2594_),
    .A1(_2597_),
    .S(_2486_),
    .X(_2598_));
 sky130_fd_sc_hd__nand4_1 _7465_ (.A(_2585_),
    .B(_2588_),
    .C(_2592_),
    .D(_2598_),
    .Y(_2599_));
 sky130_fd_sc_hd__a211o_1 _7466_ (.A1(_2522_),
    .A2(_2581_),
    .B1(_2582_),
    .C1(_2514_),
    .X(_2600_));
 sky130_fd_sc_hd__a211o_1 _7467_ (.A1(_2522_),
    .A2(_2523_),
    .B1(_2527_),
    .C1(_2486_),
    .X(_2601_));
 sky130_fd_sc_hd__mux2_1 _7468_ (.A0(_2594_),
    .A1(_2567_),
    .S(_2514_),
    .X(_2602_));
 sky130_fd_sc_hd__a21bo_1 _7469_ (.A1(_2600_),
    .A2(_2601_),
    .B1_N(_2602_),
    .X(_2603_));
 sky130_fd_sc_hd__buf_2 _7470_ (.A(_2520_),
    .X(_2604_));
 sky130_fd_sc_hd__o41a_1 _7471_ (.A1(_2487_),
    .A2(_2576_),
    .A3(_2599_),
    .A4(_2603_),
    .B1(_2604_),
    .X(_2605_));
 sky130_fd_sc_hd__or4_1 _7472_ (.A(_2521_),
    .B(_2571_),
    .C(_2575_),
    .D(_2605_),
    .X(_2607_));
 sky130_fd_sc_hd__and3_1 _7473_ (.A(_2379_),
    .B(_2448_),
    .C(_2516_),
    .X(_2608_));
 sky130_fd_sc_hd__a21oi_1 _7474_ (.A1(_2520_),
    .A2(_2569_),
    .B1(_2608_),
    .Y(_2609_));
 sky130_fd_sc_hd__a21o_1 _7475_ (.A1(_2607_),
    .A2(_2609_),
    .B1(_1308_),
    .X(_2610_));
 sky130_fd_sc_hd__inv_2 _7476_ (.A(_2520_),
    .Y(_2611_));
 sky130_fd_sc_hd__o21a_1 _7477_ (.A1(_2381_),
    .A2(_2410_),
    .B1(_2589_),
    .X(_2612_));
 sky130_fd_sc_hd__mux2_1 _7478_ (.A0(_2488_),
    .A1(_2392_),
    .S(_2410_),
    .X(_2613_));
 sky130_fd_sc_hd__mux2_1 _7479_ (.A0(_2612_),
    .A1(_2613_),
    .S(_2494_),
    .X(_2614_));
 sky130_fd_sc_hd__mux2_1 _7480_ (.A0(_2579_),
    .A1(_2614_),
    .S(_2486_),
    .X(_2615_));
 sky130_fd_sc_hd__a21o_1 _7481_ (.A1(_2600_),
    .A2(_2601_),
    .B1(_2520_),
    .X(_2616_));
 sky130_fd_sc_hd__o21a_1 _7482_ (.A1(_2611_),
    .A2(_2615_),
    .B1(_2616_),
    .X(_2618_));
 sky130_fd_sc_hd__and3_1 _7483_ (.A(_2521_),
    .B(_2610_),
    .C(_2618_),
    .X(_2619_));
 sky130_fd_sc_hd__or3b_1 _7484_ (.A(\cmd[6] ),
    .B(_0092_),
    .C_N(\cmd[7] ),
    .X(_2620_));
 sky130_fd_sc_hd__buf_2 _7485_ (.A(_2620_),
    .X(_2621_));
 sky130_fd_sc_hd__a21oi_1 _7486_ (.A1(_2610_),
    .A2(_2618_),
    .B1(_2521_),
    .Y(_2622_));
 sky130_fd_sc_hd__nand2_1 _7487_ (.A(_3328_),
    .B(_0347_),
    .Y(_2623_));
 sky130_fd_sc_hd__inv_2 _7488_ (.A(_3035_),
    .Y(_2624_));
 sky130_fd_sc_hd__or2_1 _7489_ (.A(_2624_),
    .B(_1539_),
    .X(_2625_));
 sky130_fd_sc_hd__xnor2_1 _7490_ (.A(\posit_add.in1[7] ),
    .B(_2683_),
    .Y(_2626_));
 sky130_fd_sc_hd__nor2_1 _7491_ (.A(_2826_),
    .B(_0402_),
    .Y(_2627_));
 sky130_fd_sc_hd__inv_2 _7492_ (.A(_1913_),
    .Y(_2629_));
 sky130_fd_sc_hd__a211o_1 _7493_ (.A1(\posit_add.in1[1] ),
    .A2(_2034_),
    .B1(_3765_),
    .C1(_2969_),
    .X(_2630_));
 sky130_fd_sc_hd__o221a_1 _7494_ (.A1(_3189_),
    .A2(_1803_),
    .B1(_2034_),
    .B2(_3232_),
    .C1(_2630_),
    .X(_2631_));
 sky130_fd_sc_hd__a22o_1 _7495_ (.A1(_2936_),
    .A2(_1836_),
    .B1(_1803_),
    .B2(_3189_),
    .X(_2632_));
 sky130_fd_sc_hd__or2_1 _7496_ (.A(_2936_),
    .B(_1836_),
    .X(_2633_));
 sky130_fd_sc_hd__o221a_1 _7497_ (.A1(_2903_),
    .A2(_1858_),
    .B1(_2631_),
    .B2(_2632_),
    .C1(_2633_),
    .X(_2634_));
 sky130_fd_sc_hd__a22o_1 _7498_ (.A1(_2859_),
    .A2(_2629_),
    .B1(_1858_),
    .B2(_2903_),
    .X(_2635_));
 sky130_fd_sc_hd__o22a_1 _7499_ (.A1(_2859_),
    .A2(_2629_),
    .B1(_2634_),
    .B2(_2635_),
    .X(_2636_));
 sky130_fd_sc_hd__a21oi_1 _7500_ (.A1(_2826_),
    .A2(_0402_),
    .B1(_2636_),
    .Y(_2637_));
 sky130_fd_sc_hd__o22a_1 _7501_ (.A1(_2626_),
    .A2(_1682_),
    .B1(_2627_),
    .B2(_2637_),
    .X(_2638_));
 sky130_fd_sc_hd__a221o_1 _7502_ (.A1(_2626_),
    .A2(_1682_),
    .B1(_3643_),
    .B2(_2639_),
    .C1(_2638_),
    .X(_2640_));
 sky130_fd_sc_hd__o2bb2a_1 _7503_ (.A1_N(_2760_),
    .A2_N(_3919_),
    .B1(_3643_),
    .B2(_2639_),
    .X(_2641_));
 sky130_fd_sc_hd__o22ai_1 _7504_ (.A1(_2727_),
    .A2(_1583_),
    .B1(_3919_),
    .B2(_2760_),
    .Y(_2642_));
 sky130_fd_sc_hd__a21oi_1 _7505_ (.A1(_2640_),
    .A2(_2641_),
    .B1(_2642_),
    .Y(_2643_));
 sky130_fd_sc_hd__a22o_1 _7506_ (.A1(_3101_),
    .A2(_1484_),
    .B1(_1583_),
    .B2(_2727_),
    .X(_2644_));
 sky130_fd_sc_hd__or2_1 _7507_ (.A(_3068_),
    .B(_1451_),
    .X(_2645_));
 sky130_fd_sc_hd__o221a_1 _7508_ (.A1(_3101_),
    .A2(_1484_),
    .B1(_2643_),
    .B2(_2644_),
    .C1(_2645_),
    .X(_2646_));
 sky130_fd_sc_hd__a221o_1 _7509_ (.A1(_3068_),
    .A2(_1451_),
    .B1(_1539_),
    .B2(_2624_),
    .C1(_2646_),
    .X(_2647_));
 sky130_fd_sc_hd__nor2_1 _7510_ (.A(_3328_),
    .B(_0347_),
    .Y(_2648_));
 sky130_fd_sc_hd__a31o_1 _7511_ (.A1(_2623_),
    .A2(_2625_),
    .A3(_2647_),
    .B1(_2648_),
    .X(_2649_));
 sky130_fd_sc_hd__clkbuf_4 _7512_ (.A(_2649_),
    .X(_2651_));
 sky130_fd_sc_hd__clkbuf_4 _7513_ (.A(_2651_),
    .X(_2652_));
 sky130_fd_sc_hd__mux2_2 _7514_ (.A0(_0420_),
    .A1(_0410_),
    .S(_2652_),
    .X(_2653_));
 sky130_fd_sc_hd__mux2_2 _7515_ (.A0(_0348_),
    .A1(_0349_),
    .S(_2651_),
    .X(_2654_));
 sky130_fd_sc_hd__a21o_1 _7516_ (.A1(_0347_),
    .A2(_3635_),
    .B1(_3830_),
    .X(_2655_));
 sky130_fd_sc_hd__and2_1 _7517_ (.A(_0419_),
    .B(_2655_),
    .X(_2656_));
 sky130_fd_sc_hd__mux2_1 _7518_ (.A0(_2656_),
    .A1(_0427_),
    .S(_2651_),
    .X(_2657_));
 sky130_fd_sc_hd__a31o_2 _7519_ (.A1(_2653_),
    .A2(_2654_),
    .A3(_2657_),
    .B1(_0399_),
    .X(_2658_));
 sky130_fd_sc_hd__mux2_2 _7520_ (.A0(_0403_),
    .A1(_0406_),
    .S(_2652_),
    .X(_2659_));
 sky130_fd_sc_hd__a21o_1 _7521_ (.A1(_2654_),
    .A2(_2657_),
    .B1(_0399_),
    .X(_2660_));
 sky130_fd_sc_hd__xnor2_4 _7522_ (.A(_2653_),
    .B(_2660_),
    .Y(_2662_));
 sky130_fd_sc_hd__or2_1 _7523_ (.A(_0399_),
    .B(_2654_),
    .X(_2663_));
 sky130_fd_sc_hd__xnor2_1 _7524_ (.A(_2657_),
    .B(_2663_),
    .Y(_2664_));
 sky130_fd_sc_hd__inv_2 _7525_ (.A(_2664_),
    .Y(_2665_));
 sky130_fd_sc_hd__nand2_1 _7526_ (.A(_2662_),
    .B(_2665_),
    .Y(_2666_));
 sky130_fd_sc_hd__nor2_1 _7527_ (.A(_0385_),
    .B(_2651_),
    .Y(_2667_));
 sky130_fd_sc_hd__a211o_1 _7528_ (.A1(_0388_),
    .A2(_2651_),
    .B1(_2667_),
    .C1(_0386_),
    .X(_2668_));
 sky130_fd_sc_hd__xnor2_1 _7529_ (.A(_0369_),
    .B(_2651_),
    .Y(_2669_));
 sky130_fd_sc_hd__mux2_1 _7530_ (.A0(_2668_),
    .A1(_2669_),
    .S(_0375_),
    .X(_2670_));
 sky130_fd_sc_hd__nor2_1 _7531_ (.A(_0363_),
    .B(_2651_),
    .Y(_2671_));
 sky130_fd_sc_hd__a21oi_2 _7532_ (.A1(_0356_),
    .A2(_2651_),
    .B1(_2671_),
    .Y(_2673_));
 sky130_fd_sc_hd__o2bb2ai_2 _7533_ (.A1_N(_0442_),
    .A2_N(_2670_),
    .B1(_2673_),
    .B2(_0395_),
    .Y(_2674_));
 sky130_fd_sc_hd__xnor2_2 _7534_ (.A(_2346_),
    .B(_2674_),
    .Y(_2675_));
 sky130_fd_sc_hd__xnor2_2 _7535_ (.A(_0442_),
    .B(_2670_),
    .Y(_2676_));
 sky130_fd_sc_hd__xor2_2 _7536_ (.A(_2658_),
    .B(_2659_),
    .X(_2677_));
 sky130_fd_sc_hd__mux2_1 _7537_ (.A0(_0345_),
    .A1(_0342_),
    .S(_2651_),
    .X(_2678_));
 sky130_fd_sc_hd__mux2_1 _7538_ (.A0(_0427_),
    .A1(_2656_),
    .S(_2651_),
    .X(_2679_));
 sky130_fd_sc_hd__inv_2 _7539_ (.A(_2679_),
    .Y(_2680_));
 sky130_fd_sc_hd__nor2_1 _7540_ (.A(_3328_),
    .B(_1781_),
    .Y(_2681_));
 sky130_fd_sc_hd__o21ba_1 _7541_ (.A1(_2678_),
    .A2(_2680_),
    .B1_N(_2681_),
    .X(_2682_));
 sky130_fd_sc_hd__mux2_1 _7542_ (.A0(_0410_),
    .A1(_0420_),
    .S(_2652_),
    .X(_2684_));
 sky130_fd_sc_hd__nor2_1 _7543_ (.A(_2681_),
    .B(_2684_),
    .Y(_2685_));
 sky130_fd_sc_hd__mux2_1 _7544_ (.A0(_0406_),
    .A1(_0403_),
    .S(_2652_),
    .X(_2686_));
 sky130_fd_sc_hd__or3_1 _7545_ (.A(_2682_),
    .B(_2685_),
    .C(_2686_),
    .X(_2687_));
 sky130_fd_sc_hd__o21ai_1 _7546_ (.A1(_2682_),
    .A2(_2685_),
    .B1(_2686_),
    .Y(_2688_));
 sky130_fd_sc_hd__xnor2_1 _7547_ (.A(_2682_),
    .B(_2684_),
    .Y(_2689_));
 sky130_fd_sc_hd__a2bb2o_1 _7548_ (.A1_N(_2654_),
    .A2_N(_2678_),
    .B1(_2674_),
    .B2(_0351_),
    .X(_2690_));
 sky130_fd_sc_hd__or2b_1 _7549_ (.A(_2681_),
    .B_N(_2678_),
    .X(_2691_));
 sky130_fd_sc_hd__xnor2_1 _7550_ (.A(_2691_),
    .B(_2679_),
    .Y(_2692_));
 sky130_fd_sc_hd__a22o_1 _7551_ (.A1(_0433_),
    .A2(_2690_),
    .B1(_2692_),
    .B2(_2665_),
    .X(_2693_));
 sky130_fd_sc_hd__a2bb2o_1 _7552_ (.A1_N(_2662_),
    .A2_N(_2689_),
    .B1(_2693_),
    .B2(_0448_),
    .X(_2695_));
 sky130_fd_sc_hd__a32o_1 _7553_ (.A1(_2677_),
    .A2(_2687_),
    .A3(_2688_),
    .B1(_2695_),
    .B2(_0415_),
    .X(_2696_));
 sky130_fd_sc_hd__xnor2_1 _7554_ (.A(_0416_),
    .B(_2695_),
    .Y(_2697_));
 sky130_fd_sc_hd__nand2_1 _7555_ (.A(_0433_),
    .B(_2690_),
    .Y(_2698_));
 sky130_fd_sc_hd__or2_1 _7556_ (.A(_0433_),
    .B(_2690_),
    .X(_2699_));
 sky130_fd_sc_hd__xnor2_1 _7557_ (.A(_0425_),
    .B(_2693_),
    .Y(_2700_));
 sky130_fd_sc_hd__a21o_1 _7558_ (.A1(_2698_),
    .A2(_2699_),
    .B1(_2700_),
    .X(_2701_));
 sky130_fd_sc_hd__a211oi_4 _7559_ (.A1(_0465_),
    .A2(_2696_),
    .B1(_2697_),
    .C1(_2701_),
    .Y(_2702_));
 sky130_fd_sc_hd__nand2_1 _7560_ (.A(_2676_),
    .B(_2702_),
    .Y(_2703_));
 sky130_fd_sc_hd__buf_2 _7561_ (.A(_2703_),
    .X(_2704_));
 sky130_fd_sc_hd__xor2_2 _7562_ (.A(_0375_),
    .B(_2668_),
    .X(_2706_));
 sky130_fd_sc_hd__and2_1 _7563_ (.A(_2702_),
    .B(_0390_),
    .X(_2707_));
 sky130_fd_sc_hd__buf_2 _7564_ (.A(_2707_),
    .X(_2708_));
 sky130_fd_sc_hd__and3_1 _7565_ (.A(_2319_),
    .B(_2706_),
    .C(_2708_),
    .X(_2709_));
 sky130_fd_sc_hd__or3b_2 _7566_ (.A(_2675_),
    .B(_2704_),
    .C_N(_2709_),
    .X(_2710_));
 sky130_fd_sc_hd__nand2_1 _7567_ (.A(_2319_),
    .B(_2708_),
    .Y(_2711_));
 sky130_fd_sc_hd__nand2_2 _7568_ (.A(_2702_),
    .B(_2706_),
    .Y(_2712_));
 sky130_fd_sc_hd__clkbuf_4 _7569_ (.A(_2652_),
    .X(_2713_));
 sky130_fd_sc_hd__mux2_1 _7570_ (.A0(_0218_),
    .A1(_4222_),
    .S(_2713_),
    .X(_2714_));
 sky130_fd_sc_hd__mux2_1 _7571_ (.A0(_3855_),
    .A1(_3802_),
    .S(_2652_),
    .X(_2715_));
 sky130_fd_sc_hd__or3b_1 _7572_ (.A(_0391_),
    .B(_2715_),
    .C_N(_2702_),
    .X(_2717_));
 sky130_fd_sc_hd__o21ai_1 _7573_ (.A1(_2708_),
    .A2(_2714_),
    .B1(_2717_),
    .Y(_2718_));
 sky130_fd_sc_hd__o22a_1 _7574_ (.A1(_2706_),
    .A2(_2711_),
    .B1(_2712_),
    .B2(_2718_),
    .X(_2719_));
 sky130_fd_sc_hd__or2_1 _7575_ (.A(_2704_),
    .B(_2719_),
    .X(_2720_));
 sky130_fd_sc_hd__buf_4 _7576_ (.A(_2713_),
    .X(_2721_));
 sky130_fd_sc_hd__mux2_1 _7577_ (.A0(_3802_),
    .A1(_4217_),
    .S(_2721_),
    .X(_2722_));
 sky130_fd_sc_hd__or3_1 _7578_ (.A(_2675_),
    .B(_2720_),
    .C(_2722_),
    .X(_2723_));
 sky130_fd_sc_hd__o21a_1 _7579_ (.A1(_2675_),
    .A2(_2720_),
    .B1(_2722_),
    .X(_2724_));
 sky130_fd_sc_hd__inv_2 _7580_ (.A(_2724_),
    .Y(_2725_));
 sky130_fd_sc_hd__nand2_1 _7581_ (.A(_2723_),
    .B(_2725_),
    .Y(_2726_));
 sky130_fd_sc_hd__inv_2 _7582_ (.A(_2726_),
    .Y(_2728_));
 sky130_fd_sc_hd__inv_2 _7583_ (.A(_2675_),
    .Y(_2729_));
 sky130_fd_sc_hd__and2_1 _7584_ (.A(_2702_),
    .B(_2706_),
    .X(_2730_));
 sky130_fd_sc_hd__buf_2 _7585_ (.A(_2730_),
    .X(_2731_));
 sky130_fd_sc_hd__mux2_1 _7586_ (.A0(_2319_),
    .A1(_2714_),
    .S(_2707_),
    .X(_2732_));
 sky130_fd_sc_hd__mux2_1 _7587_ (.A0(_4153_),
    .A1(_0113_),
    .S(_2652_),
    .X(_2733_));
 sky130_fd_sc_hd__mux2_1 _7588_ (.A0(_2715_),
    .A1(_2733_),
    .S(_2707_),
    .X(_2734_));
 sky130_fd_sc_hd__or2_1 _7589_ (.A(_2712_),
    .B(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__o21ai_1 _7590_ (.A1(_2731_),
    .A2(_2732_),
    .B1(_2735_),
    .Y(_2736_));
 sky130_fd_sc_hd__nor2_1 _7591_ (.A(_2704_),
    .B(_2736_),
    .Y(_2737_));
 sky130_fd_sc_hd__nand2_1 _7592_ (.A(_2729_),
    .B(_2737_),
    .Y(_2739_));
 sky130_fd_sc_hd__mux2_2 _7593_ (.A0(_0113_),
    .A1(_4153_),
    .S(_2721_),
    .X(_2740_));
 sky130_fd_sc_hd__xnor2_1 _7594_ (.A(_2739_),
    .B(_2740_),
    .Y(_2741_));
 sky130_fd_sc_hd__and2_1 _7595_ (.A(_2729_),
    .B(_2702_),
    .X(_2742_));
 sky130_fd_sc_hd__clkbuf_4 _7596_ (.A(_2742_),
    .X(_2743_));
 sky130_fd_sc_hd__mux2_1 _7597_ (.A0(_1355_),
    .A1(_3881_),
    .S(_2713_),
    .X(_2744_));
 sky130_fd_sc_hd__mux2_1 _7598_ (.A0(_2733_),
    .A1(_2744_),
    .S(_2708_),
    .X(_2745_));
 sky130_fd_sc_hd__nor2_1 _7599_ (.A(_2712_),
    .B(_2745_),
    .Y(_2746_));
 sky130_fd_sc_hd__a21oi_1 _7600_ (.A1(_2712_),
    .A2(_2718_),
    .B1(_2746_),
    .Y(_2747_));
 sky130_fd_sc_hd__and2_2 _7601_ (.A(_2676_),
    .B(_2702_),
    .X(_2748_));
 sky130_fd_sc_hd__mux2_1 _7602_ (.A0(_2709_),
    .A1(_2747_),
    .S(_2748_),
    .X(_2750_));
 sky130_fd_sc_hd__and2_1 _7603_ (.A(_2743_),
    .B(_2750_),
    .X(_2751_));
 sky130_fd_sc_hd__mux2_1 _7604_ (.A0(_3881_),
    .A1(_1355_),
    .S(_2721_),
    .X(_2752_));
 sky130_fd_sc_hd__nand2_1 _7605_ (.A(_2731_),
    .B(_2732_),
    .Y(_2753_));
 sky130_fd_sc_hd__mux2_1 _7606_ (.A0(_3986_),
    .A1(_3901_),
    .S(_2652_),
    .X(_2754_));
 sky130_fd_sc_hd__mux2_1 _7607_ (.A0(_2744_),
    .A1(_2754_),
    .S(_2708_),
    .X(_2755_));
 sky130_fd_sc_hd__mux2_1 _7608_ (.A0(_2734_),
    .A1(_2755_),
    .S(_2731_),
    .X(_2756_));
 sky130_fd_sc_hd__a2bb2o_1 _7609_ (.A1_N(_2676_),
    .A2_N(_2753_),
    .B1(_2756_),
    .B2(_2748_),
    .X(_2757_));
 sky130_fd_sc_hd__nand2_1 _7610_ (.A(_2743_),
    .B(_2757_),
    .Y(_2758_));
 sky130_fd_sc_hd__mux2_1 _7611_ (.A0(_3816_),
    .A1(_1384_),
    .S(_2721_),
    .X(_2759_));
 sky130_fd_sc_hd__and2_1 _7612_ (.A(_2758_),
    .B(_2759_),
    .X(_2761_));
 sky130_fd_sc_hd__nand2_2 _7613_ (.A(_2729_),
    .B(_2702_),
    .Y(_2762_));
 sky130_fd_sc_hd__mux2_1 _7614_ (.A0(_0147_),
    .A1(_4045_),
    .S(_2652_),
    .X(_2763_));
 sky130_fd_sc_hd__mux2_1 _7615_ (.A0(_2754_),
    .A1(_2763_),
    .S(_2707_),
    .X(_2764_));
 sky130_fd_sc_hd__or2_1 _7616_ (.A(_2712_),
    .B(_2764_),
    .X(_2765_));
 sky130_fd_sc_hd__o21ai_1 _7617_ (.A1(_2731_),
    .A2(_2745_),
    .B1(_2765_),
    .Y(_2766_));
 sky130_fd_sc_hd__mux2_1 _7618_ (.A0(_2719_),
    .A1(_2766_),
    .S(_2748_),
    .X(_2767_));
 sky130_fd_sc_hd__or2_1 _7619_ (.A(_2762_),
    .B(_2767_),
    .X(_2768_));
 sky130_fd_sc_hd__mux2_1 _7620_ (.A0(_4045_),
    .A1(_0147_),
    .S(_2721_),
    .X(_2769_));
 sky130_fd_sc_hd__or2_1 _7621_ (.A(_2768_),
    .B(_2769_),
    .X(_2770_));
 sky130_fd_sc_hd__nand2_1 _7622_ (.A(_2768_),
    .B(_2769_),
    .Y(_2772_));
 sky130_fd_sc_hd__nand2_1 _7623_ (.A(_2770_),
    .B(_2772_),
    .Y(_2773_));
 sky130_fd_sc_hd__mux2_1 _7624_ (.A0(_3883_),
    .A1(_3776_),
    .S(_2652_),
    .X(_2774_));
 sky130_fd_sc_hd__mux2_1 _7625_ (.A0(_2763_),
    .A1(_2774_),
    .S(_2707_),
    .X(_2775_));
 sky130_fd_sc_hd__or2_1 _7626_ (.A(_2712_),
    .B(_2775_),
    .X(_2776_));
 sky130_fd_sc_hd__o21ai_1 _7627_ (.A1(_2731_),
    .A2(_2755_),
    .B1(_2776_),
    .Y(_2777_));
 sky130_fd_sc_hd__mux2_1 _7628_ (.A0(_2736_),
    .A1(_2777_),
    .S(_2748_),
    .X(_2778_));
 sky130_fd_sc_hd__nor2_1 _7629_ (.A(_2762_),
    .B(_2778_),
    .Y(_2779_));
 sky130_fd_sc_hd__mux2_1 _7630_ (.A0(_3793_),
    .A1(_3795_),
    .S(_2713_),
    .X(_2780_));
 sky130_fd_sc_hd__inv_2 _7631_ (.A(_2780_),
    .Y(_2781_));
 sky130_fd_sc_hd__nand2_1 _7632_ (.A(_2779_),
    .B(_2781_),
    .Y(_2783_));
 sky130_fd_sc_hd__mux2_1 _7633_ (.A0(_3868_),
    .A1(_3893_),
    .S(_2713_),
    .X(_2784_));
 sky130_fd_sc_hd__mux2_1 _7634_ (.A0(_2774_),
    .A1(_2784_),
    .S(_2708_),
    .X(_2785_));
 sky130_fd_sc_hd__mux2_1 _7635_ (.A0(_2764_),
    .A1(_2785_),
    .S(_2731_),
    .X(_2786_));
 sky130_fd_sc_hd__o221a_1 _7636_ (.A1(_2676_),
    .A2(_2747_),
    .B1(_2786_),
    .B2(_2704_),
    .C1(_2743_),
    .X(_2787_));
 sky130_fd_sc_hd__a31o_1 _7637_ (.A1(_2675_),
    .A2(_2748_),
    .A3(_2709_),
    .B1(_2787_),
    .X(_2788_));
 sky130_fd_sc_hd__mux2_1 _7638_ (.A0(_3893_),
    .A1(_3868_),
    .S(_2713_),
    .X(_2789_));
 sky130_fd_sc_hd__and2_1 _7639_ (.A(_2788_),
    .B(_2789_),
    .X(_2790_));
 sky130_fd_sc_hd__mux2_1 _7640_ (.A0(_1531_),
    .A1(_3878_),
    .S(_2713_),
    .X(_2791_));
 sky130_fd_sc_hd__mux2_1 _7641_ (.A0(_2784_),
    .A1(_2791_),
    .S(_2708_),
    .X(_2792_));
 sky130_fd_sc_hd__mux2_1 _7642_ (.A0(_2775_),
    .A1(_2792_),
    .S(_2731_),
    .X(_2794_));
 sky130_fd_sc_hd__mux2_1 _7643_ (.A0(_2756_),
    .A1(_2794_),
    .S(_2748_),
    .X(_2795_));
 sky130_fd_sc_hd__or2_1 _7644_ (.A(_2762_),
    .B(_2795_),
    .X(_2796_));
 sky130_fd_sc_hd__and3_1 _7645_ (.A(_2676_),
    .B(_2731_),
    .C(_2732_),
    .X(_2797_));
 sky130_fd_sc_hd__or2_1 _7646_ (.A(_2742_),
    .B(_2797_),
    .X(_2798_));
 sky130_fd_sc_hd__nand2_1 _7647_ (.A(_2796_),
    .B(_2798_),
    .Y(_2799_));
 sky130_fd_sc_hd__mux2_1 _7648_ (.A0(_3771_),
    .A1(_3703_),
    .S(_2713_),
    .X(_2800_));
 sky130_fd_sc_hd__nor2_1 _7649_ (.A(_2799_),
    .B(_2800_),
    .Y(_2801_));
 sky130_fd_sc_hd__mux2_1 _7650_ (.A0(_3845_),
    .A1(_4126_),
    .S(_2713_),
    .X(_2802_));
 sky130_fd_sc_hd__mux2_1 _7651_ (.A0(_3726_),
    .A1(_3845_),
    .S(_2713_),
    .X(_2803_));
 sky130_fd_sc_hd__nand2_1 _7652_ (.A(_2708_),
    .B(_2803_),
    .Y(_2805_));
 sky130_fd_sc_hd__o21ai_1 _7653_ (.A1(_2708_),
    .A2(_2791_),
    .B1(_2805_),
    .Y(_2806_));
 sky130_fd_sc_hd__nand2_1 _7654_ (.A(_2712_),
    .B(_2785_),
    .Y(_2807_));
 sky130_fd_sc_hd__o21ai_1 _7655_ (.A1(_2712_),
    .A2(_2806_),
    .B1(_2807_),
    .Y(_2808_));
 sky130_fd_sc_hd__nand2_1 _7656_ (.A(_2704_),
    .B(_2766_),
    .Y(_2809_));
 sky130_fd_sc_hd__o211a_1 _7657_ (.A1(_2704_),
    .A2(_2808_),
    .B1(_2809_),
    .C1(_2742_),
    .X(_2810_));
 sky130_fd_sc_hd__o21bai_1 _7658_ (.A1(_2729_),
    .A2(_2720_),
    .B1_N(_2810_),
    .Y(_2811_));
 sky130_fd_sc_hd__and2b_1 _7659_ (.A_N(_2802_),
    .B(_2811_),
    .X(_2812_));
 sky130_fd_sc_hd__nand2_1 _7660_ (.A(_2799_),
    .B(_2800_),
    .Y(_2813_));
 sky130_fd_sc_hd__o21a_1 _7661_ (.A1(_2801_),
    .A2(_2812_),
    .B1(_2813_),
    .X(_2814_));
 sky130_fd_sc_hd__nor2_1 _7662_ (.A(_2788_),
    .B(_2789_),
    .Y(_2816_));
 sky130_fd_sc_hd__o21bai_1 _7663_ (.A1(_2790_),
    .A2(_2814_),
    .B1_N(_2816_),
    .Y(_2817_));
 sky130_fd_sc_hd__or2_1 _7664_ (.A(_2779_),
    .B(_2781_),
    .X(_2818_));
 sky130_fd_sc_hd__a21boi_1 _7665_ (.A1(_2783_),
    .A2(_2817_),
    .B1_N(_2818_),
    .Y(_2819_));
 sky130_fd_sc_hd__and2b_1 _7666_ (.A_N(_2768_),
    .B(_2769_),
    .X(_2820_));
 sky130_fd_sc_hd__a21oi_1 _7667_ (.A1(_2773_),
    .A2(_2819_),
    .B1(_2820_),
    .Y(_2821_));
 sky130_fd_sc_hd__or2_1 _7668_ (.A(_2758_),
    .B(_2759_),
    .X(_2822_));
 sky130_fd_sc_hd__o21a_1 _7669_ (.A1(_2761_),
    .A2(_2821_),
    .B1(_2822_),
    .X(_2823_));
 sky130_fd_sc_hd__nand2_1 _7670_ (.A(_2743_),
    .B(_2750_),
    .Y(_2824_));
 sky130_fd_sc_hd__or2_1 _7671_ (.A(_2824_),
    .B(_2752_),
    .X(_2825_));
 sky130_fd_sc_hd__and2_1 _7672_ (.A(_2824_),
    .B(_2752_),
    .X(_2827_));
 sky130_fd_sc_hd__inv_2 _7673_ (.A(_2827_),
    .Y(_2828_));
 sky130_fd_sc_hd__nand2_1 _7674_ (.A(_2825_),
    .B(_2828_),
    .Y(_2829_));
 sky130_fd_sc_hd__or2b_1 _7675_ (.A(_2823_),
    .B_N(_2829_),
    .X(_2830_));
 sky130_fd_sc_hd__a21bo_1 _7676_ (.A1(_2751_),
    .A2(_2752_),
    .B1_N(_2830_),
    .X(_2831_));
 sky130_fd_sc_hd__and3_1 _7677_ (.A(_2729_),
    .B(_2737_),
    .C(_2740_),
    .X(_2832_));
 sky130_fd_sc_hd__a21oi_1 _7678_ (.A1(_2741_),
    .A2(_2831_),
    .B1(_2832_),
    .Y(_2833_));
 sky130_fd_sc_hd__or3b_1 _7679_ (.A(_2675_),
    .B(_2720_),
    .C_N(_2722_),
    .X(_2834_));
 sky130_fd_sc_hd__o21ai_1 _7680_ (.A1(_2728_),
    .A2(_2833_),
    .B1(_2834_),
    .Y(_2835_));
 sky130_fd_sc_hd__nand2_1 _7681_ (.A(_2743_),
    .B(_2797_),
    .Y(_2836_));
 sky130_fd_sc_hd__mux2_1 _7682_ (.A0(_3925_),
    .A1(_0080_),
    .S(_2721_),
    .X(_2838_));
 sky130_fd_sc_hd__nand2_1 _7683_ (.A(_2836_),
    .B(_2838_),
    .Y(_2839_));
 sky130_fd_sc_hd__nor2_1 _7684_ (.A(_2836_),
    .B(_2838_),
    .Y(_2840_));
 sky130_fd_sc_hd__a21oi_2 _7685_ (.A1(_2835_),
    .A2(_2839_),
    .B1(_2840_),
    .Y(_2841_));
 sky130_fd_sc_hd__a21oi_4 _7686_ (.A1(_2710_),
    .A2(_2841_),
    .B1(_1297_),
    .Y(_2842_));
 sky130_fd_sc_hd__a21bo_1 _7687_ (.A1(_4250_),
    .A2(_0082_),
    .B1_N(_2710_),
    .X(_2843_));
 sky130_fd_sc_hd__and2b_1 _7688_ (.A_N(_2840_),
    .B(_2839_),
    .X(_2844_));
 sky130_fd_sc_hd__or2b_1 _7689_ (.A(_2761_),
    .B_N(_2822_),
    .X(_2845_));
 sky130_fd_sc_hd__nand2_1 _7690_ (.A(_2783_),
    .B(_2818_),
    .Y(_2846_));
 sky130_fd_sc_hd__inv_2 _7691_ (.A(_2846_),
    .Y(_2847_));
 sky130_fd_sc_hd__or2_1 _7692_ (.A(_2790_),
    .B(_2816_),
    .X(_2849_));
 sky130_fd_sc_hd__and2b_1 _7693_ (.A_N(_2801_),
    .B(_2813_),
    .X(_2850_));
 sky130_fd_sc_hd__nor2_1 _7694_ (.A(_2811_),
    .B(_2802_),
    .Y(_2851_));
 sky130_fd_sc_hd__nor2_1 _7695_ (.A(_2708_),
    .B(_2803_),
    .Y(_2852_));
 sky130_fd_sc_hd__mux2_1 _7696_ (.A0(_2792_),
    .A1(_2852_),
    .S(_2731_),
    .X(_2853_));
 sky130_fd_sc_hd__nor2_1 _7697_ (.A(_2704_),
    .B(_2853_),
    .Y(_2854_));
 sky130_fd_sc_hd__a21oi_1 _7698_ (.A1(_2704_),
    .A2(_2777_),
    .B1(_2854_),
    .Y(_2855_));
 sky130_fd_sc_hd__a22o_1 _7699_ (.A1(_2675_),
    .A2(_2737_),
    .B1(_2855_),
    .B2(_2743_),
    .X(_2856_));
 sky130_fd_sc_hd__nor2_1 _7700_ (.A(_2676_),
    .B(_2762_),
    .Y(_2857_));
 sky130_fd_sc_hd__o2bb2a_1 _7701_ (.A1_N(_2808_),
    .A2_N(_2857_),
    .B1(_2742_),
    .B2(_2767_),
    .X(_2858_));
 sky130_fd_sc_hd__o2bb2a_1 _7702_ (.A1_N(_2853_),
    .A2_N(_2857_),
    .B1(_2742_),
    .B2(_2778_),
    .X(_2860_));
 sky130_fd_sc_hd__nand2_1 _7703_ (.A(_2858_),
    .B(_2860_),
    .Y(_2861_));
 sky130_fd_sc_hd__nor2_1 _7704_ (.A(_2703_),
    .B(_2706_),
    .Y(_2862_));
 sky130_fd_sc_hd__a221o_1 _7705_ (.A1(_2704_),
    .A2(_2794_),
    .B1(_2852_),
    .B2(_2862_),
    .C1(_2762_),
    .X(_2863_));
 sky130_fd_sc_hd__o21ai_2 _7706_ (.A1(_2743_),
    .A2(_2757_),
    .B1(_2863_),
    .Y(_2864_));
 sky130_fd_sc_hd__and2b_1 _7707_ (.A_N(_2806_),
    .B(_2862_),
    .X(_2865_));
 sky130_fd_sc_hd__a211o_1 _7708_ (.A1(_2704_),
    .A2(_2786_),
    .B1(_2865_),
    .C1(_2762_),
    .X(_2866_));
 sky130_fd_sc_hd__o21ai_2 _7709_ (.A1(_2743_),
    .A2(_2750_),
    .B1(_2866_),
    .Y(_2867_));
 sky130_fd_sc_hd__nand3b_1 _7710_ (.A_N(_2861_),
    .B(_2864_),
    .C(_2867_),
    .Y(_2868_));
 sky130_fd_sc_hd__nor2_1 _7711_ (.A(_2856_),
    .B(_2868_),
    .Y(_2869_));
 sky130_fd_sc_hd__and2_1 _7712_ (.A(_2811_),
    .B(_2802_),
    .X(_2871_));
 sky130_fd_sc_hd__o21bai_1 _7713_ (.A1(_2851_),
    .A2(_2869_),
    .B1_N(_2871_),
    .Y(_2872_));
 sky130_fd_sc_hd__a21o_1 _7714_ (.A1(_2796_),
    .A2(_2798_),
    .B1(_2800_),
    .X(_2873_));
 sky130_fd_sc_hd__o21ai_1 _7715_ (.A1(_2850_),
    .A2(_2872_),
    .B1(_2873_),
    .Y(_2874_));
 sky130_fd_sc_hd__and2b_1 _7716_ (.A_N(_2788_),
    .B(_2789_),
    .X(_2875_));
 sky130_fd_sc_hd__a21oi_1 _7717_ (.A1(_2849_),
    .A2(_2874_),
    .B1(_2875_),
    .Y(_2876_));
 sky130_fd_sc_hd__or2_1 _7718_ (.A(_2779_),
    .B(_2780_),
    .X(_2877_));
 sky130_fd_sc_hd__o21ai_1 _7719_ (.A1(_2847_),
    .A2(_2876_),
    .B1(_2877_),
    .Y(_2878_));
 sky130_fd_sc_hd__and2_1 _7720_ (.A(_2768_),
    .B(_2769_),
    .X(_2879_));
 sky130_fd_sc_hd__a21o_1 _7721_ (.A1(_2770_),
    .A2(_2878_),
    .B1(_2879_),
    .X(_2880_));
 sky130_fd_sc_hd__a21oi_1 _7722_ (.A1(_2743_),
    .A2(_2757_),
    .B1(_2759_),
    .Y(_2882_));
 sky130_fd_sc_hd__a21o_1 _7723_ (.A1(_2845_),
    .A2(_2880_),
    .B1(_2882_),
    .X(_2883_));
 sky130_fd_sc_hd__a221o_1 _7724_ (.A1(_2739_),
    .A2(_2740_),
    .B1(_2825_),
    .B2(_2883_),
    .C1(_2827_),
    .X(_2884_));
 sky130_fd_sc_hd__o21a_1 _7725_ (.A1(_2739_),
    .A2(_2740_),
    .B1(_2884_),
    .X(_2885_));
 sky130_fd_sc_hd__a21oi_1 _7726_ (.A1(_2723_),
    .A2(_2885_),
    .B1(_2724_),
    .Y(_2886_));
 sky130_fd_sc_hd__a21o_1 _7727_ (.A1(_2743_),
    .A2(_2797_),
    .B1(_2838_),
    .X(_2887_));
 sky130_fd_sc_hd__o211a_1 _7728_ (.A1(_2844_),
    .A2(_2886_),
    .B1(_2887_),
    .C1(_1286_),
    .X(_2888_));
 sky130_fd_sc_hd__o21bai_1 _7729_ (.A1(_1297_),
    .A2(_2841_),
    .B1_N(_2888_),
    .Y(_2889_));
 sky130_fd_sc_hd__xor2_1 _7730_ (.A(_2843_),
    .B(_2889_),
    .X(_2890_));
 sky130_fd_sc_hd__or2b_1 _7731_ (.A(_2842_),
    .B_N(_2890_),
    .X(_2891_));
 sky130_fd_sc_hd__mux2_1 _7732_ (.A0(_2835_),
    .A1(_2886_),
    .S(_1297_),
    .X(_2893_));
 sky130_fd_sc_hd__xnor2_1 _7733_ (.A(_2844_),
    .B(_2893_),
    .Y(_2894_));
 sky130_fd_sc_hd__or2b_1 _7734_ (.A(_2891_),
    .B_N(_2894_),
    .X(_2895_));
 sky130_fd_sc_hd__a21oi_1 _7735_ (.A1(_2825_),
    .A2(_2883_),
    .B1(_2827_),
    .Y(_2896_));
 sky130_fd_sc_hd__mux2_1 _7736_ (.A0(_2831_),
    .A1(_2896_),
    .S(_1286_),
    .X(_2897_));
 sky130_fd_sc_hd__xnor2_1 _7737_ (.A(_2741_),
    .B(_2897_),
    .Y(_2898_));
 sky130_fd_sc_hd__inv_2 _7738_ (.A(_2898_),
    .Y(_2899_));
 sky130_fd_sc_hd__mux2_1 _7739_ (.A0(_2833_),
    .A1(_2885_),
    .S(_1297_),
    .X(_2900_));
 sky130_fd_sc_hd__xnor2_1 _7740_ (.A(_2726_),
    .B(_2900_),
    .Y(_2901_));
 sky130_fd_sc_hd__or2_1 _7741_ (.A(_2899_),
    .B(_2901_),
    .X(_2902_));
 sky130_fd_sc_hd__or2_1 _7742_ (.A(_2895_),
    .B(_2902_),
    .X(_2904_));
 sky130_fd_sc_hd__mux2_1 _7743_ (.A0(_2823_),
    .A1(_2883_),
    .S(_1297_),
    .X(_2905_));
 sky130_fd_sc_hd__xnor2_2 _7744_ (.A(_2829_),
    .B(_2905_),
    .Y(_2906_));
 sky130_fd_sc_hd__mux2_1 _7745_ (.A0(_2821_),
    .A1(_2880_),
    .S(_1297_),
    .X(_2907_));
 sky130_fd_sc_hd__xor2_2 _7746_ (.A(_2845_),
    .B(_2907_),
    .X(_2908_));
 sky130_fd_sc_hd__nor2_1 _7747_ (.A(_1297_),
    .B(_2819_),
    .Y(_2909_));
 sky130_fd_sc_hd__a21oi_1 _7748_ (.A1(_1297_),
    .A2(_2878_),
    .B1(_2909_),
    .Y(_2910_));
 sky130_fd_sc_hd__xor2_2 _7749_ (.A(_2773_),
    .B(_2910_),
    .X(_2911_));
 sky130_fd_sc_hd__clkinv_2 _7750_ (.A(_2817_),
    .Y(_2912_));
 sky130_fd_sc_hd__mux2_1 _7751_ (.A0(_2912_),
    .A1(_2876_),
    .S(_1297_),
    .X(_2913_));
 sky130_fd_sc_hd__xnor2_2 _7752_ (.A(_2846_),
    .B(_2913_),
    .Y(_2915_));
 sky130_fd_sc_hd__or2_1 _7753_ (.A(_2911_),
    .B(_2915_),
    .X(_2916_));
 sky130_fd_sc_hd__or3_1 _7754_ (.A(_2906_),
    .B(_2908_),
    .C(_2916_),
    .X(_2917_));
 sky130_fd_sc_hd__or2_2 _7755_ (.A(_2904_),
    .B(_2917_),
    .X(_2918_));
 sky130_fd_sc_hd__nor2_1 _7756_ (.A(_1308_),
    .B(_2814_),
    .Y(_2919_));
 sky130_fd_sc_hd__a21oi_1 _7757_ (.A1(_1308_),
    .A2(_2874_),
    .B1(_2919_),
    .Y(_2920_));
 sky130_fd_sc_hd__xor2_2 _7758_ (.A(_2849_),
    .B(_2920_),
    .X(_2921_));
 sky130_fd_sc_hd__mux2_1 _7759_ (.A0(_2812_),
    .A1(_2872_),
    .S(_1308_),
    .X(_2922_));
 sky130_fd_sc_hd__xor2_2 _7760_ (.A(_2850_),
    .B(_2922_),
    .X(_2923_));
 sky130_fd_sc_hd__inv_2 _7761_ (.A(_2923_),
    .Y(_2924_));
 sky130_fd_sc_hd__nand2_1 _7762_ (.A(_2921_),
    .B(_2924_),
    .Y(_2926_));
 sky130_fd_sc_hd__and2_1 _7763_ (.A(_1308_),
    .B(_2868_),
    .X(_2927_));
 sky130_fd_sc_hd__xnor2_1 _7764_ (.A(_2856_),
    .B(_2927_),
    .Y(_2928_));
 sky130_fd_sc_hd__xnor2_2 _7765_ (.A(_1253_),
    .B(_1275_),
    .Y(_2929_));
 sky130_fd_sc_hd__or4_1 _7766_ (.A(_2929_),
    .B(_2851_),
    .C(_2871_),
    .D(_2869_),
    .X(_2930_));
 sky130_fd_sc_hd__o22ai_1 _7767_ (.A1(_2851_),
    .A2(_2871_),
    .B1(_2869_),
    .B2(_2929_),
    .Y(_2931_));
 sky130_fd_sc_hd__nand2_1 _7768_ (.A(_2930_),
    .B(_2931_),
    .Y(_2932_));
 sky130_fd_sc_hd__inv_2 _7769_ (.A(_2932_),
    .Y(_2933_));
 sky130_fd_sc_hd__nand2_1 _7770_ (.A(_2928_),
    .B(_2933_),
    .Y(_2934_));
 sky130_fd_sc_hd__nor2_1 _7771_ (.A(_2926_),
    .B(_2934_),
    .Y(_2935_));
 sky130_fd_sc_hd__nor2_4 _7772_ (.A(_2918_),
    .B(_2935_),
    .Y(_2937_));
 sky130_fd_sc_hd__or2_1 _7773_ (.A(_2654_),
    .B(_2937_),
    .X(_2938_));
 sky130_fd_sc_hd__nor2_1 _7774_ (.A(_2665_),
    .B(_2938_),
    .Y(_2939_));
 sky130_fd_sc_hd__a21oi_1 _7775_ (.A1(_2868_),
    .A2(_2935_),
    .B1(_2917_),
    .Y(_2940_));
 sky130_fd_sc_hd__nor2_2 _7776_ (.A(_2904_),
    .B(_2940_),
    .Y(_2941_));
 sky130_fd_sc_hd__or2_1 _7777_ (.A(_2673_),
    .B(_2941_),
    .X(_2942_));
 sky130_fd_sc_hd__nand2_1 _7778_ (.A(_2654_),
    .B(_2937_),
    .Y(_2943_));
 sky130_fd_sc_hd__and2_1 _7779_ (.A(_2938_),
    .B(_2943_),
    .X(_2944_));
 sky130_fd_sc_hd__and2b_1 _7780_ (.A_N(_2942_),
    .B(_2944_),
    .X(_2945_));
 sky130_fd_sc_hd__a31o_1 _7781_ (.A1(_2858_),
    .A2(_2860_),
    .A3(_2864_),
    .B1(_2929_),
    .X(_2946_));
 sky130_fd_sc_hd__xnor2_1 _7782_ (.A(_2867_),
    .B(_2946_),
    .Y(_2948_));
 sky130_fd_sc_hd__nand2_1 _7783_ (.A(_1308_),
    .B(_2861_),
    .Y(_2949_));
 sky130_fd_sc_hd__xnor2_1 _7784_ (.A(_2864_),
    .B(_2949_),
    .Y(_2950_));
 sky130_fd_sc_hd__a31oi_2 _7785_ (.A1(_2861_),
    .A2(_2948_),
    .A3(_2950_),
    .B1(_2934_),
    .Y(_2951_));
 sky130_fd_sc_hd__nor2_1 _7786_ (.A(_2906_),
    .B(_2908_),
    .Y(_2952_));
 sky130_fd_sc_hd__a21oi_1 _7787_ (.A1(_2952_),
    .A2(_2916_),
    .B1(_2902_),
    .Y(_2953_));
 sky130_fd_sc_hd__o32ai_4 _7788_ (.A1(_2918_),
    .A2(_2926_),
    .A3(_2951_),
    .B1(_2953_),
    .B2(_2895_),
    .Y(_2954_));
 sky130_fd_sc_hd__mux2_1 _7789_ (.A0(_0370_),
    .A1(_2340_),
    .S(_2721_),
    .X(_2955_));
 sky130_fd_sc_hd__or2b_1 _7790_ (.A(_2954_),
    .B_N(_2955_),
    .X(_2956_));
 sky130_fd_sc_hd__nand2_1 _7791_ (.A(_2673_),
    .B(_2941_),
    .Y(_2957_));
 sky130_fd_sc_hd__nand2_1 _7792_ (.A(_2942_),
    .B(_2957_),
    .Y(_2959_));
 sky130_fd_sc_hd__nor2_1 _7793_ (.A(_2956_),
    .B(_2959_),
    .Y(_2960_));
 sky130_fd_sc_hd__xor2_1 _7794_ (.A(_2954_),
    .B(_2955_),
    .X(_2961_));
 sky130_fd_sc_hd__a21o_1 _7795_ (.A1(_0388_),
    .A2(_2721_),
    .B1(_2667_),
    .X(_2962_));
 sky130_fd_sc_hd__nor2_1 _7796_ (.A(_2928_),
    .B(_2932_),
    .Y(_2963_));
 sky130_fd_sc_hd__o21a_1 _7797_ (.A1(_2923_),
    .A2(_2963_),
    .B1(_2921_),
    .X(_2964_));
 sky130_fd_sc_hd__inv_2 _7798_ (.A(_2911_),
    .Y(_2965_));
 sky130_fd_sc_hd__a21oi_1 _7799_ (.A1(_2965_),
    .A2(_2915_),
    .B1(_2908_),
    .Y(_2966_));
 sky130_fd_sc_hd__o21a_1 _7800_ (.A1(_2898_),
    .A2(_2901_),
    .B1(_2894_),
    .X(_2967_));
 sky130_fd_sc_hd__o32ai_1 _7801_ (.A1(_2904_),
    .A2(_2906_),
    .A3(_2966_),
    .B1(_2967_),
    .B2(_2891_),
    .Y(_2968_));
 sky130_fd_sc_hd__mux2_1 _7802_ (.A0(_2964_),
    .A1(_2968_),
    .S(_2918_),
    .X(_2970_));
 sky130_fd_sc_hd__clkbuf_4 _7803_ (.A(_2970_),
    .X(_2971_));
 sky130_fd_sc_hd__and2b_1 _7804_ (.A_N(_2962_),
    .B(_2971_),
    .X(_2972_));
 sky130_fd_sc_hd__xor2_1 _7805_ (.A(_2962_),
    .B(_2971_),
    .X(_2973_));
 sky130_fd_sc_hd__nand2_1 _7806_ (.A(_2842_),
    .B(_2973_),
    .Y(_2974_));
 sky130_fd_sc_hd__xnor2_1 _7807_ (.A(_2961_),
    .B(_2972_),
    .Y(_2975_));
 sky130_fd_sc_hd__o22a_1 _7808_ (.A1(_2961_),
    .A2(_2972_),
    .B1(_2974_),
    .B2(_2975_),
    .X(_2976_));
 sky130_fd_sc_hd__and2_1 _7809_ (.A(_2956_),
    .B(_2959_),
    .X(_2977_));
 sky130_fd_sc_hd__or2_1 _7810_ (.A(_2960_),
    .B(_2977_),
    .X(_2978_));
 sky130_fd_sc_hd__nor2_1 _7811_ (.A(_2976_),
    .B(_2978_),
    .Y(_2979_));
 sky130_fd_sc_hd__xnor2_1 _7812_ (.A(_2942_),
    .B(_2944_),
    .Y(_2981_));
 sky130_fd_sc_hd__o21a_1 _7813_ (.A1(_2960_),
    .A2(_2979_),
    .B1(_2981_),
    .X(_2982_));
 sky130_fd_sc_hd__and2_1 _7814_ (.A(_2665_),
    .B(_2938_),
    .X(_2983_));
 sky130_fd_sc_hd__nor2_1 _7815_ (.A(_2939_),
    .B(_2983_),
    .Y(_2984_));
 sky130_fd_sc_hd__o21a_1 _7816_ (.A1(_2945_),
    .A2(_2982_),
    .B1(_2984_),
    .X(_2985_));
 sky130_fd_sc_hd__xnor2_1 _7817_ (.A(_2662_),
    .B(_2664_),
    .Y(_2986_));
 sky130_fd_sc_hd__o21ai_1 _7818_ (.A1(_2939_),
    .A2(_2985_),
    .B1(_2986_),
    .Y(_2987_));
 sky130_fd_sc_hd__xnor2_1 _7819_ (.A(_2662_),
    .B(_2677_),
    .Y(_2988_));
 sky130_fd_sc_hd__a21oi_2 _7820_ (.A1(_2666_),
    .A2(_2987_),
    .B1(_2988_),
    .Y(_2989_));
 sky130_fd_sc_hd__nor2_1 _7821_ (.A(_2980_),
    .B(_0347_),
    .Y(_2990_));
 sky130_fd_sc_hd__o22ai_2 _7822_ (.A1(_2990_),
    .A2(_2659_),
    .B1(_2677_),
    .B2(_2662_),
    .Y(_2992_));
 sky130_fd_sc_hd__o22ai_4 _7823_ (.A1(_2658_),
    .A2(_2659_),
    .B1(_2989_),
    .B2(_2992_),
    .Y(_2993_));
 sky130_fd_sc_hd__nor3_1 _7824_ (.A(_2981_),
    .B(_2960_),
    .C(_2979_),
    .Y(_2994_));
 sky130_fd_sc_hd__nor2_1 _7825_ (.A(_2982_),
    .B(_2994_),
    .Y(_2995_));
 sky130_fd_sc_hd__or2_1 _7826_ (.A(_2993_),
    .B(_2995_),
    .X(_2996_));
 sky130_fd_sc_hd__nand2_1 _7827_ (.A(_2993_),
    .B(_2995_),
    .Y(_2997_));
 sky130_fd_sc_hd__nand2_4 _7828_ (.A(_2996_),
    .B(_2997_),
    .Y(_2998_));
 sky130_fd_sc_hd__clkbuf_4 _7829_ (.A(_2998_),
    .X(_2999_));
 sky130_fd_sc_hd__nor3_1 _7830_ (.A(_2984_),
    .B(_2945_),
    .C(_2982_),
    .Y(_3000_));
 sky130_fd_sc_hd__or2_1 _7831_ (.A(_2985_),
    .B(_3000_),
    .X(_3001_));
 sky130_fd_sc_hd__nand2_1 _7832_ (.A(_2995_),
    .B(_3001_),
    .Y(_3003_));
 sky130_fd_sc_hd__nor2_1 _7833_ (.A(_2995_),
    .B(_3001_),
    .Y(_3004_));
 sky130_fd_sc_hd__inv_2 _7834_ (.A(_3004_),
    .Y(_3005_));
 sky130_fd_sc_hd__nand2_2 _7835_ (.A(_3003_),
    .B(_3005_),
    .Y(_3006_));
 sky130_fd_sc_hd__and2_1 _7836_ (.A(_2976_),
    .B(_2978_),
    .X(_3007_));
 sky130_fd_sc_hd__nor2_1 _7837_ (.A(_2979_),
    .B(_3007_),
    .Y(_3008_));
 sky130_fd_sc_hd__xor2_1 _7838_ (.A(_2974_),
    .B(_2975_),
    .X(_3009_));
 sky130_fd_sc_hd__or2_1 _7839_ (.A(_2842_),
    .B(_2973_),
    .X(_3010_));
 sky130_fd_sc_hd__and2_1 _7840_ (.A(_2974_),
    .B(_3010_),
    .X(_3011_));
 sky130_fd_sc_hd__or4_1 _7841_ (.A(_2995_),
    .B(_3008_),
    .C(_3009_),
    .D(_3011_),
    .X(_3012_));
 sky130_fd_sc_hd__or3b_1 _7842_ (.A(_2998_),
    .B(_3006_),
    .C_N(_3012_),
    .X(_3014_));
 sky130_fd_sc_hd__inv_2 _7843_ (.A(_3001_),
    .Y(_3015_));
 sky130_fd_sc_hd__o21ai_1 _7844_ (.A1(_3012_),
    .A2(_3015_),
    .B1(_2993_),
    .Y(_3016_));
 sky130_fd_sc_hd__or3_1 _7845_ (.A(_2986_),
    .B(_2939_),
    .C(_2985_),
    .X(_3017_));
 sky130_fd_sc_hd__and2_1 _7846_ (.A(_2987_),
    .B(_3017_),
    .X(_3018_));
 sky130_fd_sc_hd__xnor2_1 _7847_ (.A(_3016_),
    .B(_3018_),
    .Y(_3019_));
 sky130_fd_sc_hd__xnor2_2 _7848_ (.A(_3014_),
    .B(_3019_),
    .Y(_3020_));
 sky130_fd_sc_hd__clkbuf_4 _7849_ (.A(_3020_),
    .X(_3021_));
 sky130_fd_sc_hd__and3_1 _7850_ (.A(_2988_),
    .B(_2666_),
    .C(_2987_),
    .X(_3022_));
 sky130_fd_sc_hd__or2_2 _7851_ (.A(_2989_),
    .B(_3022_),
    .X(_3023_));
 sky130_fd_sc_hd__clkinv_2 _7852_ (.A(_3020_),
    .Y(_3025_));
 sky130_fd_sc_hd__and2_1 _7853_ (.A(_2993_),
    .B(_2995_),
    .X(_3026_));
 sky130_fd_sc_hd__a21o_1 _7854_ (.A1(_2996_),
    .A2(_3015_),
    .B1(_3026_),
    .X(_3027_));
 sky130_fd_sc_hd__and2_1 _7855_ (.A(_2993_),
    .B(_3020_),
    .X(_3028_));
 sky130_fd_sc_hd__a21o_1 _7856_ (.A1(_3025_),
    .A2(_3027_),
    .B1(_3028_),
    .X(_3029_));
 sky130_fd_sc_hd__xnor2_2 _7857_ (.A(_3023_),
    .B(_3029_),
    .Y(_3030_));
 sky130_fd_sc_hd__or2_1 _7858_ (.A(_3006_),
    .B(_3020_),
    .X(_3031_));
 sky130_fd_sc_hd__o211a_1 _7859_ (.A1(_2999_),
    .A2(_3021_),
    .B1(_3030_),
    .C1(_3031_),
    .X(_3032_));
 sky130_fd_sc_hd__inv_2 _7860_ (.A(_3032_),
    .Y(_3033_));
 sky130_fd_sc_hd__buf_2 _7861_ (.A(_2971_),
    .X(_3034_));
 sky130_fd_sc_hd__or2b_1 _7862_ (.A(_2950_),
    .B_N(_3034_),
    .X(_3036_));
 sky130_fd_sc_hd__o21ai_1 _7863_ (.A1(_2948_),
    .A2(_3034_),
    .B1(_3036_),
    .Y(_3037_));
 sky130_fd_sc_hd__buf_2 _7864_ (.A(_2941_),
    .X(_3038_));
 sky130_fd_sc_hd__mux2_1 _7865_ (.A0(_2928_),
    .A1(_2948_),
    .S(_2971_),
    .X(_3039_));
 sky130_fd_sc_hd__or2_1 _7866_ (.A(_2954_),
    .B(_3039_),
    .X(_3040_));
 sky130_fd_sc_hd__nor2_1 _7867_ (.A(_3038_),
    .B(_3040_),
    .Y(_3041_));
 sky130_fd_sc_hd__clkbuf_4 _7868_ (.A(_2842_),
    .X(_3042_));
 sky130_fd_sc_hd__mux2_1 _7869_ (.A0(_3037_),
    .A1(_3041_),
    .S(_3042_),
    .X(_3043_));
 sky130_fd_sc_hd__buf_2 _7870_ (.A(_2954_),
    .X(_3044_));
 sky130_fd_sc_hd__mux2_1 _7871_ (.A0(_2933_),
    .A1(_2928_),
    .S(_3034_),
    .X(_3045_));
 sky130_fd_sc_hd__or2_1 _7872_ (.A(_3044_),
    .B(_3045_),
    .X(_3047_));
 sky130_fd_sc_hd__nor2_1 _7873_ (.A(_3038_),
    .B(_3047_),
    .Y(_3048_));
 sky130_fd_sc_hd__nor2_1 _7874_ (.A(_3042_),
    .B(_2937_),
    .Y(_3049_));
 sky130_fd_sc_hd__a22o_1 _7875_ (.A1(_3042_),
    .A2(_3048_),
    .B1(_3041_),
    .B2(_3049_),
    .X(_3050_));
 sky130_fd_sc_hd__mux2_1 _7876_ (.A0(_3043_),
    .A1(_3050_),
    .S(_2999_),
    .X(_3051_));
 sky130_fd_sc_hd__mux2_1 _7877_ (.A0(_2923_),
    .A1(_2932_),
    .S(_2971_),
    .X(_3052_));
 sky130_fd_sc_hd__clkinv_2 _7878_ (.A(_3052_),
    .Y(_3053_));
 sky130_fd_sc_hd__mux2_1 _7879_ (.A0(_3053_),
    .A1(_3039_),
    .S(_2954_),
    .X(_3054_));
 sky130_fd_sc_hd__or2_1 _7880_ (.A(_2941_),
    .B(_3054_),
    .X(_3055_));
 sky130_fd_sc_hd__inv_2 _7881_ (.A(_3055_),
    .Y(_3056_));
 sky130_fd_sc_hd__a22o_1 _7882_ (.A1(_3042_),
    .A2(_3056_),
    .B1(_3049_),
    .B2(_3048_),
    .X(_3058_));
 sky130_fd_sc_hd__or2_1 _7883_ (.A(_2937_),
    .B(_2941_),
    .X(_3059_));
 sky130_fd_sc_hd__mux2_1 _7884_ (.A0(_2921_),
    .A1(_2924_),
    .S(_3034_),
    .X(_3060_));
 sky130_fd_sc_hd__mux2_1 _7885_ (.A0(_3060_),
    .A1(_3045_),
    .S(_3044_),
    .X(_3061_));
 sky130_fd_sc_hd__nor2_1 _7886_ (.A(_3059_),
    .B(_3061_),
    .Y(_3062_));
 sky130_fd_sc_hd__a22o_1 _7887_ (.A1(_3042_),
    .A2(_3062_),
    .B1(_3056_),
    .B2(_3049_),
    .X(_3063_));
 sky130_fd_sc_hd__mux2_1 _7888_ (.A0(_3058_),
    .A1(_3063_),
    .S(_2999_),
    .X(_3064_));
 sky130_fd_sc_hd__clkbuf_4 _7889_ (.A(_3006_),
    .X(_3065_));
 sky130_fd_sc_hd__inv_2 _7890_ (.A(_2915_),
    .Y(_3066_));
 sky130_fd_sc_hd__mux2_1 _7891_ (.A0(_3066_),
    .A1(_2921_),
    .S(_2971_),
    .X(_3067_));
 sky130_fd_sc_hd__clkinv_2 _7892_ (.A(_3067_),
    .Y(_3069_));
 sky130_fd_sc_hd__mux2_1 _7893_ (.A0(_3069_),
    .A1(_3052_),
    .S(_2954_),
    .X(_3070_));
 sky130_fd_sc_hd__clkinv_2 _7894_ (.A(_3040_),
    .Y(_3071_));
 sky130_fd_sc_hd__mux2_1 _7895_ (.A0(_3070_),
    .A1(_3071_),
    .S(_3038_),
    .X(_3072_));
 sky130_fd_sc_hd__mux2_1 _7896_ (.A0(_3062_),
    .A1(_3072_),
    .S(_2842_),
    .X(_3073_));
 sky130_fd_sc_hd__clkinv_2 _7897_ (.A(_3073_),
    .Y(_3074_));
 sky130_fd_sc_hd__clkinv_2 _7898_ (.A(_3072_),
    .Y(_3075_));
 sky130_fd_sc_hd__mux2_1 _7899_ (.A0(_2965_),
    .A1(_3066_),
    .S(_2971_),
    .X(_3076_));
 sky130_fd_sc_hd__and2b_1 _7900_ (.A_N(_2954_),
    .B(_3076_),
    .X(_3077_));
 sky130_fd_sc_hd__a21oi_1 _7901_ (.A1(_3044_),
    .A2(_3060_),
    .B1(_3077_),
    .Y(_3078_));
 sky130_fd_sc_hd__clkinv_2 _7902_ (.A(_3078_),
    .Y(_3080_));
 sky130_fd_sc_hd__mux2_1 _7903_ (.A0(_3080_),
    .A1(_3047_),
    .S(_3038_),
    .X(_3081_));
 sky130_fd_sc_hd__mux2_1 _7904_ (.A0(_3075_),
    .A1(_3081_),
    .S(_2842_),
    .X(_3082_));
 sky130_fd_sc_hd__mux2_1 _7905_ (.A0(_3074_),
    .A1(_3082_),
    .S(_2998_),
    .X(_3083_));
 sky130_fd_sc_hd__inv_2 _7906_ (.A(_3083_),
    .Y(_3084_));
 sky130_fd_sc_hd__and2_1 _7907_ (.A(_3065_),
    .B(_3084_),
    .X(_3085_));
 sky130_fd_sc_hd__mux2_1 _7908_ (.A0(_3063_),
    .A1(_3073_),
    .S(_2999_),
    .X(_3086_));
 sky130_fd_sc_hd__mux2_1 _7909_ (.A0(_2908_),
    .A1(_2911_),
    .S(_2971_),
    .X(_3087_));
 sky130_fd_sc_hd__clkinv_2 _7910_ (.A(_3087_),
    .Y(_3088_));
 sky130_fd_sc_hd__mux2_1 _7911_ (.A0(_3088_),
    .A1(_3067_),
    .S(_3044_),
    .X(_3089_));
 sky130_fd_sc_hd__and2b_1 _7912_ (.A_N(_3038_),
    .B(_3089_),
    .X(_3091_));
 sky130_fd_sc_hd__a21oi_1 _7913_ (.A1(_3038_),
    .A2(_3054_),
    .B1(_3091_),
    .Y(_3092_));
 sky130_fd_sc_hd__nand2_1 _7914_ (.A(_3042_),
    .B(_3092_),
    .Y(_3093_));
 sky130_fd_sc_hd__o21ai_1 _7915_ (.A1(_3042_),
    .A2(_3081_),
    .B1(_3093_),
    .Y(_3094_));
 sky130_fd_sc_hd__nand2_1 _7916_ (.A(_2998_),
    .B(_3094_),
    .Y(_3095_));
 sky130_fd_sc_hd__o21a_1 _7917_ (.A1(_2998_),
    .A2(_3082_),
    .B1(_3095_),
    .X(_3096_));
 sky130_fd_sc_hd__inv_2 _7918_ (.A(_3096_),
    .Y(_3097_));
 sky130_fd_sc_hd__and2_1 _7919_ (.A(_3065_),
    .B(_3097_),
    .X(_3098_));
 sky130_fd_sc_hd__o41a_1 _7920_ (.A1(_3064_),
    .A2(_3085_),
    .A3(_3086_),
    .A4(_3098_),
    .B1(_3021_),
    .X(_3099_));
 sky130_fd_sc_hd__mux2_1 _7921_ (.A0(_3050_),
    .A1(_3058_),
    .S(_2999_),
    .X(_3100_));
 sky130_fd_sc_hd__o31a_1 _7922_ (.A1(_3051_),
    .A2(_3099_),
    .A3(_3100_),
    .B1(_3031_),
    .X(_3102_));
 sky130_fd_sc_hd__inv_2 _7923_ (.A(_3031_),
    .Y(_3103_));
 sky130_fd_sc_hd__mux2_1 _7924_ (.A0(_2906_),
    .A1(_2908_),
    .S(_3034_),
    .X(_3104_));
 sky130_fd_sc_hd__a2bb2o_1 _7925_ (.A1_N(_3044_),
    .A2_N(_3104_),
    .B1(_3061_),
    .B2(_3038_),
    .X(_3105_));
 sky130_fd_sc_hd__a21oi_1 _7926_ (.A1(_3044_),
    .A2(_3076_),
    .B1(_3105_),
    .Y(_3106_));
 sky130_fd_sc_hd__mux2_1 _7927_ (.A0(_3092_),
    .A1(_3106_),
    .S(_2842_),
    .X(_3107_));
 sky130_fd_sc_hd__mux2_1 _7928_ (.A0(_3094_),
    .A1(_3107_),
    .S(_2998_),
    .X(_3108_));
 sky130_fd_sc_hd__mux2_1 _7929_ (.A0(_2899_),
    .A1(_2906_),
    .S(_2971_),
    .X(_3109_));
 sky130_fd_sc_hd__mux2_1 _7930_ (.A0(_3109_),
    .A1(_3087_),
    .S(_3044_),
    .X(_3110_));
 sky130_fd_sc_hd__mux2_1 _7931_ (.A0(_3110_),
    .A1(_3070_),
    .S(_3038_),
    .X(_3111_));
 sky130_fd_sc_hd__a21o_1 _7932_ (.A1(_2937_),
    .A2(_3041_),
    .B1(_3111_),
    .X(_3113_));
 sky130_fd_sc_hd__mux2_1 _7933_ (.A0(_3106_),
    .A1(_3113_),
    .S(_2842_),
    .X(_3114_));
 sky130_fd_sc_hd__mux2_1 _7934_ (.A0(_2901_),
    .A1(_2899_),
    .S(_3034_),
    .X(_3115_));
 sky130_fd_sc_hd__mux2_1 _7935_ (.A0(_3115_),
    .A1(_3104_),
    .S(_3044_),
    .X(_3116_));
 sky130_fd_sc_hd__a21o_1 _7936_ (.A1(_3038_),
    .A2(_3078_),
    .B1(_3116_),
    .X(_3117_));
 sky130_fd_sc_hd__mux2_1 _7937_ (.A0(_3117_),
    .A1(_3048_),
    .S(_2937_),
    .X(_3118_));
 sky130_fd_sc_hd__mux2_1 _7938_ (.A0(_3113_),
    .A1(_3118_),
    .S(_2842_),
    .X(_3119_));
 sky130_fd_sc_hd__mux2_1 _7939_ (.A0(_3114_),
    .A1(_3119_),
    .S(_2998_),
    .X(_3120_));
 sky130_fd_sc_hd__mux2_1 _7940_ (.A0(_3108_),
    .A1(_3120_),
    .S(_3006_),
    .X(_3121_));
 sky130_fd_sc_hd__and2_1 _7941_ (.A(_3020_),
    .B(_3121_),
    .X(_3122_));
 sky130_fd_sc_hd__a221o_1 _7942_ (.A1(_3103_),
    .A2(_3064_),
    .B1(_3085_),
    .B2(_3025_),
    .C1(_3122_),
    .X(_3124_));
 sky130_fd_sc_hd__mux2_1 _7943_ (.A0(_3107_),
    .A1(_3114_),
    .S(_2998_),
    .X(_3125_));
 sky130_fd_sc_hd__nor2_1 _7944_ (.A(_2894_),
    .B(_3034_),
    .Y(_3126_));
 sky130_fd_sc_hd__a221o_1 _7945_ (.A1(_2901_),
    .A2(_3034_),
    .B1(_3109_),
    .B2(_3044_),
    .C1(_2941_),
    .X(_3127_));
 sky130_fd_sc_hd__a2bb2o_1 _7946_ (.A1_N(_3126_),
    .A2_N(_3127_),
    .B1(_3038_),
    .B2(_3089_),
    .X(_3128_));
 sky130_fd_sc_hd__a21bo_1 _7947_ (.A1(_2937_),
    .A2(_3056_),
    .B1_N(_3128_),
    .X(_3129_));
 sky130_fd_sc_hd__mux2_1 _7948_ (.A0(_3118_),
    .A1(_3129_),
    .S(_2842_),
    .X(_3130_));
 sky130_fd_sc_hd__mux2_1 _7949_ (.A0(_3119_),
    .A1(_3130_),
    .S(_2998_),
    .X(_3131_));
 sky130_fd_sc_hd__mux2_1 _7950_ (.A0(_3125_),
    .A1(_3131_),
    .S(_3006_),
    .X(_3132_));
 sky130_fd_sc_hd__and2_1 _7951_ (.A(_3020_),
    .B(_3132_),
    .X(_3133_));
 sky130_fd_sc_hd__a221o_1 _7952_ (.A1(_3103_),
    .A2(_3086_),
    .B1(_3098_),
    .B2(_3025_),
    .C1(_3133_),
    .X(_3135_));
 sky130_fd_sc_hd__mux2_1 _7953_ (.A0(_2890_),
    .A1(_2894_),
    .S(_3034_),
    .X(_3136_));
 sky130_fd_sc_hd__inv_2 _7954_ (.A(_3136_),
    .Y(_3137_));
 sky130_fd_sc_hd__a211o_1 _7955_ (.A1(_3044_),
    .A2(_3115_),
    .B1(_3137_),
    .C1(_3059_),
    .X(_3138_));
 sky130_fd_sc_hd__mux2_1 _7956_ (.A0(_3129_),
    .A1(_3138_),
    .S(_3042_),
    .X(_3139_));
 sky130_fd_sc_hd__mux2_1 _7957_ (.A0(_3139_),
    .A1(_3011_),
    .S(_2999_),
    .X(_3140_));
 sky130_fd_sc_hd__mux2_1 _7958_ (.A0(_3009_),
    .A1(_3008_),
    .S(_2999_),
    .X(_3141_));
 sky130_fd_sc_hd__mux2_1 _7959_ (.A0(_3140_),
    .A1(_3141_),
    .S(_3065_),
    .X(_3142_));
 sky130_fd_sc_hd__mux2_1 _7960_ (.A0(_3132_),
    .A1(_3142_),
    .S(_3021_),
    .X(_3143_));
 sky130_fd_sc_hd__mux2_1 _7961_ (.A0(_3084_),
    .A1(_3108_),
    .S(_3006_),
    .X(_3144_));
 sky130_fd_sc_hd__mux2_1 _7962_ (.A0(_3130_),
    .A1(_3139_),
    .S(_2999_),
    .X(_3146_));
 sky130_fd_sc_hd__mux2_1 _7963_ (.A0(_3120_),
    .A1(_3146_),
    .S(_3065_),
    .X(_3147_));
 sky130_fd_sc_hd__mux2_1 _7964_ (.A0(_3144_),
    .A1(_3147_),
    .S(_3021_),
    .X(_3148_));
 sky130_fd_sc_hd__or4_1 _7965_ (.A(_3124_),
    .B(_3135_),
    .C(_3143_),
    .D(_3148_),
    .X(_3149_));
 sky130_fd_sc_hd__mux2_1 _7966_ (.A0(_3011_),
    .A1(_3009_),
    .S(_2999_),
    .X(_3150_));
 sky130_fd_sc_hd__mux2_1 _7967_ (.A0(_3146_),
    .A1(_3150_),
    .S(_3006_),
    .X(_3151_));
 sky130_fd_sc_hd__mux2_1 _7968_ (.A0(_3121_),
    .A1(_3151_),
    .S(_3021_),
    .X(_3152_));
 sky130_fd_sc_hd__mux2_1 _7969_ (.A0(_3051_),
    .A1(_3064_),
    .S(_3065_),
    .X(_3153_));
 sky130_fd_sc_hd__mux2_1 _7970_ (.A0(_3144_),
    .A1(_3153_),
    .S(_3025_),
    .X(_3154_));
 sky130_fd_sc_hd__mux2_1 _7971_ (.A0(_3097_),
    .A1(_3125_),
    .S(_3065_),
    .X(_3155_));
 sky130_fd_sc_hd__mux2_1 _7972_ (.A0(_3131_),
    .A1(_3140_),
    .S(_3065_),
    .X(_3157_));
 sky130_fd_sc_hd__mux2_1 _7973_ (.A0(_3155_),
    .A1(_3157_),
    .S(_3021_),
    .X(_3158_));
 sky130_fd_sc_hd__mux2_1 _7974_ (.A0(_3100_),
    .A1(_3086_),
    .S(_3065_),
    .X(_3159_));
 sky130_fd_sc_hd__mux2_1 _7975_ (.A0(_3155_),
    .A1(_3159_),
    .S(_3025_),
    .X(_3160_));
 sky130_fd_sc_hd__or4_1 _7976_ (.A(_3152_),
    .B(_3154_),
    .C(_3158_),
    .D(_3160_),
    .X(_3161_));
 sky130_fd_sc_hd__o21a_1 _7977_ (.A1(_3149_),
    .A2(_3161_),
    .B1(_3030_),
    .X(_3162_));
 sky130_fd_sc_hd__a21o_1 _7978_ (.A1(_3003_),
    .A2(_3141_),
    .B1(_3004_),
    .X(_3163_));
 sky130_fd_sc_hd__mux2_1 _7979_ (.A0(_3157_),
    .A1(_3163_),
    .S(_3021_),
    .X(_3164_));
 sky130_fd_sc_hd__mux2_1 _7980_ (.A0(_3160_),
    .A1(_3164_),
    .S(_3030_),
    .X(_3165_));
 sky130_fd_sc_hd__buf_2 _7981_ (.A(_2929_),
    .X(_3166_));
 sky130_fd_sc_hd__nor2_1 _7982_ (.A(_3166_),
    .B(_2860_),
    .Y(_3168_));
 sky130_fd_sc_hd__xnor2_1 _7983_ (.A(_2858_),
    .B(_3168_),
    .Y(_3169_));
 sky130_fd_sc_hd__a221o_1 _7984_ (.A1(_3042_),
    .A2(_3037_),
    .B1(_3043_),
    .B2(_2999_),
    .C1(_3169_),
    .X(_3170_));
 sky130_fd_sc_hd__o21ba_1 _7985_ (.A1(_2950_),
    .A2(_3034_),
    .B1_N(_3170_),
    .X(_3171_));
 sky130_fd_sc_hd__or4b_1 _7986_ (.A(_3102_),
    .B(_3162_),
    .C(_3165_),
    .D_N(_3171_),
    .X(_3172_));
 sky130_fd_sc_hd__clkinv_2 _7987_ (.A(_3154_),
    .Y(_3173_));
 sky130_fd_sc_hd__clkinv_2 _7988_ (.A(_3147_),
    .Y(_3174_));
 sky130_fd_sc_hd__clkinv_2 _7989_ (.A(_3150_),
    .Y(_3175_));
 sky130_fd_sc_hd__o21ai_1 _7990_ (.A1(_3026_),
    .A2(_3008_),
    .B1(_2996_),
    .Y(_3176_));
 sky130_fd_sc_hd__mux2_1 _7991_ (.A0(_3175_),
    .A1(_3176_),
    .S(_3065_),
    .X(_3177_));
 sky130_fd_sc_hd__mux2_1 _7992_ (.A0(_3174_),
    .A1(_3177_),
    .S(_3021_),
    .X(_3179_));
 sky130_fd_sc_hd__mux2_1 _7993_ (.A0(_3173_),
    .A1(_3179_),
    .S(_3030_),
    .X(_3180_));
 sky130_fd_sc_hd__a21o_1 _7994_ (.A1(_3033_),
    .A2(_3172_),
    .B1(_3180_),
    .X(_3181_));
 sky130_fd_sc_hd__mux2_4 _7995_ (.A0(_1275_),
    .A1(_1253_),
    .S(_2721_),
    .X(_3182_));
 sky130_fd_sc_hd__xor2_1 _7996_ (.A(_3165_),
    .B(_3180_),
    .X(_3183_));
 sky130_fd_sc_hd__o21ai_1 _7997_ (.A1(_3181_),
    .A2(_3182_),
    .B1(_3183_),
    .Y(_3184_));
 sky130_fd_sc_hd__inv_2 _7998_ (.A(_1253_),
    .Y(_3185_));
 sky130_fd_sc_hd__nand2_1 _7999_ (.A(_1275_),
    .B(_4250_),
    .Y(_3186_));
 sky130_fd_sc_hd__o21a_1 _8000_ (.A1(_3185_),
    .A2(_0121_),
    .B1(_3186_),
    .X(_3187_));
 sky130_fd_sc_hd__o21ai_2 _8001_ (.A1(_3042_),
    .A2(_3138_),
    .B1(_3187_),
    .Y(_3188_));
 sky130_fd_sc_hd__nor3_4 _8002_ (.A(\cmd[7] ),
    .B(\cmd[6] ),
    .C(_3188_),
    .Y(_3190_));
 sky130_fd_sc_hd__o31a_1 _8003_ (.A1(_3165_),
    .A2(_3181_),
    .A3(_3182_),
    .B1(_3190_),
    .X(_3191_));
 sky130_fd_sc_hd__nand2_1 _8004_ (.A(_3184_),
    .B(_3191_),
    .Y(_3192_));
 sky130_fd_sc_hd__o31a_1 _8005_ (.A1(_2619_),
    .A2(_2621_),
    .A3(_2622_),
    .B1(_3192_),
    .X(_3193_));
 sky130_fd_sc_hd__o31a_1 _8006_ (.A1(_0598_),
    .A2(_0600_),
    .A3(_0602_),
    .B1(_3193_),
    .X(_3194_));
 sky130_fd_sc_hd__clkbuf_4 _8007_ (.A(_1177_),
    .X(_3195_));
 sky130_fd_sc_hd__o2bb2a_1 _8008_ (.A1_N(\out_reg[0] ),
    .A2_N(_1231_),
    .B1(_3194_),
    .B2(_3195_),
    .X(_3196_));
 sky130_fd_sc_hd__nor2_1 _8009_ (.A(_1220_),
    .B(_3196_),
    .Y(_0020_));
 sky130_fd_sc_hd__buf_2 _8010_ (.A(_1231_),
    .X(_3197_));
 sky130_fd_sc_hd__o211a_1 _8011_ (.A1(_2611_),
    .A2(_2615_),
    .B1(_2616_),
    .C1(_2609_),
    .X(_3198_));
 sky130_fd_sc_hd__nand2_2 _8012_ (.A(_2521_),
    .B(_3198_),
    .Y(_3200_));
 sky130_fd_sc_hd__or2_1 _8013_ (.A(_2521_),
    .B(_2618_),
    .X(_3201_));
 sky130_fd_sc_hd__and3_1 _8014_ (.A(_1319_),
    .B(_3200_),
    .C(_3201_),
    .X(_3202_));
 sky130_fd_sc_hd__a21o_1 _8015_ (.A1(_2451_),
    .A2(_2578_),
    .B1(_2590_),
    .X(_3203_));
 sky130_fd_sc_hd__nand2_1 _8016_ (.A(_2392_),
    .B(_2494_),
    .Y(_3204_));
 sky130_fd_sc_hd__o211a_1 _8017_ (.A1(_2494_),
    .A2(_2613_),
    .B1(_3204_),
    .C1(_2486_),
    .X(_3205_));
 sky130_fd_sc_hd__a211o_1 _8018_ (.A1(_2514_),
    .A2(_3203_),
    .B1(_3205_),
    .C1(_2611_),
    .X(_3206_));
 sky130_fd_sc_hd__a21boi_2 _8019_ (.A1(_2611_),
    .A2(_2588_),
    .B1_N(_3206_),
    .Y(_3207_));
 sky130_fd_sc_hd__xnor2_1 _8020_ (.A(_3200_),
    .B(_3207_),
    .Y(_3208_));
 sky130_fd_sc_hd__nand2_1 _8021_ (.A(_3202_),
    .B(_3207_),
    .Y(_3209_));
 sky130_fd_sc_hd__and3b_1 _8022_ (.A_N(\cmd[6] ),
    .B(_2319_),
    .C(\cmd[7] ),
    .X(_3211_));
 sky130_fd_sc_hd__buf_2 _8023_ (.A(_3211_),
    .X(_3212_));
 sky130_fd_sc_hd__o211a_1 _8024_ (.A1(_3202_),
    .A2(_3208_),
    .B1(_3209_),
    .C1(_3212_),
    .X(_3213_));
 sky130_fd_sc_hd__or2_1 _8025_ (.A(_0594_),
    .B(_0597_),
    .X(_3214_));
 sky130_fd_sc_hd__mux2_1 _8026_ (.A0(_0451_),
    .A1(_0512_),
    .S(_0515_),
    .X(_3215_));
 sky130_fd_sc_hd__nand2_1 _8027_ (.A(_0557_),
    .B(_3215_),
    .Y(_3216_));
 sky130_fd_sc_hd__o21ai_2 _8028_ (.A1(_0557_),
    .A2(_0569_),
    .B1(_3216_),
    .Y(_3217_));
 sky130_fd_sc_hd__clkinv_2 _8029_ (.A(_3217_),
    .Y(_3218_));
 sky130_fd_sc_hd__mux2_1 _8030_ (.A0(_0583_),
    .A1(_3218_),
    .S(_0519_),
    .X(_3219_));
 sky130_fd_sc_hd__xnor2_1 _8031_ (.A(_0595_),
    .B(_3219_),
    .Y(_3220_));
 sky130_fd_sc_hd__and3_1 _8032_ (.A(_0601_),
    .B(_3214_),
    .C(_3220_),
    .X(_3222_));
 sky130_fd_sc_hd__a21oi_1 _8033_ (.A1(_1330_),
    .A2(_3214_),
    .B1(_3220_),
    .Y(_3223_));
 sky130_fd_sc_hd__nor3_2 _8034_ (.A(_0600_),
    .B(_3222_),
    .C(_3223_),
    .Y(_3224_));
 sky130_fd_sc_hd__inv_2 _8035_ (.A(_1275_),
    .Y(_3225_));
 sky130_fd_sc_hd__mux2_1 _8036_ (.A0(_3225_),
    .A1(_3185_),
    .S(_2721_),
    .X(_3226_));
 sky130_fd_sc_hd__buf_2 _8037_ (.A(_3226_),
    .X(_3227_));
 sky130_fd_sc_hd__and2_1 _8038_ (.A(_3181_),
    .B(_3183_),
    .X(_3228_));
 sky130_fd_sc_hd__and3b_1 _8039_ (.A_N(_3180_),
    .B(_3033_),
    .C(_3165_),
    .X(_3229_));
 sky130_fd_sc_hd__mux2_1 _8040_ (.A0(_3176_),
    .A1(_2993_),
    .S(_3065_),
    .X(_3230_));
 sky130_fd_sc_hd__clkinv_2 _8041_ (.A(_3230_),
    .Y(_3231_));
 sky130_fd_sc_hd__mux2_1 _8042_ (.A0(_3151_),
    .A1(_3231_),
    .S(_3021_),
    .X(_3233_));
 sky130_fd_sc_hd__buf_2 _8043_ (.A(_3030_),
    .X(_3234_));
 sky130_fd_sc_hd__mux2_1 _8044_ (.A0(_3124_),
    .A1(_3233_),
    .S(_3234_),
    .X(_3235_));
 sky130_fd_sc_hd__nand2_1 _8045_ (.A(_3229_),
    .B(_3235_),
    .Y(_3236_));
 sky130_fd_sc_hd__or2_1 _8046_ (.A(_3229_),
    .B(_3235_),
    .X(_3237_));
 sky130_fd_sc_hd__nand2_1 _8047_ (.A(_3236_),
    .B(_3237_),
    .Y(_3238_));
 sky130_fd_sc_hd__or3_1 _8048_ (.A(_3227_),
    .B(_3228_),
    .C(_3238_),
    .X(_3239_));
 sky130_fd_sc_hd__o21ai_1 _8049_ (.A1(_3227_),
    .A2(_3228_),
    .B1(_3238_),
    .Y(_3240_));
 sky130_fd_sc_hd__a31o_1 _8050_ (.A1(_3190_),
    .A2(_3239_),
    .A3(_3240_),
    .B1(_0701_),
    .X(_3241_));
 sky130_fd_sc_hd__buf_2 _8051_ (.A(_0786_),
    .X(_3242_));
 sky130_fd_sc_hd__a21bo_1 _8052_ (.A1(\out_reg[0] ),
    .A2(_3242_),
    .B1_N(_0701_),
    .X(_3244_));
 sky130_fd_sc_hd__o31a_1 _8053_ (.A1(_3213_),
    .A2(_3224_),
    .A3(_3241_),
    .B1(_3244_),
    .X(_3245_));
 sky130_fd_sc_hd__a21oi_1 _8054_ (.A1(\out_reg[1] ),
    .A2(_3197_),
    .B1(_3245_),
    .Y(_3246_));
 sky130_fd_sc_hd__nor2_1 _8055_ (.A(_1220_),
    .B(_3246_),
    .Y(_0021_));
 sky130_fd_sc_hd__a21o_1 _8056_ (.A1(_3200_),
    .A2(_3201_),
    .B1(_3208_),
    .X(_3247_));
 sky130_fd_sc_hd__and2_1 _8057_ (.A(_1319_),
    .B(_3247_),
    .X(_3248_));
 sky130_fd_sc_hd__nand3_2 _8058_ (.A(_2521_),
    .B(_3198_),
    .C(_3207_),
    .Y(_3249_));
 sky130_fd_sc_hd__o21ai_1 _8059_ (.A1(_2348_),
    .A2(_2522_),
    .B1(_3204_),
    .Y(_3250_));
 sky130_fd_sc_hd__mux2_1 _8060_ (.A0(_2597_),
    .A1(_3250_),
    .S(_2486_),
    .X(_3251_));
 sky130_fd_sc_hd__mux2_2 _8061_ (.A0(_2602_),
    .A1(_3251_),
    .S(_2520_),
    .X(_3252_));
 sky130_fd_sc_hd__xor2_4 _8062_ (.A(_3249_),
    .B(_3252_),
    .X(_3254_));
 sky130_fd_sc_hd__o21ai_1 _8063_ (.A1(_3248_),
    .A2(_3254_),
    .B1(_3212_),
    .Y(_3255_));
 sky130_fd_sc_hd__a21oi_2 _8064_ (.A1(_3248_),
    .A2(_3254_),
    .B1(_3255_),
    .Y(_3256_));
 sky130_fd_sc_hd__nor2_1 _8065_ (.A(_3214_),
    .B(_3220_),
    .Y(_3257_));
 sky130_fd_sc_hd__or2b_1 _8066_ (.A(_0595_),
    .B_N(_3219_),
    .X(_3258_));
 sky130_fd_sc_hd__clkbuf_4 _8067_ (.A(_0519_),
    .X(_3259_));
 sky130_fd_sc_hd__mux2_1 _8068_ (.A0(_0440_),
    .A1(_0398_),
    .S(_0515_),
    .X(_3260_));
 sky130_fd_sc_hd__mux2_1 _8069_ (.A0(_0572_),
    .A1(_3260_),
    .S(_0557_),
    .X(_3261_));
 sky130_fd_sc_hd__or2_1 _8070_ (.A(_0521_),
    .B(_3261_),
    .X(_3262_));
 sky130_fd_sc_hd__o21ai_1 _8071_ (.A1(_3259_),
    .A2(_0585_),
    .B1(_3262_),
    .Y(_3263_));
 sky130_fd_sc_hd__nor2_2 _8072_ (.A(_3258_),
    .B(_3263_),
    .Y(_3265_));
 sky130_fd_sc_hd__and2_1 _8073_ (.A(_3258_),
    .B(_3263_),
    .X(_3266_));
 sky130_fd_sc_hd__or2_1 _8074_ (.A(_3265_),
    .B(_3266_),
    .X(_3267_));
 sky130_fd_sc_hd__o21a_1 _8075_ (.A1(_3166_),
    .A2(_3257_),
    .B1(_3267_),
    .X(_3268_));
 sky130_fd_sc_hd__nor2_1 _8076_ (.A(_0600_),
    .B(_3268_),
    .Y(_3269_));
 sky130_fd_sc_hd__o31a_1 _8077_ (.A1(_3166_),
    .A2(_3257_),
    .A3(_3267_),
    .B1(_3269_),
    .X(_3270_));
 sky130_fd_sc_hd__and2_1 _8078_ (.A(_3228_),
    .B(_3238_),
    .X(_3271_));
 sky130_fd_sc_hd__clkinv_2 _8079_ (.A(_3142_),
    .Y(_3272_));
 sky130_fd_sc_hd__mux2_1 _8080_ (.A0(_3027_),
    .A1(_3272_),
    .S(_3025_),
    .X(_3273_));
 sky130_fd_sc_hd__clkinv_2 _8081_ (.A(_3273_),
    .Y(_3274_));
 sky130_fd_sc_hd__mux2_1 _8082_ (.A0(_3135_),
    .A1(_3274_),
    .S(_3030_),
    .X(_3276_));
 sky130_fd_sc_hd__xor2_1 _8083_ (.A(_3236_),
    .B(_3276_),
    .X(_3277_));
 sky130_fd_sc_hd__o21ai_1 _8084_ (.A1(_3227_),
    .A2(_3271_),
    .B1(_3277_),
    .Y(_3278_));
 sky130_fd_sc_hd__or3_1 _8085_ (.A(_3227_),
    .B(_3271_),
    .C(_3277_),
    .X(_3279_));
 sky130_fd_sc_hd__a31o_1 _8086_ (.A1(_3190_),
    .A2(_3278_),
    .A3(_3279_),
    .B1(_0701_),
    .X(_3280_));
 sky130_fd_sc_hd__a21bo_1 _8087_ (.A1(\out_reg[1] ),
    .A2(_3242_),
    .B1_N(_0701_),
    .X(_3281_));
 sky130_fd_sc_hd__o31a_1 _8088_ (.A1(_3256_),
    .A2(_3270_),
    .A3(_3280_),
    .B1(_3281_),
    .X(_3282_));
 sky130_fd_sc_hd__a21oi_1 _8089_ (.A1(\out_reg[2] ),
    .A2(_3197_),
    .B1(_3282_),
    .Y(_3283_));
 sky130_fd_sc_hd__nor2_1 _8090_ (.A(_1220_),
    .B(_3283_),
    .Y(_0022_));
 sky130_fd_sc_hd__and4b_2 _8091_ (.A_N(_3252_),
    .B(_3207_),
    .C(_3198_),
    .D(_2521_),
    .X(_3284_));
 sky130_fd_sc_hd__nand2_2 _8092_ (.A(_2392_),
    .B(_2486_),
    .Y(_3286_));
 sky130_fd_sc_hd__o21a_1 _8093_ (.A1(_2486_),
    .A2(_2614_),
    .B1(_3286_),
    .X(_3287_));
 sky130_fd_sc_hd__clkinv_2 _8094_ (.A(_3287_),
    .Y(_3288_));
 sky130_fd_sc_hd__mux2_2 _8095_ (.A0(_2585_),
    .A1(_3288_),
    .S(_2604_),
    .X(_3289_));
 sky130_fd_sc_hd__xnor2_2 _8096_ (.A(_3284_),
    .B(_3289_),
    .Y(_3290_));
 sky130_fd_sc_hd__o21a_1 _8097_ (.A1(_3247_),
    .A2(_3254_),
    .B1(_0601_),
    .X(_3291_));
 sky130_fd_sc_hd__a21oi_1 _8098_ (.A1(_3290_),
    .A2(_3291_),
    .B1(_2621_),
    .Y(_3292_));
 sky130_fd_sc_hd__o21ai_1 _8099_ (.A1(_3290_),
    .A2(_3291_),
    .B1(_3292_),
    .Y(_3293_));
 sky130_fd_sc_hd__and3_1 _8100_ (.A(_3228_),
    .B(_3238_),
    .C(_3277_),
    .X(_3294_));
 sky130_fd_sc_hd__or2_1 _8101_ (.A(_3227_),
    .B(_3294_),
    .X(_3295_));
 sky130_fd_sc_hd__and3_1 _8102_ (.A(_3229_),
    .B(_3235_),
    .C(_3276_),
    .X(_3297_));
 sky130_fd_sc_hd__a21o_1 _8103_ (.A1(_3025_),
    .A2(_3177_),
    .B1(_3028_),
    .X(_3298_));
 sky130_fd_sc_hd__clkinv_2 _8104_ (.A(_3298_),
    .Y(_3299_));
 sky130_fd_sc_hd__mux2_1 _8105_ (.A0(_3148_),
    .A1(_3299_),
    .S(_3234_),
    .X(_3300_));
 sky130_fd_sc_hd__xnor2_1 _8106_ (.A(_3297_),
    .B(_3300_),
    .Y(_3301_));
 sky130_fd_sc_hd__nor2_1 _8107_ (.A(_3295_),
    .B(_3301_),
    .Y(_3302_));
 sky130_fd_sc_hd__or3_2 _8108_ (.A(\cmd[7] ),
    .B(\cmd[6] ),
    .C(_3188_),
    .X(_3303_));
 sky130_fd_sc_hd__a211o_1 _8109_ (.A1(_3295_),
    .A2(_3301_),
    .B1(_3302_),
    .C1(_3303_),
    .X(_3304_));
 sky130_fd_sc_hd__nand2_1 _8110_ (.A(_3257_),
    .B(_3267_),
    .Y(_3305_));
 sky130_fd_sc_hd__nand2_1 _8111_ (.A(_0451_),
    .B(_0557_),
    .Y(_3306_));
 sky130_fd_sc_hd__a21boi_1 _8112_ (.A1(_0535_),
    .A2(_0516_),
    .B1_N(_3306_),
    .Y(_3308_));
 sky130_fd_sc_hd__mux2_1 _8113_ (.A0(_0586_),
    .A1(_3308_),
    .S(_3259_),
    .X(_3309_));
 sky130_fd_sc_hd__xor2_2 _8114_ (.A(_3265_),
    .B(_3309_),
    .X(_3310_));
 sky130_fd_sc_hd__a21oi_1 _8115_ (.A1(_1330_),
    .A2(_3305_),
    .B1(_3310_),
    .Y(_3311_));
 sky130_fd_sc_hd__a31o_1 _8116_ (.A1(_0601_),
    .A2(_3305_),
    .A3(_3310_),
    .B1(_0600_),
    .X(_3312_));
 sky130_fd_sc_hd__or2_1 _8117_ (.A(_3311_),
    .B(_3312_),
    .X(_3313_));
 sky130_fd_sc_hd__a31o_1 _8118_ (.A1(_3293_),
    .A2(_3304_),
    .A3(_3313_),
    .B1(_3195_),
    .X(_3314_));
 sky130_fd_sc_hd__and2_1 _8119_ (.A(_0701_),
    .B(_0786_),
    .X(_3315_));
 sky130_fd_sc_hd__clkbuf_2 _8120_ (.A(_3315_),
    .X(_3316_));
 sky130_fd_sc_hd__a22oi_1 _8121_ (.A1(\out_reg[2] ),
    .A2(_3316_),
    .B1(_3197_),
    .B2(\out_reg[3] ),
    .Y(_3317_));
 sky130_fd_sc_hd__a21oi_1 _8122_ (.A1(_3314_),
    .A2(_3317_),
    .B1(_0635_),
    .Y(_0023_));
 sky130_fd_sc_hd__or3_2 _8123_ (.A(_3249_),
    .B(_3252_),
    .C(_3289_),
    .X(_3319_));
 sky130_fd_sc_hd__o211a_1 _8124_ (.A1(_2569_),
    .A2(_2495_),
    .B1(_3286_),
    .C1(_2520_),
    .X(_3320_));
 sky130_fd_sc_hd__a21oi_4 _8125_ (.A1(_2611_),
    .A2(_2576_),
    .B1(_3320_),
    .Y(_3321_));
 sky130_fd_sc_hd__xor2_4 _8126_ (.A(_3319_),
    .B(_3321_),
    .X(_3322_));
 sky130_fd_sc_hd__a2111oi_2 _8127_ (.A1(_3200_),
    .A2(_3201_),
    .B1(_3208_),
    .C1(_3254_),
    .D1(_3290_),
    .Y(_3323_));
 sky130_fd_sc_hd__or2_1 _8128_ (.A(_3166_),
    .B(_3323_),
    .X(_3324_));
 sky130_fd_sc_hd__xnor2_2 _8129_ (.A(_3322_),
    .B(_3324_),
    .Y(_3325_));
 sky130_fd_sc_hd__o21ba_1 _8130_ (.A1(_3021_),
    .A2(_3163_),
    .B1_N(_3028_),
    .X(_3326_));
 sky130_fd_sc_hd__mux2_1 _8131_ (.A0(_3158_),
    .A1(_3326_),
    .S(_3234_),
    .X(_3327_));
 sky130_fd_sc_hd__nand3_1 _8132_ (.A(_3297_),
    .B(_3300_),
    .C(_3327_),
    .Y(_3329_));
 sky130_fd_sc_hd__a21o_1 _8133_ (.A1(_3297_),
    .A2(_3300_),
    .B1(_3327_),
    .X(_3330_));
 sky130_fd_sc_hd__and2_1 _8134_ (.A(_3329_),
    .B(_3330_),
    .X(_3331_));
 sky130_fd_sc_hd__a21oi_1 _8135_ (.A1(_3294_),
    .A2(_3301_),
    .B1(_3226_),
    .Y(_3332_));
 sky130_fd_sc_hd__nand2_1 _8136_ (.A(_3331_),
    .B(_3332_),
    .Y(_3333_));
 sky130_fd_sc_hd__or2_1 _8137_ (.A(_3331_),
    .B(_3332_),
    .X(_3334_));
 sky130_fd_sc_hd__and3_1 _8138_ (.A(_3190_),
    .B(_3333_),
    .C(_3334_),
    .X(_3335_));
 sky130_fd_sc_hd__nor2_1 _8139_ (.A(_3305_),
    .B(_3310_),
    .Y(_3336_));
 sky130_fd_sc_hd__o21a_1 _8140_ (.A1(_0557_),
    .A2(_0527_),
    .B1(_3306_),
    .X(_3337_));
 sky130_fd_sc_hd__mux2_1 _8141_ (.A0(_0584_),
    .A1(_3337_),
    .S(_3259_),
    .X(_3338_));
 sky130_fd_sc_hd__nand3_1 _8142_ (.A(_3265_),
    .B(_3309_),
    .C(_3338_),
    .Y(_3340_));
 sky130_fd_sc_hd__a21o_1 _8143_ (.A1(_3265_),
    .A2(_3309_),
    .B1(_3338_),
    .X(_3341_));
 sky130_fd_sc_hd__nand2_1 _8144_ (.A(_3340_),
    .B(_3341_),
    .Y(_3342_));
 sky130_fd_sc_hd__o21a_1 _8145_ (.A1(_3166_),
    .A2(_3336_),
    .B1(_3342_),
    .X(_3343_));
 sky130_fd_sc_hd__nor2_1 _8146_ (.A(_0599_),
    .B(_3343_),
    .Y(_3344_));
 sky130_fd_sc_hd__o31a_1 _8147_ (.A1(_3166_),
    .A2(_3336_),
    .A3(_3342_),
    .B1(_3344_),
    .X(_3345_));
 sky130_fd_sc_hd__a2111oi_4 _8148_ (.A1(_3212_),
    .A2(_3325_),
    .B1(_3335_),
    .C1(_3345_),
    .D1(_1177_),
    .Y(_3346_));
 sky130_fd_sc_hd__a21boi_1 _8149_ (.A1(\out_reg[3] ),
    .A2(_3242_),
    .B1_N(_1177_),
    .Y(_3347_));
 sky130_fd_sc_hd__o2bb2a_1 _8150_ (.A1_N(\out_reg[4] ),
    .A2_N(_1231_),
    .B1(_3346_),
    .B2(_3347_),
    .X(_3348_));
 sky130_fd_sc_hd__nor2_1 _8151_ (.A(_1220_),
    .B(_3348_),
    .Y(_0024_));
 sky130_fd_sc_hd__or2b_1 _8152_ (.A(_3322_),
    .B_N(_3323_),
    .X(_3350_));
 sky130_fd_sc_hd__or3b_1 _8153_ (.A(_3289_),
    .B(_3321_),
    .C_N(_3284_),
    .X(_3351_));
 sky130_fd_sc_hd__o21a_1 _8154_ (.A1(_2522_),
    .A2(_2613_),
    .B1(_3204_),
    .X(_3352_));
 sky130_fd_sc_hd__o211ai_1 _8155_ (.A1(_2569_),
    .A2(_3352_),
    .B1(_3286_),
    .C1(_2520_),
    .Y(_3353_));
 sky130_fd_sc_hd__o21ai_2 _8156_ (.A1(_2604_),
    .A2(_2592_),
    .B1(_3353_),
    .Y(_3354_));
 sky130_fd_sc_hd__xnor2_2 _8157_ (.A(_3351_),
    .B(_3354_),
    .Y(_3355_));
 sky130_fd_sc_hd__a21oi_1 _8158_ (.A1(_1330_),
    .A2(_3350_),
    .B1(_3355_),
    .Y(_3356_));
 sky130_fd_sc_hd__a31o_1 _8159_ (.A1(_0601_),
    .A2(_3350_),
    .A3(_3355_),
    .B1(_2621_),
    .X(_3357_));
 sky130_fd_sc_hd__or2_1 _8160_ (.A(_3356_),
    .B(_3357_),
    .X(_3358_));
 sky130_fd_sc_hd__nand2_1 _8161_ (.A(_3336_),
    .B(_3342_),
    .Y(_3359_));
 sky130_fd_sc_hd__clkinv_2 _8162_ (.A(_0570_),
    .Y(_3361_));
 sky130_fd_sc_hd__a21boi_1 _8163_ (.A1(_0535_),
    .A2(_3215_),
    .B1_N(_3306_),
    .Y(_3362_));
 sky130_fd_sc_hd__inv_2 _8164_ (.A(_3362_),
    .Y(_3363_));
 sky130_fd_sc_hd__mux2_1 _8165_ (.A0(_3361_),
    .A1(_3363_),
    .S(_3259_),
    .X(_3364_));
 sky130_fd_sc_hd__nor2_1 _8166_ (.A(_3340_),
    .B(_3364_),
    .Y(_3365_));
 sky130_fd_sc_hd__and2_1 _8167_ (.A(_3340_),
    .B(_3364_),
    .X(_3366_));
 sky130_fd_sc_hd__nor2_1 _8168_ (.A(_3365_),
    .B(_3366_),
    .Y(_3367_));
 sky130_fd_sc_hd__a21oi_1 _8169_ (.A1(_1330_),
    .A2(_3359_),
    .B1(_3367_),
    .Y(_3368_));
 sky130_fd_sc_hd__a311o_1 _8170_ (.A1(_1330_),
    .A2(_3359_),
    .A3(_3367_),
    .B1(_3368_),
    .C1(_0600_),
    .X(_3369_));
 sky130_fd_sc_hd__a21o_1 _8171_ (.A1(_3025_),
    .A2(_3230_),
    .B1(_3028_),
    .X(_3370_));
 sky130_fd_sc_hd__clkinv_2 _8172_ (.A(_3370_),
    .Y(_3372_));
 sky130_fd_sc_hd__mux2_1 _8173_ (.A0(_3152_),
    .A1(_3372_),
    .S(_3234_),
    .X(_3373_));
 sky130_fd_sc_hd__xnor2_1 _8174_ (.A(_3329_),
    .B(_3373_),
    .Y(_3374_));
 sky130_fd_sc_hd__and2_1 _8175_ (.A(_3182_),
    .B(_3334_),
    .X(_3375_));
 sky130_fd_sc_hd__o21ai_1 _8176_ (.A1(_3374_),
    .A2(_3375_),
    .B1(_3190_),
    .Y(_3376_));
 sky130_fd_sc_hd__a21o_1 _8177_ (.A1(_3374_),
    .A2(_3375_),
    .B1(_3376_),
    .X(_3377_));
 sky130_fd_sc_hd__a31o_2 _8178_ (.A1(_3358_),
    .A2(_3369_),
    .A3(_3377_),
    .B1(_3195_),
    .X(_3378_));
 sky130_fd_sc_hd__a22oi_1 _8179_ (.A1(\out_reg[4] ),
    .A2(_3316_),
    .B1(_3197_),
    .B2(\out_reg[5] ),
    .Y(_3379_));
 sky130_fd_sc_hd__a21oi_1 _8180_ (.A1(_3378_),
    .A2(_3379_),
    .B1(_0635_),
    .Y(_0025_));
 sky130_fd_sc_hd__or2_1 _8181_ (.A(_3359_),
    .B(_3367_),
    .X(_3380_));
 sky130_fd_sc_hd__nand2_1 _8182_ (.A(_0601_),
    .B(_3380_),
    .Y(_3382_));
 sky130_fd_sc_hd__clkinv_2 _8183_ (.A(_0573_),
    .Y(_3383_));
 sky130_fd_sc_hd__o21ai_1 _8184_ (.A1(_0557_),
    .A2(_3260_),
    .B1(_3306_),
    .Y(_3384_));
 sky130_fd_sc_hd__mux2_1 _8185_ (.A0(_3383_),
    .A1(_3384_),
    .S(_3259_),
    .X(_3385_));
 sky130_fd_sc_hd__xnor2_1 _8186_ (.A(_3365_),
    .B(_3385_),
    .Y(_3386_));
 sky130_fd_sc_hd__xor2_1 _8187_ (.A(_3382_),
    .B(_3386_),
    .X(_3387_));
 sky130_fd_sc_hd__and2b_1 _8188_ (.A_N(_3329_),
    .B(_3373_),
    .X(_3388_));
 sky130_fd_sc_hd__nand2_1 _8189_ (.A(_3023_),
    .B(_3029_),
    .Y(_3389_));
 sky130_fd_sc_hd__o21a_1 _8190_ (.A1(_3234_),
    .A2(_3143_),
    .B1(_3389_),
    .X(_3390_));
 sky130_fd_sc_hd__and2_1 _8191_ (.A(_3388_),
    .B(_3390_),
    .X(_3391_));
 sky130_fd_sc_hd__nor2_1 _8192_ (.A(_3388_),
    .B(_3390_),
    .Y(_3393_));
 sky130_fd_sc_hd__nor2_1 _8193_ (.A(_3391_),
    .B(_3393_),
    .Y(_3394_));
 sky130_fd_sc_hd__o21a_1 _8194_ (.A1(_3334_),
    .A2(_3374_),
    .B1(_3182_),
    .X(_3395_));
 sky130_fd_sc_hd__or2_1 _8195_ (.A(_3394_),
    .B(_3395_),
    .X(_3396_));
 sky130_fd_sc_hd__a21oi_1 _8196_ (.A1(_3394_),
    .A2(_3395_),
    .B1(_3303_),
    .Y(_3397_));
 sky130_fd_sc_hd__nand2_1 _8197_ (.A(_3396_),
    .B(_3397_),
    .Y(_3398_));
 sky130_fd_sc_hd__or3b_1 _8198_ (.A(_3322_),
    .B(_3355_),
    .C_N(_3323_),
    .X(_3399_));
 sky130_fd_sc_hd__nand2_1 _8199_ (.A(_0601_),
    .B(_3399_),
    .Y(_3400_));
 sky130_fd_sc_hd__or2b_1 _8200_ (.A(_3321_),
    .B_N(_3354_),
    .X(_3401_));
 sky130_fd_sc_hd__or3b_1 _8201_ (.A(_3289_),
    .B(_3401_),
    .C_N(_3284_),
    .X(_3402_));
 sky130_fd_sc_hd__a21bo_1 _8202_ (.A1(_2514_),
    .A2(_3250_),
    .B1_N(_3286_),
    .X(_3404_));
 sky130_fd_sc_hd__mux2_1 _8203_ (.A0(_2598_),
    .A1(_3404_),
    .S(_2520_),
    .X(_3405_));
 sky130_fd_sc_hd__nor3b_1 _8204_ (.A(_3321_),
    .B(_3405_),
    .C_N(_3354_),
    .Y(_3406_));
 sky130_fd_sc_hd__and3b_1 _8205_ (.A_N(_3289_),
    .B(_3406_),
    .C(_3284_),
    .X(_3407_));
 sky130_fd_sc_hd__a21o_1 _8206_ (.A1(_3402_),
    .A2(_3405_),
    .B1(_3407_),
    .X(_3408_));
 sky130_fd_sc_hd__a21oi_1 _8207_ (.A1(_3400_),
    .A2(_3408_),
    .B1(_2621_),
    .Y(_3409_));
 sky130_fd_sc_hd__o21ai_1 _8208_ (.A1(_3400_),
    .A2(_3408_),
    .B1(_3409_),
    .Y(_3410_));
 sky130_fd_sc_hd__o211a_1 _8209_ (.A1(_0600_),
    .A2(_3387_),
    .B1(_3398_),
    .C1(_3410_),
    .X(_3411_));
 sky130_fd_sc_hd__a22o_1 _8210_ (.A1(\out_reg[5] ),
    .A2(_3316_),
    .B1(_1231_),
    .B2(\out_reg[6] ),
    .X(_3412_));
 sky130_fd_sc_hd__o21ba_1 _8211_ (.A1(_3195_),
    .A2(_3411_),
    .B1_N(_3412_),
    .X(_3413_));
 sky130_fd_sc_hd__nor2_1 _8212_ (.A(_1220_),
    .B(_3413_),
    .Y(_0026_));
 sky130_fd_sc_hd__or4bb_1 _8213_ (.A(_3322_),
    .B(_3355_),
    .C_N(_3408_),
    .D_N(_3323_),
    .X(_3415_));
 sky130_fd_sc_hd__nor2_4 _8214_ (.A(_2491_),
    .B(_2611_),
    .Y(_3416_));
 sky130_fd_sc_hd__o21ba_1 _8215_ (.A1(_2604_),
    .A2(_2615_),
    .B1_N(_3416_),
    .X(_3417_));
 sky130_fd_sc_hd__and4b_1 _8216_ (.A_N(_3289_),
    .B(_3406_),
    .C(_3417_),
    .D(_3284_),
    .X(_3418_));
 sky130_fd_sc_hd__buf_2 _8217_ (.A(_3418_),
    .X(_3419_));
 sky130_fd_sc_hd__nor2_1 _8218_ (.A(_3407_),
    .B(_3417_),
    .Y(_3420_));
 sky130_fd_sc_hd__nor2_1 _8219_ (.A(_3419_),
    .B(_3420_),
    .Y(_3421_));
 sky130_fd_sc_hd__a21oi_1 _8220_ (.A1(_1330_),
    .A2(_3415_),
    .B1(_3421_),
    .Y(_3422_));
 sky130_fd_sc_hd__a31o_1 _8221_ (.A1(_0601_),
    .A2(_3421_),
    .A3(_3415_),
    .B1(_2621_),
    .X(_3423_));
 sky130_fd_sc_hd__or2_1 _8222_ (.A(_3422_),
    .B(_3423_),
    .X(_3425_));
 sky130_fd_sc_hd__nor2_1 _8223_ (.A(_3380_),
    .B(_3386_),
    .Y(_3426_));
 sky130_fd_sc_hd__or2_1 _8224_ (.A(_3166_),
    .B(_3426_),
    .X(_3427_));
 sky130_fd_sc_hd__or3_1 _8225_ (.A(_3340_),
    .B(_3364_),
    .C(_3385_),
    .X(_3428_));
 sky130_fd_sc_hd__nor2_2 _8226_ (.A(_0440_),
    .B(_0521_),
    .Y(_3429_));
 sky130_fd_sc_hd__a21o_1 _8227_ (.A1(_0521_),
    .A2(_0517_),
    .B1(_3429_),
    .X(_3430_));
 sky130_fd_sc_hd__or2_1 _8228_ (.A(_3428_),
    .B(_3430_),
    .X(_3431_));
 sky130_fd_sc_hd__nand2_1 _8229_ (.A(_3428_),
    .B(_3430_),
    .Y(_3432_));
 sky130_fd_sc_hd__nand2_1 _8230_ (.A(_3431_),
    .B(_3432_),
    .Y(_3433_));
 sky130_fd_sc_hd__a21oi_1 _8231_ (.A1(_3427_),
    .A2(_3433_),
    .B1(_0600_),
    .Y(_3434_));
 sky130_fd_sc_hd__o21ai_1 _8232_ (.A1(_3427_),
    .A2(_3433_),
    .B1(_3434_),
    .Y(_3436_));
 sky130_fd_sc_hd__inv_2 _8233_ (.A(_3234_),
    .Y(_3437_));
 sky130_fd_sc_hd__and2_1 _8234_ (.A(_2993_),
    .B(_3234_),
    .X(_3438_));
 sky130_fd_sc_hd__a21oi_1 _8235_ (.A1(_3437_),
    .A2(_3179_),
    .B1(_3438_),
    .Y(_3439_));
 sky130_fd_sc_hd__and2_1 _8236_ (.A(_3391_),
    .B(_3439_),
    .X(_3440_));
 sky130_fd_sc_hd__nor2_1 _8237_ (.A(_3391_),
    .B(_3439_),
    .Y(_3441_));
 sky130_fd_sc_hd__nor2_1 _8238_ (.A(_3440_),
    .B(_3441_),
    .Y(_3442_));
 sky130_fd_sc_hd__a21oi_1 _8239_ (.A1(_3182_),
    .A2(_3396_),
    .B1(_3442_),
    .Y(_3443_));
 sky130_fd_sc_hd__a311o_1 _8240_ (.A1(_3182_),
    .A2(_3396_),
    .A3(_3442_),
    .B1(_3443_),
    .C1(_3303_),
    .X(_3444_));
 sky130_fd_sc_hd__a31o_1 _8241_ (.A1(_3425_),
    .A2(_3436_),
    .A3(_3444_),
    .B1(_3195_),
    .X(_3445_));
 sky130_fd_sc_hd__a22oi_1 _8242_ (.A1(\out_reg[6] ),
    .A2(_3316_),
    .B1(_3197_),
    .B2(\out_reg[7] ),
    .Y(_3447_));
 sky130_fd_sc_hd__a21oi_1 _8243_ (.A1(_3445_),
    .A2(_3447_),
    .B1(_0635_),
    .Y(_0027_));
 sky130_fd_sc_hd__o21a_1 _8244_ (.A1(_3421_),
    .A2(_3415_),
    .B1(_0601_),
    .X(_3448_));
 sky130_fd_sc_hd__or2_1 _8245_ (.A(_2604_),
    .B(_2515_),
    .X(_3449_));
 sky130_fd_sc_hd__buf_2 _8246_ (.A(_3449_),
    .X(_3450_));
 sky130_fd_sc_hd__o21bai_1 _8247_ (.A1(_3419_),
    .A2(_3450_),
    .B1_N(_3416_),
    .Y(_3451_));
 sky130_fd_sc_hd__a21oi_2 _8248_ (.A1(_3419_),
    .A2(_3450_),
    .B1(_3451_),
    .Y(_3452_));
 sky130_fd_sc_hd__xor2_1 _8249_ (.A(_3448_),
    .B(_3452_),
    .X(_3453_));
 sky130_fd_sc_hd__or2_1 _8250_ (.A(_3234_),
    .B(_3164_),
    .X(_3454_));
 sky130_fd_sc_hd__and3_1 _8251_ (.A(_3391_),
    .B(_3439_),
    .C(_3454_),
    .X(_3455_));
 sky130_fd_sc_hd__o21bai_1 _8252_ (.A1(_3440_),
    .A2(_3454_),
    .B1_N(_3438_),
    .Y(_3457_));
 sky130_fd_sc_hd__nor2_1 _8253_ (.A(_3455_),
    .B(_3457_),
    .Y(_3458_));
 sky130_fd_sc_hd__o31a_1 _8254_ (.A1(_3394_),
    .A2(_3395_),
    .A3(_3442_),
    .B1(_3182_),
    .X(_3459_));
 sky130_fd_sc_hd__nor2_2 _8255_ (.A(_3458_),
    .B(_3459_),
    .Y(_3460_));
 sky130_fd_sc_hd__a21o_1 _8256_ (.A1(_3458_),
    .A2(_3459_),
    .B1(_3303_),
    .X(_3461_));
 sky130_fd_sc_hd__nand2_1 _8257_ (.A(_3426_),
    .B(_3433_),
    .Y(_3462_));
 sky130_fd_sc_hd__nand2_1 _8258_ (.A(_1319_),
    .B(_3462_),
    .Y(_3463_));
 sky130_fd_sc_hd__nor2_1 _8259_ (.A(_3259_),
    .B(_0528_),
    .Y(_3464_));
 sky130_fd_sc_hd__or2_1 _8260_ (.A(_3431_),
    .B(_3464_),
    .X(_3465_));
 sky130_fd_sc_hd__o21ai_1 _8261_ (.A1(_3429_),
    .A2(_3464_),
    .B1(_3431_),
    .Y(_3466_));
 sky130_fd_sc_hd__and2_1 _8262_ (.A(_3465_),
    .B(_3466_),
    .X(_3468_));
 sky130_fd_sc_hd__xor2_1 _8263_ (.A(_3463_),
    .B(_3468_),
    .X(_3469_));
 sky130_fd_sc_hd__o22ai_1 _8264_ (.A1(_3460_),
    .A2(_3461_),
    .B1(_3469_),
    .B2(_0600_),
    .Y(_3470_));
 sky130_fd_sc_hd__a211o_2 _8265_ (.A1(_3212_),
    .A2(_3453_),
    .B1(_3470_),
    .C1(_1177_),
    .X(_3471_));
 sky130_fd_sc_hd__a21bo_1 _8266_ (.A1(\out_reg[7] ),
    .A2(_3242_),
    .B1_N(_1177_),
    .X(_3472_));
 sky130_fd_sc_hd__a22oi_1 _8267_ (.A1(\out_reg[8] ),
    .A2(_3197_),
    .B1(_3471_),
    .B2(_3472_),
    .Y(_3473_));
 sky130_fd_sc_hd__nor2_1 _8268_ (.A(_1220_),
    .B(_3473_),
    .Y(_0028_));
 sky130_fd_sc_hd__o21ba_1 _8269_ (.A1(_3234_),
    .A2(_3233_),
    .B1_N(_3438_),
    .X(_3474_));
 sky130_fd_sc_hd__nand2_1 _8270_ (.A(_3455_),
    .B(_3474_),
    .Y(_3475_));
 sky130_fd_sc_hd__or2_1 _8271_ (.A(_3455_),
    .B(_3474_),
    .X(_3476_));
 sky130_fd_sc_hd__nand2_1 _8272_ (.A(_3475_),
    .B(_3476_),
    .Y(_3478_));
 sky130_fd_sc_hd__o21ai_1 _8273_ (.A1(_3227_),
    .A2(_3460_),
    .B1(_3478_),
    .Y(_3479_));
 sky130_fd_sc_hd__o31a_1 _8274_ (.A1(_3227_),
    .A2(_3460_),
    .A3(_3478_),
    .B1(_3190_),
    .X(_3480_));
 sky130_fd_sc_hd__o31a_2 _8275_ (.A1(_3421_),
    .A2(_3415_),
    .A3(_3452_),
    .B1(_1308_),
    .X(_3481_));
 sky130_fd_sc_hd__a211o_2 _8276_ (.A1(_2514_),
    .A2(_3203_),
    .B1(_3205_),
    .C1(_2604_),
    .X(_3482_));
 sky130_fd_sc_hd__and2b_1 _8277_ (.A_N(_3416_),
    .B(_3482_),
    .X(_3483_));
 sky130_fd_sc_hd__a21oi_1 _8278_ (.A1(_3419_),
    .A2(_3450_),
    .B1(_3483_),
    .Y(_3484_));
 sky130_fd_sc_hd__a31oi_4 _8279_ (.A1(_3419_),
    .A2(_3450_),
    .A3(_3482_),
    .B1(_3484_),
    .Y(_3485_));
 sky130_fd_sc_hd__nand2_1 _8280_ (.A(_3481_),
    .B(_3485_),
    .Y(_3486_));
 sky130_fd_sc_hd__or2_1 _8281_ (.A(_3481_),
    .B(_3485_),
    .X(_3487_));
 sky130_fd_sc_hd__o21a_1 _8282_ (.A1(_3462_),
    .A2(_3468_),
    .B1(_1319_),
    .X(_3489_));
 sky130_fd_sc_hd__a21oi_1 _8283_ (.A1(_0521_),
    .A2(_3217_),
    .B1(_3429_),
    .Y(_3490_));
 sky130_fd_sc_hd__xnor2_2 _8284_ (.A(_3465_),
    .B(_3490_),
    .Y(_3491_));
 sky130_fd_sc_hd__o21bai_1 _8285_ (.A1(_3489_),
    .A2(_3491_),
    .B1_N(_0599_),
    .Y(_3492_));
 sky130_fd_sc_hd__a21oi_1 _8286_ (.A1(_3489_),
    .A2(_3491_),
    .B1(_3492_),
    .Y(_3493_));
 sky130_fd_sc_hd__a31o_1 _8287_ (.A1(_3212_),
    .A2(_3486_),
    .A3(_3487_),
    .B1(_3493_),
    .X(_3494_));
 sky130_fd_sc_hd__a21oi_2 _8288_ (.A1(_3479_),
    .A2(_3480_),
    .B1(_3494_),
    .Y(_3495_));
 sky130_fd_sc_hd__a22o_1 _8289_ (.A1(\out_reg[8] ),
    .A2(_3316_),
    .B1(_1231_),
    .B2(\out_reg[9] ),
    .X(_3496_));
 sky130_fd_sc_hd__o21ba_1 _8290_ (.A1(_3195_),
    .A2(_3495_),
    .B1_N(_3496_),
    .X(_3497_));
 sky130_fd_sc_hd__nor2_1 _8291_ (.A(_1220_),
    .B(_3497_),
    .Y(_0029_));
 sky130_fd_sc_hd__and2_1 _8292_ (.A(_1319_),
    .B(_3485_),
    .X(_3499_));
 sky130_fd_sc_hd__and2_1 _8293_ (.A(_2611_),
    .B(_3251_),
    .X(_3500_));
 sky130_fd_sc_hd__clkinv_2 _8294_ (.A(_3500_),
    .Y(_3501_));
 sky130_fd_sc_hd__and4_1 _8295_ (.A(_3419_),
    .B(_3450_),
    .C(_3482_),
    .D(_3501_),
    .X(_3502_));
 sky130_fd_sc_hd__nor2_1 _8296_ (.A(_3416_),
    .B(_3500_),
    .Y(_3503_));
 sky130_fd_sc_hd__a31o_1 _8297_ (.A1(_3419_),
    .A2(_3450_),
    .A3(_3482_),
    .B1(_3503_),
    .X(_3504_));
 sky130_fd_sc_hd__and2b_1 _8298_ (.A_N(_3502_),
    .B(_3504_),
    .X(_3505_));
 sky130_fd_sc_hd__o21ai_1 _8299_ (.A1(_3481_),
    .A2(_3499_),
    .B1(_3505_),
    .Y(_3506_));
 sky130_fd_sc_hd__or3_1 _8300_ (.A(_3481_),
    .B(_3505_),
    .C(_3499_),
    .X(_3507_));
 sky130_fd_sc_hd__a21oi_1 _8301_ (.A1(_3437_),
    .A2(_3273_),
    .B1(_3475_),
    .Y(_3508_));
 sky130_fd_sc_hd__a31o_1 _8302_ (.A1(_3437_),
    .A2(_3273_),
    .A3(_3475_),
    .B1(_3438_),
    .X(_3510_));
 sky130_fd_sc_hd__or2_1 _8303_ (.A(_3508_),
    .B(_3510_),
    .X(_3511_));
 sky130_fd_sc_hd__a21o_1 _8304_ (.A1(_3460_),
    .A2(_3478_),
    .B1(_3227_),
    .X(_3512_));
 sky130_fd_sc_hd__nand2_1 _8305_ (.A(_3511_),
    .B(_3512_),
    .Y(_3513_));
 sky130_fd_sc_hd__o21a_1 _8306_ (.A1(_3511_),
    .A2(_3512_),
    .B1(_3190_),
    .X(_3514_));
 sky130_fd_sc_hd__o31a_1 _8307_ (.A1(_3462_),
    .A2(_3468_),
    .A3(_3491_),
    .B1(_1319_),
    .X(_3515_));
 sky130_fd_sc_hd__and2b_1 _8308_ (.A_N(_3465_),
    .B(_3490_),
    .X(_3516_));
 sky130_fd_sc_hd__or2_1 _8309_ (.A(_3259_),
    .B(_3261_),
    .X(_3517_));
 sky130_fd_sc_hd__nand2_1 _8310_ (.A(_3516_),
    .B(_3517_),
    .Y(_3518_));
 sky130_fd_sc_hd__o221a_1 _8311_ (.A1(_0440_),
    .A2(_0521_),
    .B1(_3516_),
    .B2(_3517_),
    .C1(_3518_),
    .X(_3519_));
 sky130_fd_sc_hd__a21oi_1 _8312_ (.A1(_3515_),
    .A2(_3519_),
    .B1(_0599_),
    .Y(_3521_));
 sky130_fd_sc_hd__o21a_1 _8313_ (.A1(_3515_),
    .A2(_3519_),
    .B1(_3521_),
    .X(_3522_));
 sky130_fd_sc_hd__a211o_1 _8314_ (.A1(_3513_),
    .A2(_3514_),
    .B1(_3522_),
    .C1(_0701_),
    .X(_3523_));
 sky130_fd_sc_hd__a31o_1 _8315_ (.A1(_3212_),
    .A2(_3506_),
    .A3(_3507_),
    .B1(_3523_),
    .X(_3524_));
 sky130_fd_sc_hd__a21bo_1 _8316_ (.A1(\out_reg[9] ),
    .A2(_3242_),
    .B1_N(_1177_),
    .X(_3525_));
 sky130_fd_sc_hd__a22oi_1 _8317_ (.A1(\out_reg[10] ),
    .A2(_3197_),
    .B1(_3524_),
    .B2(_3525_),
    .Y(_3526_));
 sky130_fd_sc_hd__nor2_1 _8318_ (.A(_1220_),
    .B(_3526_),
    .Y(_0030_));
 sky130_fd_sc_hd__nand2_1 _8319_ (.A(\out_reg[11] ),
    .B(_3197_),
    .Y(_3527_));
 sky130_fd_sc_hd__or2_1 _8320_ (.A(_2604_),
    .B(_3287_),
    .X(_3528_));
 sky130_fd_sc_hd__xnor2_1 _8321_ (.A(_3502_),
    .B(_3528_),
    .Y(_3529_));
 sky130_fd_sc_hd__nor2_1 _8322_ (.A(_3416_),
    .B(_3529_),
    .Y(_3531_));
 sky130_fd_sc_hd__o21a_1 _8323_ (.A1(_3485_),
    .A2(_3505_),
    .B1(_1308_),
    .X(_3532_));
 sky130_fd_sc_hd__o21ai_1 _8324_ (.A1(_3481_),
    .A2(_3532_),
    .B1(_3531_),
    .Y(_3533_));
 sky130_fd_sc_hd__o311a_1 _8325_ (.A1(_3481_),
    .A2(_3531_),
    .A3(_3532_),
    .B1(_3533_),
    .C1(_3212_),
    .X(_3534_));
 sky130_fd_sc_hd__a21oi_1 _8326_ (.A1(_3437_),
    .A2(_3298_),
    .B1(_3438_),
    .Y(_3535_));
 sky130_fd_sc_hd__and2_1 _8327_ (.A(_3508_),
    .B(_3535_),
    .X(_3536_));
 sky130_fd_sc_hd__nor2_1 _8328_ (.A(_3508_),
    .B(_3535_),
    .Y(_3537_));
 sky130_fd_sc_hd__or2_1 _8329_ (.A(_3536_),
    .B(_3537_),
    .X(_3538_));
 sky130_fd_sc_hd__a31o_1 _8330_ (.A1(_3460_),
    .A2(_3478_),
    .A3(_3511_),
    .B1(_3226_),
    .X(_3539_));
 sky130_fd_sc_hd__xor2_1 _8331_ (.A(_3538_),
    .B(_3539_),
    .X(_3540_));
 sky130_fd_sc_hd__o21bai_1 _8332_ (.A1(_3259_),
    .A2(_3308_),
    .B1_N(_3429_),
    .Y(_3542_));
 sky130_fd_sc_hd__xnor2_1 _8333_ (.A(_3518_),
    .B(_3542_),
    .Y(_3543_));
 sky130_fd_sc_hd__inv_2 _8334_ (.A(_3543_),
    .Y(_3544_));
 sky130_fd_sc_hd__or4_1 _8335_ (.A(_3462_),
    .B(_3468_),
    .C(_3491_),
    .D(_3519_),
    .X(_3545_));
 sky130_fd_sc_hd__a31o_1 _8336_ (.A1(_1319_),
    .A2(_3544_),
    .A3(_3545_),
    .B1(_0599_),
    .X(_3546_));
 sky130_fd_sc_hd__a21o_1 _8337_ (.A1(_1308_),
    .A2(_3545_),
    .B1(_3544_),
    .X(_3547_));
 sky130_fd_sc_hd__and2b_1 _8338_ (.A_N(_3546_),
    .B(_3547_),
    .X(_3548_));
 sky130_fd_sc_hd__a211o_1 _8339_ (.A1(_3190_),
    .A2(_3540_),
    .B1(_3548_),
    .C1(_1177_),
    .X(_3549_));
 sky130_fd_sc_hd__nand2_1 _8340_ (.A(\out_reg[10] ),
    .B(_3242_),
    .Y(_3550_));
 sky130_fd_sc_hd__a2bb2o_1 _8341_ (.A1_N(_3534_),
    .A2_N(_3549_),
    .B1(_3550_),
    .B2(_3195_),
    .X(_3551_));
 sky130_fd_sc_hd__a21oi_1 _8342_ (.A1(_3527_),
    .A2(_3551_),
    .B1(_0635_),
    .Y(_0031_));
 sky130_fd_sc_hd__or2_1 _8343_ (.A(_3518_),
    .B(_3542_),
    .X(_3553_));
 sky130_fd_sc_hd__nor2_1 _8344_ (.A(_3259_),
    .B(_3337_),
    .Y(_3554_));
 sky130_fd_sc_hd__nor2_1 _8345_ (.A(_3553_),
    .B(_3554_),
    .Y(_3555_));
 sky130_fd_sc_hd__a221oi_4 _8346_ (.A1(_0451_),
    .A2(_3259_),
    .B1(_3553_),
    .B2(_3554_),
    .C1(_3555_),
    .Y(_3556_));
 sky130_fd_sc_hd__a21oi_1 _8347_ (.A1(_1330_),
    .A2(_3547_),
    .B1(_3556_),
    .Y(_3557_));
 sky130_fd_sc_hd__a311o_1 _8348_ (.A1(_1330_),
    .A2(_3547_),
    .A3(_3556_),
    .B1(_3557_),
    .C1(_0600_),
    .X(_3558_));
 sky130_fd_sc_hd__or2_1 _8349_ (.A(_3234_),
    .B(_3326_),
    .X(_3559_));
 sky130_fd_sc_hd__and3_1 _8350_ (.A(_3508_),
    .B(_3535_),
    .C(_3559_),
    .X(_3560_));
 sky130_fd_sc_hd__o21bai_1 _8351_ (.A1(_3536_),
    .A2(_3559_),
    .B1_N(_3438_),
    .Y(_3561_));
 sky130_fd_sc_hd__nor2_1 _8352_ (.A(_3560_),
    .B(_3561_),
    .Y(_3563_));
 sky130_fd_sc_hd__o21ai_1 _8353_ (.A1(_3227_),
    .A2(_3538_),
    .B1(_3539_),
    .Y(_3564_));
 sky130_fd_sc_hd__or2_1 _8354_ (.A(_3563_),
    .B(_3564_),
    .X(_3565_));
 sky130_fd_sc_hd__a21oi_1 _8355_ (.A1(_3563_),
    .A2(_3564_),
    .B1(_3303_),
    .Y(_3566_));
 sky130_fd_sc_hd__o21ai_1 _8356_ (.A1(_2569_),
    .A2(_2495_),
    .B1(_3286_),
    .Y(_3567_));
 sky130_fd_sc_hd__a21oi_2 _8357_ (.A1(_2611_),
    .A2(_3567_),
    .B1(_3416_),
    .Y(_3568_));
 sky130_fd_sc_hd__and3_1 _8358_ (.A(_3502_),
    .B(_3528_),
    .C(_3568_),
    .X(_3569_));
 sky130_fd_sc_hd__a21oi_1 _8359_ (.A1(_3502_),
    .A2(_3528_),
    .B1(_3568_),
    .Y(_3570_));
 sky130_fd_sc_hd__nor2_1 _8360_ (.A(_3569_),
    .B(_3570_),
    .Y(_3571_));
 sky130_fd_sc_hd__or3_1 _8361_ (.A(_3166_),
    .B(_3416_),
    .C(_3529_),
    .X(_3572_));
 sky130_fd_sc_hd__or3b_1 _8362_ (.A(_3481_),
    .B(_3532_),
    .C_N(_3572_),
    .X(_3574_));
 sky130_fd_sc_hd__xnor2_1 _8363_ (.A(_3571_),
    .B(_3574_),
    .Y(_3575_));
 sky130_fd_sc_hd__o2bb2a_1 _8364_ (.A1_N(_3565_),
    .A2_N(_3566_),
    .B1(_2621_),
    .B2(_3575_),
    .X(_3576_));
 sky130_fd_sc_hd__a21oi_2 _8365_ (.A1(_3558_),
    .A2(_3576_),
    .B1(_3195_),
    .Y(_3577_));
 sky130_fd_sc_hd__a22o_1 _8366_ (.A1(\out_reg[11] ),
    .A2(_3316_),
    .B1(_3197_),
    .B2(\out_reg[12] ),
    .X(_3578_));
 sky130_fd_sc_hd__o21ba_1 _8367_ (.A1(_3577_),
    .A2(_3578_),
    .B1_N(_1220_),
    .X(_0032_));
 sky130_fd_sc_hd__o21a_1 _8368_ (.A1(_2569_),
    .A2(_3352_),
    .B1(_3286_),
    .X(_3579_));
 sky130_fd_sc_hd__o2111a_1 _8369_ (.A1(_2604_),
    .A2(_3579_),
    .B1(_3502_),
    .C1(_3528_),
    .D1(_3568_),
    .X(_3580_));
 sky130_fd_sc_hd__a311o_1 _8370_ (.A1(_3287_),
    .A2(_3502_),
    .A3(_3568_),
    .B1(_3579_),
    .C1(_2604_),
    .X(_3581_));
 sky130_fd_sc_hd__or3b_1 _8371_ (.A(_3416_),
    .B(_3580_),
    .C_N(_3581_),
    .X(_3582_));
 sky130_fd_sc_hd__or3_1 _8372_ (.A(_3166_),
    .B(_3569_),
    .C(_3570_),
    .X(_3584_));
 sky130_fd_sc_hd__and4bb_1 _8373_ (.A_N(_3481_),
    .B_N(_3532_),
    .C(_3572_),
    .D(_3584_),
    .X(_3585_));
 sky130_fd_sc_hd__xnor2_1 _8374_ (.A(_3582_),
    .B(_3585_),
    .Y(_3586_));
 sky130_fd_sc_hd__a21o_1 _8375_ (.A1(_0521_),
    .A2(_3363_),
    .B1(_3429_),
    .X(_3587_));
 sky130_fd_sc_hd__xor2_1 _8376_ (.A(_3555_),
    .B(_3587_),
    .X(_3588_));
 sky130_fd_sc_hd__o21ai_1 _8377_ (.A1(_3547_),
    .A2(_3556_),
    .B1(_1319_),
    .Y(_3589_));
 sky130_fd_sc_hd__nor2_1 _8378_ (.A(_3588_),
    .B(_3589_),
    .Y(_3590_));
 sky130_fd_sc_hd__nand2_1 _8379_ (.A(_3588_),
    .B(_3589_),
    .Y(_3591_));
 sky130_fd_sc_hd__or3b_1 _8380_ (.A(_3590_),
    .B(_0599_),
    .C_N(_3591_),
    .X(_3592_));
 sky130_fd_sc_hd__a21o_1 _8381_ (.A1(_3437_),
    .A2(_3370_),
    .B1(_3438_),
    .X(_3593_));
 sky130_fd_sc_hd__xnor2_1 _8382_ (.A(_3560_),
    .B(_3593_),
    .Y(_3595_));
 sky130_fd_sc_hd__a21o_1 _8383_ (.A1(_3182_),
    .A2(_3565_),
    .B1(_3595_),
    .X(_3596_));
 sky130_fd_sc_hd__nand2_1 _8384_ (.A(_3190_),
    .B(_3596_),
    .Y(_3597_));
 sky130_fd_sc_hd__a31o_1 _8385_ (.A1(_3182_),
    .A2(_3565_),
    .A3(_3595_),
    .B1(_3597_),
    .X(_3598_));
 sky130_fd_sc_hd__o211a_1 _8386_ (.A1(_2621_),
    .A2(_3586_),
    .B1(_3592_),
    .C1(_3598_),
    .X(_3599_));
 sky130_fd_sc_hd__a22o_1 _8387_ (.A1(\out_reg[12] ),
    .A2(_3316_),
    .B1(_1231_),
    .B2(\out_reg[13] ),
    .X(_3600_));
 sky130_fd_sc_hd__o21ba_1 _8388_ (.A1(_3195_),
    .A2(_3599_),
    .B1_N(_3600_),
    .X(_3601_));
 sky130_fd_sc_hd__nor2_1 _8389_ (.A(_1220_),
    .B(_3601_),
    .Y(_0033_));
 sky130_fd_sc_hd__or2_1 _8390_ (.A(_3166_),
    .B(_3582_),
    .X(_3602_));
 sky130_fd_sc_hd__nor2_1 _8391_ (.A(_2604_),
    .B(_3580_),
    .Y(_3603_));
 sky130_fd_sc_hd__a21o_1 _8392_ (.A1(_3404_),
    .A2(_3603_),
    .B1(_3416_),
    .X(_3605_));
 sky130_fd_sc_hd__a21oi_1 _8393_ (.A1(_3585_),
    .A2(_3602_),
    .B1(_3605_),
    .Y(_3606_));
 sky130_fd_sc_hd__a31o_1 _8394_ (.A1(_3585_),
    .A2(_3602_),
    .A3(_3605_),
    .B1(_2621_),
    .X(_3607_));
 sky130_fd_sc_hd__or2_1 _8395_ (.A(_3606_),
    .B(_3607_),
    .X(_3608_));
 sky130_fd_sc_hd__clkinv_2 _8396_ (.A(_3560_),
    .Y(_3609_));
 sky130_fd_sc_hd__or2_1 _8397_ (.A(_3609_),
    .B(_3593_),
    .X(_3610_));
 sky130_fd_sc_hd__nand2_1 _8398_ (.A(_3182_),
    .B(_3596_),
    .Y(_3611_));
 sky130_fd_sc_hd__a21oi_1 _8399_ (.A1(_2993_),
    .A2(_3610_),
    .B1(_3611_),
    .Y(_3612_));
 sky130_fd_sc_hd__a311o_1 _8400_ (.A1(_2993_),
    .A2(_3610_),
    .A3(_3611_),
    .B1(_3612_),
    .C1(_3303_),
    .X(_3613_));
 sky130_fd_sc_hd__or3_1 _8401_ (.A(_3553_),
    .B(_3554_),
    .C(_3587_),
    .X(_3614_));
 sky130_fd_sc_hd__a31o_1 _8402_ (.A1(_0521_),
    .A2(_3384_),
    .A3(_3614_),
    .B1(_3429_),
    .X(_3616_));
 sky130_fd_sc_hd__nand2_1 _8403_ (.A(_0601_),
    .B(_3591_),
    .Y(_3617_));
 sky130_fd_sc_hd__xnor2_1 _8404_ (.A(_3616_),
    .B(_3617_),
    .Y(_3618_));
 sky130_fd_sc_hd__o21ba_1 _8405_ (.A1(_0600_),
    .A2(_3618_),
    .B1_N(_1177_),
    .X(_3619_));
 sky130_fd_sc_hd__nand2_1 _8406_ (.A(\out_reg[13] ),
    .B(_3242_),
    .Y(_3620_));
 sky130_fd_sc_hd__a32o_1 _8407_ (.A1(_3608_),
    .A2(_3613_),
    .A3(_3619_),
    .B1(_3620_),
    .B2(_3195_),
    .X(_3621_));
 sky130_fd_sc_hd__nand2_1 _8408_ (.A(\out_reg[14] ),
    .B(_3197_),
    .Y(_3622_));
 sky130_fd_sc_hd__a21oi_1 _8409_ (.A1(_3621_),
    .A2(_3622_),
    .B1(_0635_),
    .Y(_0034_));
 sky130_fd_sc_hd__o21ai_1 _8410_ (.A1(_3227_),
    .A2(_3188_),
    .B1(_3187_),
    .Y(_3623_));
 sky130_fd_sc_hd__or3_1 _8411_ (.A(\cmd[7] ),
    .B(\cmd[6] ),
    .C(_3623_),
    .X(_3624_));
 sky130_fd_sc_hd__nand2_1 _8412_ (.A(\cmd[7] ),
    .B(\cmd[6] ),
    .Y(_3626_));
 sky130_fd_sc_hd__nand2_1 _8413_ (.A(_3225_),
    .B(_4250_),
    .Y(_3627_));
 sky130_fd_sc_hd__a22oi_1 _8414_ (.A1(\cmd[6] ),
    .A2(_3186_),
    .B1(_3627_),
    .B2(\cmd[7] ),
    .Y(_3628_));
 sky130_fd_sc_hd__a221o_1 _8415_ (.A1(_1253_),
    .A2(_0082_),
    .B1(_2319_),
    .B2(_1330_),
    .C1(_3628_),
    .X(_3629_));
 sky130_fd_sc_hd__a31o_1 _8416_ (.A1(_3624_),
    .A2(_3626_),
    .A3(_3629_),
    .B1(_1177_),
    .X(_3630_));
 sky130_fd_sc_hd__inv_2 _8417_ (.A(_1231_),
    .Y(_3631_));
 sky130_fd_sc_hd__o22a_1 _8418_ (.A1(\out_reg[14] ),
    .A2(_0797_),
    .B1(_3631_),
    .B2(\out_reg[15] ),
    .X(_3632_));
 sky130_fd_sc_hd__and3b_1 _8419_ (.A_N(_0635_),
    .B(_3630_),
    .C(_3632_),
    .X(_3633_));
 sky130_fd_sc_hd__clkbuf_1 _8420_ (.A(_3633_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _8421_ (.A0(\out_reg[15] ),
    .A1(io_out[3]),
    .S(_0819_),
    .X(_3634_));
 sky130_fd_sc_hd__clkbuf_1 _8422_ (.A(_3634_),
    .X(_0036_));
 sky130_fd_sc_hd__clkinv_2 _8423_ (.A(mode),
    .Y(_3636_));
 sky130_fd_sc_hd__or4b_1 _8424_ (.A(\counter[3] ),
    .B(_3636_),
    .C(_0668_),
    .D_N(\counter[4] ),
    .X(_3637_));
 sky130_fd_sc_hd__inv_2 _8425_ (.A(_3637_),
    .Y(_3638_));
 sky130_fd_sc_hd__or3b_1 _8426_ (.A(_0635_),
    .B(_3638_),
    .C_N(_0701_),
    .X(_3639_));
 sky130_fd_sc_hd__a21oi_1 _8427_ (.A1(\in_reg[1] ),
    .A2(_0679_),
    .B1(mode),
    .Y(_3640_));
 sky130_fd_sc_hd__nor2_1 _8428_ (.A(_3639_),
    .B(_3640_),
    .Y(_0037_));
 sky130_fd_sc_hd__nor2_1 _8429_ (.A(_0679_),
    .B(_3639_),
    .Y(_3641_));
 sky130_fd_sc_hd__o21ai_1 _8430_ (.A1(\counter[0] ),
    .A2(_3242_),
    .B1(_3641_),
    .Y(_3642_));
 sky130_fd_sc_hd__a21oi_1 _8431_ (.A1(\counter[0] ),
    .A2(_3242_),
    .B1(_3642_),
    .Y(_0038_));
 sky130_fd_sc_hd__and3_1 _8432_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .C(_0786_),
    .X(_3644_));
 sky130_fd_sc_hd__a21o_1 _8433_ (.A1(\counter[0] ),
    .A2(_3242_),
    .B1(\counter[1] ),
    .X(_3645_));
 sky130_fd_sc_hd__and3b_1 _8434_ (.A_N(_3644_),
    .B(_3645_),
    .C(_3641_),
    .X(_3646_));
 sky130_fd_sc_hd__clkbuf_1 _8435_ (.A(_3646_),
    .X(_0039_));
 sky130_fd_sc_hd__o21ai_1 _8436_ (.A1(\counter[2] ),
    .A2(_3644_),
    .B1(_3641_),
    .Y(_3647_));
 sky130_fd_sc_hd__a21oi_1 _8437_ (.A1(\counter[2] ),
    .A2(_3644_),
    .B1(_3647_),
    .Y(_0040_));
 sky130_fd_sc_hd__and3_1 _8438_ (.A(\counter[3] ),
    .B(\counter[2] ),
    .C(_3644_),
    .X(_3648_));
 sky130_fd_sc_hd__a21o_1 _8439_ (.A1(\counter[2] ),
    .A2(_3644_),
    .B1(\counter[3] ),
    .X(_3649_));
 sky130_fd_sc_hd__and3b_1 _8440_ (.A_N(_3648_),
    .B(_3641_),
    .C(_3649_),
    .X(_3650_));
 sky130_fd_sc_hd__clkbuf_1 _8441_ (.A(_3650_),
    .X(_0041_));
 sky130_fd_sc_hd__a211o_1 _8442_ (.A1(\counter[4] ),
    .A2(_3648_),
    .B1(_3639_),
    .C1(_0679_),
    .X(_3652_));
 sky130_fd_sc_hd__o21ba_1 _8443_ (.A1(\counter[4] ),
    .A2(_3648_),
    .B1_N(_3652_),
    .X(_0042_));
 sky130_fd_sc_hd__or4b_1 _8444_ (.A(net4),
    .B(\cmd[0] ),
    .C(_3637_),
    .D_N(net1),
    .X(_3653_));
 sky130_fd_sc_hd__clkbuf_4 _8445_ (.A(_3653_),
    .X(_3654_));
 sky130_fd_sc_hd__buf_4 _8446_ (.A(_3654_),
    .X(_3655_));
 sky130_fd_sc_hd__mux2_1 _8447_ (.A0(\in_reg[0] ),
    .A1(_2969_),
    .S(_3655_),
    .X(_3656_));
 sky130_fd_sc_hd__clkbuf_1 _8448_ (.A(_3656_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _8449_ (.A0(\in_reg[1] ),
    .A1(\posit_add.in1[1] ),
    .S(_3655_),
    .X(_3657_));
 sky130_fd_sc_hd__clkbuf_1 _8450_ (.A(_3657_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _8451_ (.A0(\in_reg[2] ),
    .A1(\posit_add.in1[2] ),
    .S(_3655_),
    .X(_3658_));
 sky130_fd_sc_hd__clkbuf_1 _8452_ (.A(_3658_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _8453_ (.A0(\in_reg[3] ),
    .A1(\posit_add.in1[3] ),
    .S(_3655_),
    .X(_3660_));
 sky130_fd_sc_hd__clkbuf_1 _8454_ (.A(_3660_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _8455_ (.A0(\in_reg[4] ),
    .A1(\posit_add.in1[4] ),
    .S(_3655_),
    .X(_3661_));
 sky130_fd_sc_hd__clkbuf_1 _8456_ (.A(_3661_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _8457_ (.A0(\in_reg[5] ),
    .A1(\posit_add.in1[5] ),
    .S(_3655_),
    .X(_3662_));
 sky130_fd_sc_hd__clkbuf_1 _8458_ (.A(_3662_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _8459_ (.A0(\in_reg[6] ),
    .A1(\posit_add.in1[6] ),
    .S(_3655_),
    .X(_3663_));
 sky130_fd_sc_hd__clkbuf_1 _8460_ (.A(_3663_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _8461_ (.A0(\in_reg[7] ),
    .A1(\posit_add.in1[7] ),
    .S(_3655_),
    .X(_3664_));
 sky130_fd_sc_hd__clkbuf_1 _8462_ (.A(_3664_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _8463_ (.A0(\in_reg[8] ),
    .A1(\posit_add.in1[8] ),
    .S(_3655_),
    .X(_3666_));
 sky130_fd_sc_hd__clkbuf_1 _8464_ (.A(_3666_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _8465_ (.A0(\in_reg[9] ),
    .A1(\posit_add.in1[9] ),
    .S(_3655_),
    .X(_3667_));
 sky130_fd_sc_hd__clkbuf_1 _8466_ (.A(_3667_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _8467_ (.A0(\in_reg[10] ),
    .A1(\posit_add.in1[10] ),
    .S(_3654_),
    .X(_3668_));
 sky130_fd_sc_hd__clkbuf_1 _8468_ (.A(_3668_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _8469_ (.A0(\in_reg[11] ),
    .A1(\posit_add.in1[11] ),
    .S(_3654_),
    .X(_3669_));
 sky130_fd_sc_hd__clkbuf_1 _8470_ (.A(_3669_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _8471_ (.A0(\in_reg[12] ),
    .A1(\posit_add.in1[12] ),
    .S(_3654_),
    .X(_3670_));
 sky130_fd_sc_hd__clkbuf_1 _8472_ (.A(_3670_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _8473_ (.A0(\in_reg[13] ),
    .A1(\posit_add.in1[13] ),
    .S(_3654_),
    .X(_3672_));
 sky130_fd_sc_hd__clkbuf_1 _8474_ (.A(_3672_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _8475_ (.A0(\in_reg[14] ),
    .A1(\posit_add.in1[14] ),
    .S(_3654_),
    .X(_3673_));
 sky130_fd_sc_hd__clkbuf_1 _8476_ (.A(_3673_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _8477_ (.A0(\in_reg[15] ),
    .A1(_1253_),
    .S(_3654_),
    .X(_3674_));
 sky130_fd_sc_hd__clkbuf_1 _8478_ (.A(_3674_),
    .X(_0058_));
 sky130_fd_sc_hd__and4b_1 _8479_ (.A_N(net4),
    .B(\cmd[0] ),
    .C(_3638_),
    .D(net1),
    .X(_3675_));
 sky130_fd_sc_hd__clkbuf_4 _8480_ (.A(_3675_),
    .X(_3676_));
 sky130_fd_sc_hd__clkbuf_4 _8481_ (.A(_3676_),
    .X(_3677_));
 sky130_fd_sc_hd__mux2_1 _8482_ (.A0(\posit_add.in2[0] ),
    .A1(\in_reg[0] ),
    .S(_3677_),
    .X(_3679_));
 sky130_fd_sc_hd__clkbuf_1 _8483_ (.A(_3679_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _8484_ (.A0(\posit_add.in2[1] ),
    .A1(\in_reg[1] ),
    .S(_3677_),
    .X(_3680_));
 sky130_fd_sc_hd__clkbuf_1 _8485_ (.A(_3680_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _8486_ (.A0(\posit_add.in2[2] ),
    .A1(\in_reg[2] ),
    .S(_3677_),
    .X(_3681_));
 sky130_fd_sc_hd__clkbuf_1 _8487_ (.A(_3681_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _8488_ (.A0(\posit_add.in2[3] ),
    .A1(\in_reg[3] ),
    .S(_3677_),
    .X(_3682_));
 sky130_fd_sc_hd__clkbuf_1 _8489_ (.A(_3682_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _8490_ (.A0(\posit_add.in2[4] ),
    .A1(\in_reg[4] ),
    .S(_3677_),
    .X(_3683_));
 sky130_fd_sc_hd__clkbuf_1 _8491_ (.A(_3683_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _8492_ (.A0(\posit_add.in2[5] ),
    .A1(\in_reg[5] ),
    .S(_3677_),
    .X(_3685_));
 sky130_fd_sc_hd__clkbuf_1 _8493_ (.A(_3685_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _8494_ (.A0(\posit_add.in2[6] ),
    .A1(\in_reg[6] ),
    .S(_3677_),
    .X(_3686_));
 sky130_fd_sc_hd__clkbuf_1 _8495_ (.A(_3686_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _8496_ (.A0(\posit_add.in2[7] ),
    .A1(\in_reg[7] ),
    .S(_3677_),
    .X(_3687_));
 sky130_fd_sc_hd__clkbuf_1 _8497_ (.A(_3687_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _8498_ (.A0(\posit_add.in2[8] ),
    .A1(\in_reg[8] ),
    .S(_3677_),
    .X(_3688_));
 sky130_fd_sc_hd__clkbuf_1 _8499_ (.A(_3688_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _8500_ (.A0(\posit_add.in2[9] ),
    .A1(\in_reg[9] ),
    .S(_3677_),
    .X(_3689_));
 sky130_fd_sc_hd__clkbuf_1 _8501_ (.A(_3689_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _8502_ (.A0(\posit_add.in2[10] ),
    .A1(\in_reg[10] ),
    .S(_3676_),
    .X(_3691_));
 sky130_fd_sc_hd__clkbuf_1 _8503_ (.A(_3691_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _8504_ (.A0(\posit_add.in2[11] ),
    .A1(\in_reg[11] ),
    .S(_3676_),
    .X(_3692_));
 sky130_fd_sc_hd__clkbuf_1 _8505_ (.A(_3692_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _8506_ (.A0(\posit_add.in2[12] ),
    .A1(\in_reg[12] ),
    .S(_3676_),
    .X(_3693_));
 sky130_fd_sc_hd__clkbuf_1 _8507_ (.A(_3693_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _8508_ (.A0(\posit_add.in2[13] ),
    .A1(\in_reg[13] ),
    .S(_3676_),
    .X(_3694_));
 sky130_fd_sc_hd__clkbuf_1 _8509_ (.A(_3694_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _8510_ (.A0(\posit_add.in2[14] ),
    .A1(\in_reg[14] ),
    .S(_3676_),
    .X(_3695_));
 sky130_fd_sc_hd__clkbuf_1 _8511_ (.A(_3695_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _8512_ (.A0(_1275_),
    .A1(\in_reg[15] ),
    .S(_3676_),
    .X(_3697_));
 sky130_fd_sc_hd__clkbuf_1 _8513_ (.A(_3697_),
    .X(_0074_));
 sky130_fd_sc_hd__dfxtp_1 _8514_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0000_),
    .Q(\cmd[0] ));
 sky130_fd_sc_hd__dfxtp_4 _8515_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0001_),
    .Q(\cmd[6] ));
 sky130_fd_sc_hd__dfxtp_4 _8516_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0002_),
    .Q(\cmd[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8517_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0003_),
    .Q(\in_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8518_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0004_),
    .Q(\in_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8519_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0005_),
    .Q(\in_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8520_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0006_),
    .Q(\in_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8521_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0007_),
    .Q(\in_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8522_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0008_),
    .Q(\in_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8523_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0009_),
    .Q(\in_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8524_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0010_),
    .Q(\in_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8525_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0011_),
    .Q(\in_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8526_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0012_),
    .Q(\in_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8527_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0013_),
    .Q(\in_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8528_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0014_),
    .Q(\in_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8529_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0015_),
    .Q(\in_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8530_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0016_),
    .Q(\in_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8531_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0017_),
    .Q(\in_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8532_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0018_),
    .Q(\in_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8533_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0019_),
    .Q(last_SCLK));
 sky130_fd_sc_hd__dfxtp_1 _8534_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0020_),
    .Q(\out_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8535_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0021_),
    .Q(\out_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8536_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0022_),
    .Q(\out_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8537_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0023_),
    .Q(\out_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8538_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0024_),
    .Q(\out_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8539_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0025_),
    .Q(\out_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8540_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0026_),
    .Q(\out_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8541_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0027_),
    .Q(\out_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8542_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0028_),
    .Q(\out_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8543_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0029_),
    .Q(\out_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8544_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0030_),
    .Q(\out_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8545_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0031_),
    .Q(\out_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8546_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0032_),
    .Q(\out_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8547_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0033_),
    .Q(\out_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8548_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0034_),
    .Q(\out_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8549_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0035_),
    .Q(\out_reg[15] ));
 sky130_fd_sc_hd__dfxtp_2 _8550_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0036_),
    .Q(io_out[3]));
 sky130_fd_sc_hd__dfxtp_1 _8551_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0037_),
    .Q(mode));
 sky130_fd_sc_hd__dfxtp_1 _8552_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0038_),
    .Q(\counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8553_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0039_),
    .Q(\counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8554_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0040_),
    .Q(\counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8555_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0041_),
    .Q(\counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8556_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0042_),
    .Q(\counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8557_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0043_),
    .Q(\posit_add.in1[0] ));
 sky130_fd_sc_hd__dfxtp_4 _8558_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0044_),
    .Q(\posit_add.in1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _8559_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0045_),
    .Q(\posit_add.in1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _8560_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0046_),
    .Q(\posit_add.in1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _8561_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0047_),
    .Q(\posit_add.in1[4] ));
 sky130_fd_sc_hd__dfxtp_2 _8562_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0048_),
    .Q(\posit_add.in1[5] ));
 sky130_fd_sc_hd__dfxtp_2 _8563_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0049_),
    .Q(\posit_add.in1[6] ));
 sky130_fd_sc_hd__dfxtp_2 _8564_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0050_),
    .Q(\posit_add.in1[7] ));
 sky130_fd_sc_hd__dfxtp_2 _8565_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0051_),
    .Q(\posit_add.in1[8] ));
 sky130_fd_sc_hd__dfxtp_2 _8566_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0052_),
    .Q(\posit_add.in1[9] ));
 sky130_fd_sc_hd__dfxtp_2 _8567_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0053_),
    .Q(\posit_add.in1[10] ));
 sky130_fd_sc_hd__dfxtp_2 _8568_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0054_),
    .Q(\posit_add.in1[11] ));
 sky130_fd_sc_hd__dfxtp_2 _8569_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0055_),
    .Q(\posit_add.in1[12] ));
 sky130_fd_sc_hd__dfxtp_2 _8570_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0056_),
    .Q(\posit_add.in1[13] ));
 sky130_fd_sc_hd__dfxtp_4 _8571_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0057_),
    .Q(\posit_add.in1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8572_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0058_),
    .Q(\posit_add.in1[15] ));
 sky130_fd_sc_hd__dfxtp_2 _8573_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0059_),
    .Q(\posit_add.in2[0] ));
 sky130_fd_sc_hd__dfxtp_2 _8574_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0060_),
    .Q(\posit_add.in2[1] ));
 sky130_fd_sc_hd__dfxtp_2 _8575_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0061_),
    .Q(\posit_add.in2[2] ));
 sky130_fd_sc_hd__dfxtp_2 _8576_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0062_),
    .Q(\posit_add.in2[3] ));
 sky130_fd_sc_hd__dfxtp_2 _8577_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0063_),
    .Q(\posit_add.in2[4] ));
 sky130_fd_sc_hd__dfxtp_2 _8578_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0064_),
    .Q(\posit_add.in2[5] ));
 sky130_fd_sc_hd__dfxtp_2 _8579_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0065_),
    .Q(\posit_add.in2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8580_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0066_),
    .Q(\posit_add.in2[7] ));
 sky130_fd_sc_hd__dfxtp_2 _8581_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0067_),
    .Q(\posit_add.in2[8] ));
 sky130_fd_sc_hd__dfxtp_2 _8582_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0068_),
    .Q(\posit_add.in2[9] ));
 sky130_fd_sc_hd__dfxtp_2 _8583_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0069_),
    .Q(\posit_add.in2[10] ));
 sky130_fd_sc_hd__dfxtp_2 _8584_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0070_),
    .Q(\posit_add.in2[11] ));
 sky130_fd_sc_hd__dfxtp_2 _8585_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0071_),
    .Q(\posit_add.in2[12] ));
 sky130_fd_sc_hd__dfxtp_2 _8586_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0072_),
    .Q(\posit_add.in2[13] ));
 sky130_fd_sc_hd__dfxtp_4 _8587_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0073_),
    .Q(\posit_add.in2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8588_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0074_),
    .Q(\posit_add.in2[15] ));
 sky130_fd_sc_hd__conb_1 posit_unit_6 (.LO(net6));
 sky130_fd_sc_hd__conb_1 posit_unit_7 (.LO(net7));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(rst),
    .X(net4));
 sky130_fd_sc_hd__conb_1 posit_unit_5 (.LO(net5));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7682__A1 (.DIODE(_0080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7172__A (.DIODE(_0080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7169__A (.DIODE(_0080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A (.DIODE(_0080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A (.DIODE(_0080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A1 (.DIODE(_0080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A (.DIODE(_0080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__A (.DIODE(_0080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__A (.DIODE(_0080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A1 (.DIODE(_0080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8415__A2 (.DIODE(_0082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7687__A2 (.DIODE(_0082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7238__B (.DIODE(_0082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7193__A1 (.DIODE(_0082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__A (.DIODE(_0082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__B (.DIODE(_0082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6502__A (.DIODE(_0082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A (.DIODE(_0082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A2 (.DIODE(_0082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A2 (.DIODE(_0082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7484__B (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7220__A2 (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A1 (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__A (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__C (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__B (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__B (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__B1 (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__C (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7593__A0 (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7587__A1 (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__A3 (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__A1 (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A1 (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__B2 (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__C (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8000__A2 (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7180__C (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__B (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__A2_N (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__B2 (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A2 (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A2 (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__B (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__D (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__B (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7620__A1 (.DIODE(_0147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7614__A0 (.DIODE(_0147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7343__A1 (.DIODE(_0147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7102__A (.DIODE(_0147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__A (.DIODE(_0147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__A (.DIODE(_0147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__C (.DIODE(_0147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__C (.DIODE(_0147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__B (.DIODE(_0147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A2 (.DIODE(_0147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7570__A0 (.DIODE(_0218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7385__A1 (.DIODE(_0218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__A (.DIODE(_0218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__A (.DIODE(_0218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__A1 (.DIODE(_0218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__A (.DIODE(_0218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A (.DIODE(_0218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A1 (.DIODE(_0218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7170__B (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__A1 (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__A (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__A (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__A (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__A (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__B (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__A (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A2 (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7548__B2 (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7270__A1 (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__A1 (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__A (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7529__A (.DIODE(_0369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7231__A (.DIODE(_0369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__A (.DIODE(_0369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A (.DIODE(_0369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7527__A (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__A (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__C1 (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8311__A1 (.DIODE(_0440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8226__A (.DIODE(_0440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8068__A0 (.DIODE(_0440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A2 (.DIODE(_0440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__A (.DIODE(_0440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__D1 (.DIODE(_0440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__A (.DIODE(_0440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__B (.DIODE(_0440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A (.DIODE(_0440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__B (.DIODE(_0440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A1 (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__A1 (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__D (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8346__A1 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8111__A (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8026__A0 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__B1 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__B (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__B (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__B1_N (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7417__B (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7414__A (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__B (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__B (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__A2 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__B (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__B (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__A (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__B (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A2 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8405__A1 (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8348__C1 (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8264__B2 (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8231__B1 (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8209__A1 (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8170__C1 (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8116__B1 (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8076__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8034__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8006__A2 (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6339__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__A1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__C (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__B (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7294__B (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7223__B (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__A1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A2 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7294__A_N (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7223__A_N (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__B2 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8426__C_N (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8314__C1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8119__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8087__B1_N (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8086__B1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8052__B1_N (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8050__B1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__B_N (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__C_N (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__B (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A1_N (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__C1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__A2 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__C (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__A2 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__B (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__C (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__B (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__A1 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__A (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__B2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__A (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__A1 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__B1 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__A4 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__A2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__S (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__S (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__S (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A1 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6320__B2 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__A (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__A (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__B (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A2 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__B2 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__A2 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6021__B1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__B (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__B1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6320__A1 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__B2 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__B (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__B (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A2 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__B (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6009__C (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__B (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__B (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A2 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__B (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__A (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__A1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__A (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__A1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__C (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__B1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__A1 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__A1 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__A1 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__A (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A1 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__A (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__A1 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__A (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__A (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__A2 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8421__S (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__S (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__S (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__S (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__S (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__S (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__S (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__A (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__S (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__S (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__S (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__S (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__S (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__S (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__S (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__S (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__S (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4276__S (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__D (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__A (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__A1 (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__B2 (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__A1 (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__D_N (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__A (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__B_N (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__A (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__B_N (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__B2 (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__A (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__B (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__B (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__A2 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__B1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__B (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A2 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__B (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__B (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__D1 (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__B (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__A2 (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__B (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__A2 (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__B (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__B (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__B2 (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__A (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__B (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8416__B1 (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8405__B1_N (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8339__C1 (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8316__B1_N (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8266__B1_N (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8265__C1 (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8149__B1_N (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8148__D1 (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8007__A (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__S (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8477__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8415__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7998__A (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7995__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7765__A (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__B1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__A (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__B1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__B1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__A (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8512__A0 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8035__A (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7999__A (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7995__A0 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7765__B (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__B (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__A (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__B1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__A (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__B (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7751__S (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7748__A1 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7747__A (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7745__S (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7743__S (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7739__S (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7732__S (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7729__A1 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7686__B1 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__A (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8337__A1 (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8323__B1 (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8275__B1 (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7783__A (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7763__A (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7759__S (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7757__A1 (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7756__A (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7475__B1 (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__A (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8415__B2 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8348__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8347__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8220__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8170__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8169__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8158__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8115__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8033__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__B (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__B (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__C (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__C (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7604__A1 (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7597__A0 (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__B (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__B (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__A1_N (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__C (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__A (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__A (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__A (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__A (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__B (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__A (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__A (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__A (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__A (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7611__A1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__A1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__A (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__A (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__A (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__B2 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__B (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__B (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__B (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__A (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__A (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__A (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__B (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__A (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__A (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__A (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__A1 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__B (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__B (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__A (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__A (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__A (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__A (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__A (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6980__A (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6979__A (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6950__A (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__A (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__B (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__B (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__B (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__B (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__B (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__A (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__A (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__A (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__A (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__A2_N (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__B (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__B (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__B1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__B (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__B (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__A (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__A (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__B1 (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__A0 (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__A (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__A (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__A1 (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__A (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__A (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__A1 (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__A (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__B (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__B (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__B (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__B (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__B (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__B (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7351__A1 (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__A (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__A (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__A1 (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__A (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__A (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__B (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__B (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__B (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__B (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7193__A2 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7169__B (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__A (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__B (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__B (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__B (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__A (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__A (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__A (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__A (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7065__A (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__A (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__A (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__A (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6978__A (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__A (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__B (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__B (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__B (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__B (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7315__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__B (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7043__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__A (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__B (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__B (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__B (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__B (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__D (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__A1 (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__A1 (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__B (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__B (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__B (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__A2 (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__B (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__B (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__B (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__B (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7640__A0 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7418__A1 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7129__A (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__A (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__B (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__B (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__B (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6881__C (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__A2 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__B1 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__A2 (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__B (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__C (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7043__A2 (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__C (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__B (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6979__B (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__B (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__B (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__A (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__A2 (.DIODE(_1538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__C (.DIODE(_1538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__C (.DIODE(_1538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6980__B (.DIODE(_1538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__A2 (.DIODE(_1538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__B (.DIODE(_1538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__B (.DIODE(_1538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__B (.DIODE(_1538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__B (.DIODE(_1538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6502__B (.DIODE(_1538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__A1 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__A1_N (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__A (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__A1 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__A (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7306__A1 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7131__A2 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__A (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__A1 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__A (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__B (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__B (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__B (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__B (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__A2 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7502__A2 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7501__A2 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__A1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__C1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__A1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__B1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4355__B1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__A (.DIODE(_1711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__A (.DIODE(_1711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__A (.DIODE(_1711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__B (.DIODE(_1711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__A (.DIODE(_1711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__B (.DIODE(_1711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__A2 (.DIODE(_1711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__B (.DIODE(_1718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__B (.DIODE(_1718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6978__B (.DIODE(_1718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6950__B (.DIODE(_1718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__B (.DIODE(_1718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__A2 (.DIODE(_1718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__B (.DIODE(_1718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__B (.DIODE(_1718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__B (.DIODE(_1718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__B (.DIODE(_1718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A1 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__B1 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A2 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__B2 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__B1 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__C (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__A (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7540__B (.DIODE(_1781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A (.DIODE(_1781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A (.DIODE(_1781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__B (.DIODE(_1781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A (.DIODE(_1781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A (.DIODE(_1781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__B (.DIODE(_1781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__A (.DIODE(_1781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__A (.DIODE(_1781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A (.DIODE(_1781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__A (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__A1 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__B (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__A (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__B (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__B (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__B (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6842__C (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__A2 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__C (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7495__B1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7494__A2 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__A1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__C (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__B (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__B (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7498__B1 (.DIODE(_1858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7497__A2 (.DIODE(_1858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A1 (.DIODE(_1858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__A1 (.DIODE(_1858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__C1 (.DIODE(_1858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__B (.DIODE(_1858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__A2 (.DIODE(_1858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__B (.DIODE(_1858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7492__A (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__A1 (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__C1 (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__A1 (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__B (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__B (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__A1 (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__A1 (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__C1 (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__B (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__C (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__C (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__B (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__C (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__C (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7154__A_N (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__B (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8415__B1 (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8022__B (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7586__A0 (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7567__A (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7565__A (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7212__B (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7312__A (.DIODE(_2333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7224__C (.DIODE(_2333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7398__B2 (.DIODE(_2335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7375__A (.DIODE(_2335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7350__A (.DIODE(_2335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7326__B2 (.DIODE(_2335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7306__B1 (.DIODE(_2335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7227__B (.DIODE(_2335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__B (.DIODE(_2335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7287__A1 (.DIODE(_2349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7277__A (.DIODE(_2349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7239__A (.DIODE(_2349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7272__B1_N (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7258__A1 (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7242__B1 (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7288__B (.DIODE(_2354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7284__A2_N (.DIODE(_2354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7272__A2 (.DIODE(_2354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7271__B (.DIODE(_2354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7247__A (.DIODE(_2354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7477__A1 (.DIODE(_2381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7457__A1 (.DIODE(_2381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7386__A1 (.DIODE(_2381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7269__A (.DIODE(_2381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7462__A1 (.DIODE(_2382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7456__B1 (.DIODE(_2382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7366__A1 (.DIODE(_2382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7269__B (.DIODE(_2382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7295__A (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7405__B1 (.DIODE(_2412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7374__A (.DIODE(_2412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7351__A2 (.DIODE(_2412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7318__B (.DIODE(_2412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7315__A2 (.DIODE(_2412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7306__A2 (.DIODE(_2412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7304__B1 (.DIODE(_2412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7426__S (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7410__B2 (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7407__B2 (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7376__B2 (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7338__A (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7322__A (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7318__A (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7314__S (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7305__A_N (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7398__A2_N (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7323__B1 (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__B (.DIODE(_2452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__B (.DIODE(_2452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__B (.DIODE(_2452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__S (.DIODE(_2452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A2 (.DIODE(_2452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__A3 (.DIODE(_2452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__C (.DIODE(_2452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__A2 (.DIODE(_2452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__A2 (.DIODE(_2452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__A2 (.DIODE(_2452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7478__A0 (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7365__B1 (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A1 (.DIODE(_2507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A1 (.DIODE(_2507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__A (.DIODE(_2507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__B2 (.DIODE(_2507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A (.DIODE(_2507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A2 (.DIODE(_2507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A2 (.DIODE(_2507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__B (.DIODE(_2507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__B (.DIODE(_2507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7407__A2 (.DIODE(_2524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7398__B1 (.DIODE(_2524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A (.DIODE(_2529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A (.DIODE(_2529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__A (.DIODE(_2529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A1 (.DIODE(_2529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A (.DIODE(_2529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__B1 (.DIODE(_2529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__A (.DIODE(_2529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__A (.DIODE(_2529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__A (.DIODE(_2529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__A (.DIODE(_2529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7409__A (.DIODE(_2534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7407__B1 (.DIODE(_2534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7424__A (.DIODE(_2536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7410__A2 (.DIODE(_2536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A1 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A1 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__B (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__A (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A1 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__A (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__A (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__A1 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7428__B1 (.DIODE(_2557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8394__B1 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8386__A1 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8364__B1 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8221__B1 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8207__B1 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8159__B1 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8098__B1 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8005__A2 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7624__S (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7614__S (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7606__S (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7587__S (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7571__S (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7569__A (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7544__S (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7542__S (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7520__S (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7514__S (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7613__B (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7601__B (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7595__B (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7584__A (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7572__C_N (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7568__A (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7563__A (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7560__B (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8036__S (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7995__S (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7795__A2 (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7789__S (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7682__S (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7620__S (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7611__S (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7604__S (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7593__S (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7577__S (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7718__B (.DIODE(_2780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7631__A (.DIODE(_2780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7714__B1 (.DIODE(_2800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7660__B (.DIODE(_2800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7649__B (.DIODE(_2800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7712__B (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7694__B (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7659__A_N (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7727__B1 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7684__B (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7683__B (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7498__B2 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7497__A1 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__A1 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__A1 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__B1 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__B (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7947__A1 (.DIODE(_2937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7937__S (.DIODE(_2937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7932__A1 (.DIODE(_2937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7883__A (.DIODE(_2937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7874__B (.DIODE(_2937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7778__B (.DIODE(_2937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7773__B (.DIODE(_2937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7945__C1 (.DIODE(_2941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7883__B (.DIODE(_2941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7880__A (.DIODE(_2941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7864__A (.DIODE(_2941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7791__B (.DIODE(_2941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7777__B (.DIODE(_2941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7900__A_N (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7893__S (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7879__S (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7870__A (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7866__A (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7794__A (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7790__A (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8447__A1 (.DIODE(_2969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7493__C1 (.DIODE(_2969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__C1 (.DIODE(_2969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A1 (.DIODE(_2969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__A1 (.DIODE(_2969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A1 (.DIODE(_2969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__A (.DIODE(_2969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A1 (.DIODE(_2969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__A (.DIODE(_2969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__A (.DIODE(_2969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7821__A (.DIODE(_2980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7238__A (.DIODE(_2980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__B1 (.DIODE(_2980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__B1 (.DIODE(_2980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A2 (.DIODE(_2980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__A (.DIODE(_2980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__A (.DIODE(_2980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__D (.DIODE(_2980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8400__A1 (.DIODE(_2993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8399__A1 (.DIODE(_2993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8234__A (.DIODE(_2993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8040__A1 (.DIODE(_2993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7855__A (.DIODE(_2993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7853__A (.DIODE(_2993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7844__B1 (.DIODE(_2993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7827__A (.DIODE(_2993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7826__A (.DIODE(_2993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7984__B2 (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7966__S (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7962__S (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7958__S (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7957__S (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7921__S (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7908__S (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7888__S (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7876__S (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7859__A1 (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8398__A (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8385__A1 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8383__A1 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8254__B1 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8240__A1 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8239__A1 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8194__B1 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8175__A (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8003__A3 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7997__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7495__B2 (.DIODE(_3189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7494__A1 (.DIODE(_3189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__B1 (.DIODE(_3189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__A1 (.DIODE(_3189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__A1 (.DIODE(_3189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__B1 (.DIODE(_3189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__B (.DIODE(_3189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8005__B1 (.DIODE(_3192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8008__B1 (.DIODE(_3194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8407__B2 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8388__A1 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8365__B1 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8341__B2 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8290__A1 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8241__B1 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8211__A1 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8178__B1 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8118__B1 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8008__B2 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8053__A1 (.DIODE(_3213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8053__A2 (.DIODE(_3224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7494__B2 (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A1 (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__B1 (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__B1 (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__A1 (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__B (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__A1 (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8088__A1 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8088__A2 (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8089__B1 (.DIODE(_3282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8122__A1 (.DIODE(_3314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8150__B1 (.DIODE(_3346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8180__A1 (.DIODE(_3378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8211__A2 (.DIODE(_3411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8243__A1 (.DIODE(_3445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8267__B1 (.DIODE(_3471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8290__A2 (.DIODE(_3495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8315__B1 (.DIODE(_3523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8317__B1 (.DIODE(_3524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8341__A1_N (.DIODE(_3534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8341__A2_N (.DIODE(_3549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8367__A1 (.DIODE(_3577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8388__A2 (.DIODE(_3599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8407__A1 (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__A (.DIODE(_3615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__A (.DIODE(_3615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__B (.DIODE(_3615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A2 (.DIODE(_3615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A2 (.DIODE(_3615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__B (.DIODE(_3615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__B (.DIODE(_3615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__B (.DIODE(_3615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__A2 (.DIODE(_3615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__B1 (.DIODE(_3615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8409__A1 (.DIODE(_3621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8419__B (.DIODE(_3630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7516__A2 (.DIODE(_3635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__B (.DIODE(_3635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A3 (.DIODE(_3635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A2 (.DIODE(_3635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A2 (.DIODE(_3635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__A2 (.DIODE(_3635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__A2 (.DIODE(_3635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A2 (.DIODE(_3635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__A2 (.DIODE(_3635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__A2 (.DIODE(_3635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8477__S (.DIODE(_3654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8475__S (.DIODE(_3654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8473__S (.DIODE(_3654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8471__S (.DIODE(_3654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8469__S (.DIODE(_3654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8467__S (.DIODE(_3654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8446__A (.DIODE(_3654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8465__S (.DIODE(_3655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8463__S (.DIODE(_3655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8461__S (.DIODE(_3655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8459__S (.DIODE(_3655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8457__S (.DIODE(_3655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8455__S (.DIODE(_3655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8453__S (.DIODE(_3655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8451__S (.DIODE(_3655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8449__S (.DIODE(_3655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8447__S (.DIODE(_3655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8512__S (.DIODE(_3676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8510__S (.DIODE(_3676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8508__S (.DIODE(_3676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8506__S (.DIODE(_3676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8504__S (.DIODE(_3676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8502__S (.DIODE(_3676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8481__A (.DIODE(_3676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A (.DIODE(_3690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A1 (.DIODE(_3690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__B1 (.DIODE(_3690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A1 (.DIODE(_3690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__B2 (.DIODE(_3690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__A (.DIODE(_3690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__A1 (.DIODE(_3690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__B1 (.DIODE(_3690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__A1_N (.DIODE(_3690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A1 (.DIODE(_3690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6021__A1 (.DIODE(_3701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A (.DIODE(_3701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A1 (.DIODE(_3701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A (.DIODE(_3701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A (.DIODE(_3701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__B (.DIODE(_3701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A (.DIODE(_3701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__A1 (.DIODE(_3701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__A (.DIODE(_3701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__A (.DIODE(_3701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__B (.DIODE(_3702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__B1 (.DIODE(_3702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__B1 (.DIODE(_3702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__B (.DIODE(_3702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__B (.DIODE(_3702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__B (.DIODE(_3702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__B (.DIODE(_3702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__B (.DIODE(_3702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__A (.DIODE(_3702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7648__A1 (.DIODE(_3703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__A2 (.DIODE(_3703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__B (.DIODE(_3703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__B (.DIODE(_3703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__B (.DIODE(_3703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__A (.DIODE(_3703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__B (.DIODE(_3703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__B (.DIODE(_3703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A2 (.DIODE(_3703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__B (.DIODE(_3703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A (.DIODE(_3719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__A1 (.DIODE(_3719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A1 (.DIODE(_3719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A (.DIODE(_3719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A (.DIODE(_3719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A (.DIODE(_3719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__A (.DIODE(_3719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A (.DIODE(_3719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__A (.DIODE(_3719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__A (.DIODE(_3719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A0 (.DIODE(_3729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__S (.DIODE(_3729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A1 (.DIODE(_3729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__B1 (.DIODE(_3729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A (.DIODE(_3729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__B2 (.DIODE(_3729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__A (.DIODE(_3729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__A (.DIODE(_3729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__C (.DIODE(_3729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A (.DIODE(_3729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A (.DIODE(_3735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__B2 (.DIODE(_3735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__A (.DIODE(_3735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A1 (.DIODE(_3735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A (.DIODE(_3735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__C (.DIODE(_3735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__B2 (.DIODE(_3735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A (.DIODE(_3735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__A (.DIODE(_3735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__A (.DIODE(_3735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A0 (.DIODE(_3736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A1 (.DIODE(_3736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__B2 (.DIODE(_3736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__C1 (.DIODE(_3736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__C1 (.DIODE(_3736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A (.DIODE(_3736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__A1 (.DIODE(_3736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__A (.DIODE(_3736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__A (.DIODE(_3736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A (.DIODE(_3736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__A2 (.DIODE(_3739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__A2 (.DIODE(_3739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__B (.DIODE(_3739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__A (.DIODE(_3739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__A1 (.DIODE(_3739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__B (.DIODE(_3739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__A (.DIODE(_3739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__A (.DIODE(_3739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__A2 (.DIODE(_3739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B (.DIODE(_3739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__B1 (.DIODE(_3750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__B (.DIODE(_3750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__B (.DIODE(_3750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__A (.DIODE(_3750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__B (.DIODE(_3750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__B (.DIODE(_3750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__B (.DIODE(_3750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__C (.DIODE(_3750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__B1 (.DIODE(_3762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__B1 (.DIODE(_3762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__B1 (.DIODE(_3762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A (.DIODE(_3762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__A (.DIODE(_3762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__B1 (.DIODE(_3762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__A (.DIODE(_3762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__A1 (.DIODE(_3762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A1 (.DIODE(_3762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A (.DIODE(_3762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__A (.DIODE(_3763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A (.DIODE(_3763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A (.DIODE(_3763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A (.DIODE(_3763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__B2 (.DIODE(_3763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A1 (.DIODE(_3763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__B (.DIODE(_3763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A (.DIODE(_3763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__A (.DIODE(_3763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__A (.DIODE(_3763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__A1 (.DIODE(_3770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A (.DIODE(_3770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A (.DIODE(_3770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A (.DIODE(_3770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__A (.DIODE(_3770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A (.DIODE(_3770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__B (.DIODE(_3770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__A (.DIODE(_3770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__C (.DIODE(_3770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__A (.DIODE(_3770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7648__A0 (.DIODE(_3771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__C (.DIODE(_3771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__B2 (.DIODE(_3771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__A (.DIODE(_3771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__A2 (.DIODE(_3771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A2 (.DIODE(_3771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__B (.DIODE(_3771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__A1 (.DIODE(_3771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__B1 (.DIODE(_3771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__C1 (.DIODE(_3771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7624__A1 (.DIODE(_3776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__B2 (.DIODE(_3776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__A1 (.DIODE(_3776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A (.DIODE(_3776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__B (.DIODE(_3776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__A (.DIODE(_3776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__B2 (.DIODE(_3776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__A (.DIODE(_3776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__B (.DIODE(_3776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__C (.DIODE(_3776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A (.DIODE(_3792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__A (.DIODE(_3792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A (.DIODE(_3792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__A1 (.DIODE(_3792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A (.DIODE(_3792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__B1 (.DIODE(_3792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A (.DIODE(_3792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__B2 (.DIODE(_3792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__A1 (.DIODE(_3792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__A (.DIODE(_3792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7630__A0 (.DIODE(_3793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A2 (.DIODE(_3793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__B2 (.DIODE(_3793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A1 (.DIODE(_3793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A1 (.DIODE(_3793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__A (.DIODE(_3793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__A (.DIODE(_3793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__A (.DIODE(_3793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__B2 (.DIODE(_3793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__A (.DIODE(_3793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7630__A1 (.DIODE(_3795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__A (.DIODE(_3795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__C (.DIODE(_3795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__B (.DIODE(_3795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A2 (.DIODE(_3795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__B (.DIODE(_3795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__A2 (.DIODE(_3795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__B (.DIODE(_3795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__B (.DIODE(_3795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__B (.DIODE(_3795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A (.DIODE(_3800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A1 (.DIODE(_3800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A (.DIODE(_3800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A1 (.DIODE(_3800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A1 (.DIODE(_3800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__A (.DIODE(_3800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__B (.DIODE(_3800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A1 (.DIODE(_3800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__A (.DIODE(_3800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A1 (.DIODE(_3800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7577__A0 (.DIODE(_3802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7571__A1 (.DIODE(_3802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__A (.DIODE(_3802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__B1 (.DIODE(_3802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A (.DIODE(_3802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A1 (.DIODE(_3802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__A (.DIODE(_3802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A (.DIODE(_3802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A1 (.DIODE(_3802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__A (.DIODE(_3802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7418__A2 (.DIODE(_3804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7415__B2 (.DIODE(_3804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7325__A (.DIODE(_3804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7132__A (.DIODE(_3804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__B (.DIODE(_3804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6930__C (.DIODE(_3804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A2 (.DIODE(_3804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__B1 (.DIODE(_3804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__B (.DIODE(_3804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__A (.DIODE(_3815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__A (.DIODE(_3815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A (.DIODE(_3815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A1 (.DIODE(_3815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__B (.DIODE(_3815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A2 (.DIODE(_3815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A2 (.DIODE(_3815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__B (.DIODE(_3815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A (.DIODE(_3815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__A (.DIODE(_3815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7611__A0 (.DIODE(_3816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A1 (.DIODE(_3816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__A1 (.DIODE(_3816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A (.DIODE(_3816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A1 (.DIODE(_3816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__B (.DIODE(_3816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A (.DIODE(_3816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A (.DIODE(_3816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A (.DIODE(_3816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A (.DIODE(_3816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__A1 (.DIODE(_3817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A (.DIODE(_3817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__B (.DIODE(_3817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__B (.DIODE(_3817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__A2 (.DIODE(_3817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A2 (.DIODE(_3817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__B (.DIODE(_3817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__B (.DIODE(_3817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__B (.DIODE(_3817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__B (.DIODE(_3817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A1 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A1 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__A (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__A1 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__A (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__B (.DIODE(_3828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A (.DIODE(_3828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__A (.DIODE(_3828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__B2 (.DIODE(_3828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__A (.DIODE(_3828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__B2 (.DIODE(_3828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A1 (.DIODE(_3828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__A (.DIODE(_3828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__B2 (.DIODE(_3828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__B (.DIODE(_3828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7516__B1 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__A (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__A (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A2 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__C1 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A2 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A2 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__S (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__B (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__B (.DIODE(_3832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__A2_N (.DIODE(_3832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__B1 (.DIODE(_3832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__D (.DIODE(_3832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__B1 (.DIODE(_3832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A1 (.DIODE(_3832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__B (.DIODE(_3832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__B (.DIODE(_3832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__A (.DIODE(_3832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__A (.DIODE(_3832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__B (.DIODE(_3838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__B (.DIODE(_3838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__C (.DIODE(_3838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A2 (.DIODE(_3838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__B (.DIODE(_3838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__B (.DIODE(_3838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__A (.DIODE(_3838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__C (.DIODE(_3838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__B (.DIODE(_3838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__B (.DIODE(_3838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__A (.DIODE(_3840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__B (.DIODE(_3840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A (.DIODE(_3840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A2 (.DIODE(_3840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A2 (.DIODE(_3840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__B (.DIODE(_3840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__B (.DIODE(_3840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__A2 (.DIODE(_3840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__B1 (.DIODE(_3840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__A (.DIODE(_3853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__B (.DIODE(_3853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7571__A0 (.DIODE(_3855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__A2 (.DIODE(_3855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A (.DIODE(_3855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A2 (.DIODE(_3855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A (.DIODE(_3855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__C (.DIODE(_3855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__B (.DIODE(_3855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__B (.DIODE(_3855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__B2 (.DIODE(_3866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A1 (.DIODE(_3866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A (.DIODE(_3866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A1 (.DIODE(_3866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__C1 (.DIODE(_3866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__C1 (.DIODE(_3866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__A (.DIODE(_3866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__A1 (.DIODE(_3866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__A (.DIODE(_3866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__A (.DIODE(_3866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7638__A1 (.DIODE(_3868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7633__A0 (.DIODE(_3868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__A (.DIODE(_3868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A2 (.DIODE(_3868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__D (.DIODE(_3868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__B1 (.DIODE(_3868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__B (.DIODE(_3868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__B (.DIODE(_3868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__B (.DIODE(_3868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7640__A1 (.DIODE(_3878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A1 (.DIODE(_3878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A2 (.DIODE(_3878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A1 (.DIODE(_3878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__B (.DIODE(_3878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A1 (.DIODE(_3878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__A (.DIODE(_3878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__A3 (.DIODE(_3878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__A (.DIODE(_3878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__A (.DIODE(_3878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7604__A0 (.DIODE(_3881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7597__A1 (.DIODE(_3881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A (.DIODE(_3881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__A1 (.DIODE(_3881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__A (.DIODE(_3881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__A (.DIODE(_3881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A (.DIODE(_3881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A1 (.DIODE(_3881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__A1 (.DIODE(_3881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__A (.DIODE(_3881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7624__A0 (.DIODE(_3883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__A2 (.DIODE(_3883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__B (.DIODE(_3883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A2 (.DIODE(_3883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__A (.DIODE(_3883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__B (.DIODE(_3883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A2 (.DIODE(_3883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__B (.DIODE(_3883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__A1 (.DIODE(_3892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__A (.DIODE(_3892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A1 (.DIODE(_3892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__A (.DIODE(_3892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__B2 (.DIODE(_3892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A2 (.DIODE(_3892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__A (.DIODE(_3892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A (.DIODE(_3892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__A (.DIODE(_3892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7638__A0 (.DIODE(_3893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7633__A1 (.DIODE(_3893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A (.DIODE(_3893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__A (.DIODE(_3893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A (.DIODE(_3893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__B2 (.DIODE(_3893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__A1 (.DIODE(_3893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__A (.DIODE(_3893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__A (.DIODE(_3893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A (.DIODE(_3893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7606__A1 (.DIODE(_3901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__A1 (.DIODE(_3901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A (.DIODE(_3901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__A2 (.DIODE(_3901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__A1 (.DIODE(_3901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A (.DIODE(_3901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A2 (.DIODE(_3901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A (.DIODE(_3901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__A (.DIODE(_3901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__A (.DIODE(_3901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A (.DIODE(_3924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A (.DIODE(_3924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A (.DIODE(_3924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__C1 (.DIODE(_3924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__C1 (.DIODE(_3924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__C1 (.DIODE(_3924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__S (.DIODE(_3924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A (.DIODE(_3924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__A (.DIODE(_3924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__A (.DIODE(_3924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7682__A0 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__A (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A1 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A1 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__B (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__A (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__A (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__B (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__A (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__B (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__B (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__C (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__B (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__B1 (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__A2 (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__B (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__B (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7606__A0 (.DIODE(_3986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7354__A1 (.DIODE(_3986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__A (.DIODE(_3986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6933__B (.DIODE(_3986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__A (.DIODE(_3986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__C (.DIODE(_3986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__B (.DIODE(_3986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__B (.DIODE(_3986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__B (.DIODE(_3986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__B (.DIODE(_3986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__A (.DIODE(_3988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__B (.DIODE(_3988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A (.DIODE(_3988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A1 (.DIODE(_3988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A1 (.DIODE(_3988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A2 (.DIODE(_3988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__B (.DIODE(_3988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A (.DIODE(_3988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A2 (.DIODE(_3988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A2 (.DIODE(_3988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7211__B (.DIODE(_3989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__B1 (.DIODE(_3989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__B (.DIODE(_3989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__B (.DIODE(_3989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A (.DIODE(_3989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__B1 (.DIODE(_3989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__B1 (.DIODE(_3989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__B1 (.DIODE(_4016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__B1 (.DIODE(_4016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__C1 (.DIODE(_4016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__A (.DIODE(_4016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__A (.DIODE(_4016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__A (.DIODE(_4016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A (.DIODE(_4016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__A (.DIODE(_4016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__A (.DIODE(_4016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__B1 (.DIODE(_4017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__A (.DIODE(_4017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__A (.DIODE(_4017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6009__A (.DIODE(_4017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A (.DIODE(_4017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__A (.DIODE(_4017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A (.DIODE(_4017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A (.DIODE(_4017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A1 (.DIODE(_4017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__A (.DIODE(_4017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__A (.DIODE(_4018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A (.DIODE(_4018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__B1 (.DIODE(_4033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__A (.DIODE(_4033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__A (.DIODE(_4037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__A (.DIODE(_4037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__A (.DIODE(_4037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__B (.DIODE(_4037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__B (.DIODE(_4037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A2 (.DIODE(_4037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__B (.DIODE(_4037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__B (.DIODE(_4037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A2 (.DIODE(_4037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__B (.DIODE(_4037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7620__A0 (.DIODE(_4045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7614__A1 (.DIODE(_4045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__A1 (.DIODE(_4045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__A (.DIODE(_4045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A (.DIODE(_4045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A1 (.DIODE(_4045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A1 (.DIODE(_4045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A (.DIODE(_4045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__A (.DIODE(_4045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__A (.DIODE(_4045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7339__A1 (.DIODE(_4089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__B (.DIODE(_4089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__A1 (.DIODE(_4089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7090__A1 (.DIODE(_4089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__A (.DIODE(_4089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__A (.DIODE(_4089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__B (.DIODE(_4089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__C (.DIODE(_4089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__C (.DIODE(_4089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__B (.DIODE(_4089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7650__A1 (.DIODE(_4126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__C (.DIODE(_4126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__A (.DIODE(_4126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__B (.DIODE(_4126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__A2 (.DIODE(_4126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6899__B (.DIODE(_4126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__B (.DIODE(_4126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__B (.DIODE(_4126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A (.DIODE(_4126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__B (.DIODE(_4126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7593__A1 (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7587__A0 (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7376__A1 (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7023__A (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__B (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__A (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__A (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__C (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A2 (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__B (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A (.DIODE(_4157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__A2 (.DIODE(_4157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__A (.DIODE(_4157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A1 (.DIODE(_4157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A (.DIODE(_4157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A (.DIODE(_4174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__D (.DIODE(_4174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__A (.DIODE(_4210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__A (.DIODE(_4210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__B (.DIODE(_4210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A (.DIODE(_4210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A (.DIODE(_4210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A (.DIODE(_4210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__A (.DIODE(_4210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A (.DIODE(_4210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A (.DIODE(_4210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A (.DIODE(_4210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7577__A1 (.DIODE(_4217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7381__A1 (.DIODE(_4217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__A (.DIODE(_4217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__A (.DIODE(_4217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__A1 (.DIODE(_4217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__A1 (.DIODE(_4217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__A (.DIODE(_4217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__A (.DIODE(_4217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__B (.DIODE(_4217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__B (.DIODE(_4217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7570__A1 (.DIODE(_4222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__A1 (.DIODE(_4222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__C1 (.DIODE(_4222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A1 (.DIODE(_4222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__A1 (.DIODE(_4222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__A1 (.DIODE(_4222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A (.DIODE(_4222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A1 (.DIODE(_4222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A1 (.DIODE(_4222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A (.DIODE(_4222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__B1 (.DIODE(_4228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__A (.DIODE(_4228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__A (.DIODE(_4228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A (.DIODE(_4228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A (.DIODE(_4228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__A (.DIODE(_4228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A (.DIODE(_4228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A (.DIODE(_4228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A (.DIODE(_4228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A (.DIODE(_4228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__A (.DIODE(_4232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__B (.DIODE(_4232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__A (.DIODE(_4232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__A (.DIODE(_4232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__B (.DIODE(_4232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__A2 (.DIODE(_4232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A (.DIODE(_4232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__B (.DIODE(_4232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A2 (.DIODE(_4232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__B (.DIODE(_4232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8413__B (.DIODE(_4250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7999__B (.DIODE(_4250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7687__A1 (.DIODE(_4250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7211__A (.DIODE(_4250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7170__A (.DIODE(_4250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__A (.DIODE(_4250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__A (.DIODE(_4250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A1 (.DIODE(_4250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__B (.DIODE(_4250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A (.DIODE(_4250_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8414__A1 (.DIODE(\cmd[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8412__B (.DIODE(\cmd[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8411__B (.DIODE(\cmd[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8108__B (.DIODE(\cmd[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8022__A_N (.DIODE(\cmd[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8002__B (.DIODE(\cmd[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7484__A (.DIODE(\cmd[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__C_N (.DIODE(\cmd[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__A1 (.DIODE(\cmd[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8414__B2 (.DIODE(\cmd[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8412__A (.DIODE(\cmd[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8411__A (.DIODE(\cmd[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8108__A (.DIODE(\cmd[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8022__C (.DIODE(\cmd[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8002__A (.DIODE(\cmd[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7484__C_N (.DIODE(\cmd[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__B (.DIODE(\cmd[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__A1 (.DIODE(\cmd[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8512__A1 (.DIODE(\in_reg[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8477__A0 (.DIODE(\in_reg[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A1 (.DIODE(\in_reg[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8484__A1 (.DIODE(\in_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8449__A0 (.DIODE(\in_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8427__A1 (.DIODE(\in_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__A0 (.DIODE(\in_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A1 (.DIODE(\in_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A (.DIODE(\in_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8486__A1 (.DIODE(\in_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8451__A0 (.DIODE(\in_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__A0 (.DIODE(\in_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__A1 (.DIODE(\in_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__D (.DIODE(\in_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8488__A1 (.DIODE(\in_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8453__A0 (.DIODE(\in_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__A0 (.DIODE(\in_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__A1 (.DIODE(\in_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__C (.DIODE(\in_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8494__A1 (.DIODE(\in_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8459__A0 (.DIODE(\in_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__A0 (.DIODE(\in_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__A1 (.DIODE(\in_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__A0 (.DIODE(\in_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__D (.DIODE(\in_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8496__A1 (.DIODE(\in_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8461__A0 (.DIODE(\in_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__A0 (.DIODE(\in_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__A1 (.DIODE(\in_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__A0 (.DIODE(\in_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__C (.DIODE(\in_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__8421__A1 (.DIODE(io_out[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__8467__A1 (.DIODE(\posit_add.in1[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__A1 (.DIODE(\posit_add.in1[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__B (.DIODE(\posit_add.in1[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__A (.DIODE(\posit_add.in1[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A2 (.DIODE(\posit_add.in1[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8469__A1 (.DIODE(\posit_add.in1[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__A (.DIODE(\posit_add.in1[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__A (.DIODE(\posit_add.in1[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A1 (.DIODE(\posit_add.in1[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8473__A1 (.DIODE(\posit_add.in1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__A (.DIODE(\posit_add.in1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__A (.DIODE(\posit_add.in1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8475__A1 (.DIODE(\posit_add.in1[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__A (.DIODE(\posit_add.in1[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__A (.DIODE(\posit_add.in1[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__A (.DIODE(\posit_add.in1[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8449__A1 (.DIODE(\posit_add.in1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7493__A1 (.DIODE(\posit_add.in1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__A (.DIODE(\posit_add.in1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__B_N (.DIODE(\posit_add.in1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__A2 (.DIODE(\posit_add.in1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__C (.DIODE(\posit_add.in1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__A3 (.DIODE(\posit_add.in1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__D (.DIODE(\posit_add.in1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8461__A1 (.DIODE(\posit_add.in1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7490__A (.DIODE(\posit_add.in1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__A (.DIODE(\posit_add.in1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__A (.DIODE(\posit_add.in1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__C (.DIODE(\posit_add.in1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8463__A1 (.DIODE(\posit_add.in1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__A (.DIODE(\posit_add.in1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A1 (.DIODE(\posit_add.in1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__A (.DIODE(\posit_add.in1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__B (.DIODE(\posit_add.in1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8465__A1 (.DIODE(\posit_add.in1[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__A (.DIODE(\posit_add.in1[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__A (.DIODE(\posit_add.in1[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8482__A0 (.DIODE(\posit_add.in2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__A (.DIODE(\posit_add.in2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__A (.DIODE(\posit_add.in2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__C1 (.DIODE(\posit_add.in2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__A (.DIODE(\posit_add.in2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__A (.DIODE(\posit_add.in2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__A (.DIODE(\posit_add.in2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__A (.DIODE(\posit_add.in2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__A (.DIODE(\posit_add.in2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8502__A0 (.DIODE(\posit_add.in2[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__A (.DIODE(\posit_add.in2[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__C (.DIODE(\posit_add.in2[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__D (.DIODE(\posit_add.in2[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8508__A0 (.DIODE(\posit_add.in2[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__A (.DIODE(\posit_add.in2[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__A (.DIODE(\posit_add.in2[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA__8479__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__8444__D_N (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__8479__A_N (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__8444__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__A (.DIODE(net4));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_729 ();
 assign io_out[0] = net5;
 assign io_out[1] = net6;
 assign io_out[2] = net7;
endmodule

