magic
tech sky130B
magscale 1 2
timestamp 1682098650
<< viali >>
rect 3065 27421 3099 27455
rect 3249 27421 3283 27455
rect 6653 27421 6687 27455
rect 9597 27421 9631 27455
rect 13093 27421 13127 27455
rect 17049 27421 17083 27455
rect 20637 27421 20671 27455
rect 22201 27421 22235 27455
rect 24685 27421 24719 27455
rect 27721 27421 27755 27455
rect 10149 27353 10183 27387
rect 13645 27353 13679 27387
rect 28089 27353 28123 27387
rect 3157 27285 3191 27319
rect 6929 27285 6963 27319
rect 16957 27285 16991 27319
rect 20913 27285 20947 27319
rect 22109 27285 22143 27319
rect 24961 27285 24995 27319
rect 4537 27013 4571 27047
rect 16957 27013 16991 27047
rect 28181 27013 28215 27047
rect 2605 26945 2639 26979
rect 2872 26945 2906 26979
rect 5089 26945 5123 26979
rect 7297 26945 7331 26979
rect 7849 26945 7883 26979
rect 10425 26945 10459 26979
rect 11897 26945 11931 26979
rect 19809 26945 19843 26979
rect 19993 26945 20027 26979
rect 22201 26945 22235 26979
rect 23029 26945 23063 26979
rect 25789 26945 25823 26979
rect 27353 26945 27387 26979
rect 27905 26945 27939 26979
rect 8769 26877 8803 26911
rect 9597 26877 9631 26911
rect 12541 26877 12575 26911
rect 12817 26877 12851 26911
rect 20361 26877 20395 26911
rect 22937 26877 22971 26911
rect 26065 26877 26099 26911
rect 26617 26877 26651 26911
rect 17233 26809 17267 26843
rect 3985 26741 4019 26775
rect 7205 26741 7239 26775
rect 7941 26741 7975 26775
rect 10517 26741 10551 26775
rect 11805 26741 11839 26775
rect 14289 26741 14323 26775
rect 22109 26741 22143 26775
rect 23397 26741 23431 26775
rect 27261 26741 27295 26775
rect 4169 26537 4203 26571
rect 13001 26537 13035 26571
rect 17693 26537 17727 26571
rect 23489 26537 23523 26571
rect 27721 26537 27755 26571
rect 4813 26469 4847 26503
rect 3433 26401 3467 26435
rect 6561 26401 6595 26435
rect 8033 26401 8067 26435
rect 10517 26401 10551 26435
rect 10793 26401 10827 26435
rect 15301 26401 15335 26435
rect 21741 26401 21775 26435
rect 22017 26401 22051 26435
rect 26249 26401 26283 26435
rect 5089 26333 5123 26367
rect 6285 26333 6319 26367
rect 9597 26333 9631 26367
rect 13093 26333 13127 26367
rect 14381 26333 14415 26367
rect 16313 26333 16347 26367
rect 18153 26333 18187 26367
rect 21281 26333 21315 26367
rect 25329 26333 25363 26367
rect 25421 26333 25455 26367
rect 25973 26333 26007 26367
rect 3166 26265 3200 26299
rect 3985 26265 4019 26299
rect 4201 26265 4235 26299
rect 4813 26265 4847 26299
rect 16580 26265 16614 26299
rect 21005 26265 21039 26299
rect 2053 26197 2087 26231
rect 4353 26197 4387 26231
rect 4997 26197 5031 26231
rect 9505 26197 9539 26231
rect 12265 26197 12299 26231
rect 18245 26197 18279 26231
rect 19533 26197 19567 26231
rect 2605 25993 2639 26027
rect 4445 25993 4479 26027
rect 4905 25993 4939 26027
rect 10149 25993 10183 26027
rect 12265 25993 12299 26027
rect 17325 25993 17359 26027
rect 20269 25993 20303 26027
rect 20913 25993 20947 26027
rect 23121 25993 23155 26027
rect 23949 25993 23983 26027
rect 3332 25925 3366 25959
rect 7665 25925 7699 25959
rect 8677 25925 8711 25959
rect 13553 25925 13587 25959
rect 14381 25925 14415 25959
rect 18797 25925 18831 25959
rect 2145 25857 2179 25891
rect 2421 25857 2455 25891
rect 4905 25857 4939 25891
rect 4997 25857 5031 25891
rect 8401 25857 8435 25891
rect 12173 25857 12207 25891
rect 13645 25857 13679 25891
rect 19717 25857 19751 25891
rect 20177 25857 20211 25891
rect 21005 25857 21039 25891
rect 22477 25857 22511 25891
rect 25789 25857 25823 25891
rect 27169 25857 27203 25891
rect 3065 25789 3099 25823
rect 5181 25789 5215 25823
rect 6837 25789 6871 25823
rect 14105 25789 14139 25823
rect 19073 25789 19107 25823
rect 19625 25789 19659 25823
rect 22201 25789 22235 25823
rect 24041 25789 24075 25823
rect 24133 25789 24167 25823
rect 26065 25789 26099 25823
rect 26525 25789 26559 25823
rect 2237 25653 2271 25687
rect 15853 25653 15887 25687
rect 23581 25653 23615 25687
rect 27261 25653 27295 25687
rect 3341 25449 3375 25483
rect 5273 25449 5307 25483
rect 6193 25449 6227 25483
rect 13645 25449 13679 25483
rect 22661 25449 22695 25483
rect 8125 25381 8159 25415
rect 9229 25313 9263 25347
rect 9689 25313 9723 25347
rect 11805 25313 11839 25347
rect 15393 25313 15427 25347
rect 18337 25313 18371 25347
rect 23581 25313 23615 25347
rect 23673 25313 23707 25347
rect 24685 25313 24719 25347
rect 25145 25313 25179 25347
rect 26065 25313 26099 25347
rect 27537 25313 27571 25347
rect 3157 25245 3191 25279
rect 3433 25245 3467 25279
rect 4169 25245 4203 25279
rect 4261 25245 4295 25279
rect 4997 25245 5031 25279
rect 6285 25245 6319 25279
rect 6745 25245 6779 25279
rect 9321 25245 9355 25279
rect 10885 25245 10919 25279
rect 13553 25245 13587 25279
rect 14381 25245 14415 25279
rect 17785 25245 17819 25279
rect 17877 25245 17911 25279
rect 21281 25245 21315 25279
rect 24777 25245 24811 25279
rect 27813 25245 27847 25279
rect 4537 25177 4571 25211
rect 5089 25177 5123 25211
rect 5273 25177 5307 25211
rect 7012 25177 7046 25211
rect 21548 25177 21582 25211
rect 2973 25109 3007 25143
rect 3985 25109 4019 25143
rect 4353 25109 4387 25143
rect 23121 25109 23155 25143
rect 23489 25109 23523 25143
rect 4261 24905 4295 24939
rect 7481 24905 7515 24939
rect 7941 24905 7975 24939
rect 12081 24905 12115 24939
rect 24225 24905 24259 24939
rect 7849 24837 7883 24871
rect 3137 24769 3171 24803
rect 10793 24769 10827 24803
rect 14657 24769 14691 24803
rect 17132 24769 17166 24803
rect 18889 24769 18923 24803
rect 23112 24769 23146 24803
rect 24869 24769 24903 24803
rect 24961 24769 24995 24803
rect 25145 24769 25179 24803
rect 26157 24769 26191 24803
rect 2881 24701 2915 24735
rect 8033 24701 8067 24735
rect 10885 24701 10919 24735
rect 12173 24701 12207 24735
rect 12357 24701 12391 24735
rect 14749 24701 14783 24735
rect 16865 24701 16899 24735
rect 18797 24701 18831 24735
rect 22845 24701 22879 24735
rect 26065 24701 26099 24735
rect 11161 24633 11195 24667
rect 11713 24565 11747 24599
rect 14289 24565 14323 24599
rect 18245 24565 18279 24599
rect 19257 24565 19291 24599
rect 24685 24565 24719 24599
rect 25053 24565 25087 24599
rect 3985 24361 4019 24395
rect 11805 24361 11839 24395
rect 12725 24361 12759 24395
rect 15669 24361 15703 24395
rect 17049 24361 17083 24395
rect 17509 24225 17543 24259
rect 17693 24225 17727 24259
rect 22569 24225 22603 24259
rect 2881 24157 2915 24191
rect 3065 24157 3099 24191
rect 3985 24157 4019 24191
rect 4169 24157 4203 24191
rect 6377 24157 6411 24191
rect 10425 24157 10459 24191
rect 10692 24157 10726 24191
rect 12449 24157 12483 24191
rect 12541 24157 12575 24191
rect 14289 24157 14323 24191
rect 18521 24157 18555 24191
rect 19625 24157 19659 24191
rect 22385 24157 22419 24191
rect 27905 24157 27939 24191
rect 12725 24089 12759 24123
rect 14534 24089 14568 24123
rect 17417 24089 17451 24123
rect 28181 24089 28215 24123
rect 2973 24021 3007 24055
rect 6469 24021 6503 24055
rect 12265 24021 12299 24055
rect 18613 24021 18647 24055
rect 19533 24021 19567 24055
rect 22017 24021 22051 24055
rect 22477 24021 22511 24055
rect 2881 23817 2915 23851
rect 8309 23817 8343 23851
rect 23397 23817 23431 23851
rect 6837 23749 6871 23783
rect 18889 23749 18923 23783
rect 22284 23749 22318 23783
rect 4353 23681 4387 23715
rect 15117 23681 15151 23715
rect 18613 23681 18647 23715
rect 22017 23681 22051 23715
rect 26433 23681 26467 23715
rect 27445 23681 27479 23715
rect 6561 23613 6595 23647
rect 14565 23613 14599 23647
rect 20637 23613 20671 23647
rect 27353 23613 27387 23647
rect 28181 23613 28215 23647
rect 26525 23477 26559 23511
rect 3341 23273 3375 23307
rect 11161 23273 11195 23307
rect 14289 23273 14323 23307
rect 25145 23273 25179 23307
rect 28181 23273 28215 23307
rect 23489 23205 23523 23239
rect 2421 23137 2455 23171
rect 7297 23137 7331 23171
rect 8125 23137 8159 23171
rect 8401 23137 8435 23171
rect 10701 23137 10735 23171
rect 14749 23137 14783 23171
rect 14841 23137 14875 23171
rect 23765 23137 23799 23171
rect 24685 23137 24719 23171
rect 26709 23137 26743 23171
rect 2329 23069 2363 23103
rect 2513 23069 2547 23103
rect 3157 23069 3191 23103
rect 3433 23069 3467 23103
rect 3985 23069 4019 23103
rect 6285 23069 6319 23103
rect 8033 23069 8067 23103
rect 10793 23069 10827 23103
rect 12265 23069 12299 23103
rect 12449 23069 12483 23103
rect 15669 23069 15703 23103
rect 23857 23069 23891 23103
rect 24777 23069 24811 23103
rect 26433 23069 26467 23103
rect 20821 23001 20855 23035
rect 22569 23001 22603 23035
rect 2973 22933 3007 22967
rect 5273 22933 5307 22967
rect 12265 22933 12299 22967
rect 14657 22933 14691 22967
rect 15577 22933 15611 22967
rect 4277 22729 4311 22763
rect 5365 22729 5399 22763
rect 8493 22729 8527 22763
rect 19441 22729 19475 22763
rect 23949 22729 23983 22763
rect 26525 22729 26559 22763
rect 4077 22661 4111 22695
rect 11989 22661 12023 22695
rect 12081 22661 12115 22695
rect 2504 22593 2538 22627
rect 5457 22593 5491 22627
rect 7113 22593 7147 22627
rect 7380 22593 7414 22627
rect 9413 22593 9447 22627
rect 9680 22593 9714 22627
rect 11851 22593 11885 22627
rect 12264 22593 12298 22627
rect 12357 22593 12391 22627
rect 13645 22593 13679 22627
rect 16221 22593 16255 22627
rect 17877 22593 17911 22627
rect 19809 22593 19843 22627
rect 20085 22593 20119 22627
rect 22661 22593 22695 22627
rect 26617 22593 26651 22627
rect 27353 22593 27387 22627
rect 2237 22525 2271 22559
rect 13369 22525 13403 22559
rect 14197 22525 14231 22559
rect 15945 22525 15979 22559
rect 17969 22525 18003 22559
rect 18061 22525 18095 22559
rect 4445 22457 4479 22491
rect 3617 22389 3651 22423
rect 4261 22389 4295 22423
rect 10793 22389 10827 22423
rect 11713 22389 11747 22423
rect 17509 22389 17543 22423
rect 27261 22389 27295 22423
rect 3433 22185 3467 22219
rect 7665 22185 7699 22219
rect 18613 22185 18647 22219
rect 24041 22185 24075 22219
rect 26512 22185 26546 22219
rect 4353 22049 4387 22083
rect 8125 22049 8159 22083
rect 8309 22049 8343 22083
rect 12449 22049 12483 22083
rect 15301 22049 15335 22083
rect 19533 22049 19567 22083
rect 19993 22049 20027 22083
rect 27997 22049 28031 22083
rect 2053 21981 2087 22015
rect 2320 21981 2354 22015
rect 3985 21981 4019 22015
rect 4169 21981 4203 22015
rect 5641 21981 5675 22015
rect 12633 21981 12667 22015
rect 12817 21981 12851 22015
rect 13277 21981 13311 22015
rect 14381 21981 14415 22015
rect 17233 21981 17267 22015
rect 17500 21981 17534 22015
rect 19625 21981 19659 22015
rect 22661 21981 22695 22015
rect 26249 21981 26283 22015
rect 6377 21913 6411 21947
rect 10241 21913 10275 21947
rect 11989 21913 12023 21947
rect 13553 21913 13587 21947
rect 22928 21913 22962 21947
rect 8033 21845 8067 21879
rect 3709 21641 3743 21675
rect 9781 21641 9815 21675
rect 11161 21641 11195 21675
rect 13737 21641 13771 21675
rect 15393 21641 15427 21675
rect 23213 21641 23247 21675
rect 23673 21641 23707 21675
rect 26341 21641 26375 21675
rect 28273 21641 28307 21675
rect 23581 21573 23615 21607
rect 2145 21505 2179 21539
rect 2329 21505 2363 21539
rect 2973 21505 3007 21539
rect 3893 21505 3927 21539
rect 4169 21505 4203 21539
rect 6745 21505 6779 21539
rect 10149 21505 10183 21539
rect 10241 21505 10275 21539
rect 10977 21505 11011 21539
rect 11161 21505 11195 21539
rect 12624 21505 12658 21539
rect 14657 21505 14691 21539
rect 15301 21505 15335 21539
rect 16957 21505 16991 21539
rect 17224 21505 17258 21539
rect 19257 21505 19291 21539
rect 22017 21505 22051 21539
rect 22201 21505 22235 21539
rect 24777 21505 24811 21539
rect 26433 21505 26467 21539
rect 27445 21505 27479 21539
rect 2237 21437 2271 21471
rect 3249 21437 3283 21471
rect 4077 21437 4111 21471
rect 10425 21437 10459 21471
rect 12357 21437 12391 21471
rect 14749 21437 14783 21471
rect 19165 21437 19199 21471
rect 23857 21437 23891 21471
rect 24685 21437 24719 21471
rect 27353 21437 27387 21471
rect 18337 21369 18371 21403
rect 2789 21301 2823 21335
rect 3157 21301 3191 21335
rect 6653 21301 6687 21335
rect 14289 21301 14323 21335
rect 19625 21301 19659 21335
rect 22109 21301 22143 21335
rect 24409 21301 24443 21335
rect 7113 21097 7147 21131
rect 13001 21097 13035 21131
rect 17325 21097 17359 21131
rect 23581 21097 23615 21131
rect 24041 21029 24075 21063
rect 5365 20961 5399 20995
rect 7941 20961 7975 20995
rect 8401 20961 8435 20995
rect 12173 20961 12207 20995
rect 13461 20961 13495 20995
rect 13645 20961 13679 20995
rect 14841 20961 14875 20995
rect 17877 20961 17911 20995
rect 23673 20961 23707 20995
rect 25053 20961 25087 20995
rect 3341 20893 3375 20927
rect 8033 20893 8067 20927
rect 17693 20893 17727 20927
rect 17785 20893 17819 20927
rect 19993 20893 20027 20927
rect 21833 20893 21867 20927
rect 21926 20893 21960 20927
rect 22109 20893 22143 20927
rect 22298 20893 22332 20927
rect 23581 20893 23615 20927
rect 23857 20893 23891 20927
rect 24593 20893 24627 20927
rect 24869 20893 24903 20927
rect 27905 20893 27939 20927
rect 5641 20825 5675 20859
rect 10425 20825 10459 20859
rect 14657 20825 14691 20859
rect 20260 20825 20294 20859
rect 22201 20825 22235 20859
rect 28181 20825 28215 20859
rect 2053 20757 2087 20791
rect 13369 20757 13403 20791
rect 14289 20757 14323 20791
rect 14749 20757 14783 20791
rect 21373 20757 21407 20791
rect 22477 20757 22511 20791
rect 24869 20757 24903 20791
rect 3433 20553 3467 20587
rect 5825 20553 5859 20587
rect 8217 20553 8251 20587
rect 11069 20553 11103 20587
rect 15117 20553 15151 20587
rect 20453 20553 20487 20587
rect 22385 20553 22419 20587
rect 2320 20485 2354 20519
rect 9597 20485 9631 20519
rect 14004 20485 14038 20519
rect 17132 20485 17166 20519
rect 20821 20485 20855 20519
rect 20913 20485 20947 20519
rect 22017 20485 22051 20519
rect 22201 20485 22235 20519
rect 23397 20485 23431 20519
rect 4353 20417 4387 20451
rect 4813 20417 4847 20451
rect 4997 20417 5031 20451
rect 5917 20417 5951 20451
rect 9873 20417 9907 20451
rect 10701 20417 10735 20451
rect 10885 20417 10919 20451
rect 11713 20417 11747 20451
rect 11989 20417 12023 20451
rect 12173 20417 12207 20451
rect 12817 20417 12851 20451
rect 27353 20417 27387 20451
rect 2053 20349 2087 20383
rect 4169 20349 4203 20383
rect 8309 20349 8343 20383
rect 8493 20349 8527 20383
rect 9781 20349 9815 20383
rect 12357 20349 12391 20383
rect 13093 20349 13127 20383
rect 13737 20349 13771 20383
rect 16865 20349 16899 20383
rect 21005 20349 21039 20383
rect 25145 20349 25179 20383
rect 10057 20281 10091 20315
rect 18245 20281 18279 20315
rect 5181 20213 5215 20247
rect 7849 20213 7883 20247
rect 9689 20213 9723 20247
rect 27261 20213 27295 20247
rect 8493 20009 8527 20043
rect 9689 20009 9723 20043
rect 10517 20009 10551 20043
rect 17693 20009 17727 20043
rect 20085 20009 20119 20043
rect 21281 20009 21315 20043
rect 28273 20009 28307 20043
rect 24041 19941 24075 19975
rect 9413 19873 9447 19907
rect 11897 19873 11931 19907
rect 13185 19873 13219 19907
rect 14565 19873 14599 19907
rect 16773 19873 16807 19907
rect 22661 19873 22695 19907
rect 25053 19873 25087 19907
rect 25145 19873 25179 19907
rect 26801 19873 26835 19907
rect 2053 19805 2087 19839
rect 3985 19805 4019 19839
rect 6745 19805 6779 19839
rect 9321 19805 9355 19839
rect 13001 19805 13035 19839
rect 13553 19805 13587 19839
rect 16589 19805 16623 19839
rect 16957 19805 16991 19839
rect 17601 19805 17635 19839
rect 17785 19805 17819 19839
rect 24961 19805 24995 19839
rect 25881 19805 25915 19839
rect 25973 19805 26007 19839
rect 26525 19805 26559 19839
rect 2320 19737 2354 19771
rect 7021 19737 7055 19771
rect 11630 19737 11664 19771
rect 15393 19737 15427 19771
rect 19809 19737 19843 19771
rect 20913 19737 20947 19771
rect 21097 19737 21131 19771
rect 22928 19737 22962 19771
rect 3433 19669 3467 19703
rect 5181 19669 5215 19703
rect 24593 19669 24627 19703
rect 5917 19465 5951 19499
rect 6653 19465 6687 19499
rect 8585 19465 8619 19499
rect 9505 19465 9539 19499
rect 11713 19465 11747 19499
rect 16221 19465 16255 19499
rect 16865 19465 16899 19499
rect 21097 19465 21131 19499
rect 22201 19465 22235 19499
rect 28273 19465 28307 19499
rect 4353 19397 4387 19431
rect 7472 19397 7506 19431
rect 12173 19397 12207 19431
rect 2973 19329 3007 19363
rect 4905 19329 4939 19363
rect 5089 19329 5123 19363
rect 5181 19329 5215 19363
rect 6009 19329 6043 19363
rect 6561 19329 6595 19363
rect 9597 19329 9631 19363
rect 10333 19329 10367 19363
rect 12081 19329 12115 19363
rect 13093 19329 13127 19363
rect 13277 19329 13311 19363
rect 13921 19329 13955 19363
rect 14197 19329 14231 19363
rect 16037 19329 16071 19363
rect 17049 19329 17083 19363
rect 19717 19329 19751 19363
rect 19984 19329 20018 19363
rect 22017 19329 22051 19363
rect 22201 19329 22235 19363
rect 22661 19329 22695 19363
rect 22928 19329 22962 19363
rect 24961 19329 24995 19363
rect 26157 19329 26191 19363
rect 27445 19329 27479 19363
rect 2789 19261 2823 19295
rect 3157 19261 3191 19295
rect 3249 19261 3283 19295
rect 7205 19261 7239 19295
rect 9689 19261 9723 19295
rect 12265 19261 12299 19295
rect 12909 19261 12943 19295
rect 14289 19261 14323 19295
rect 15853 19261 15887 19295
rect 17233 19261 17267 19295
rect 24593 19261 24627 19295
rect 24869 19261 24903 19295
rect 27353 19261 27387 19295
rect 4905 19193 4939 19227
rect 10517 19193 10551 19227
rect 24041 19193 24075 19227
rect 4077 19125 4111 19159
rect 9137 19125 9171 19159
rect 26065 19125 26099 19159
rect 10517 18921 10551 18955
rect 13001 18921 13035 18955
rect 21281 18921 21315 18955
rect 22937 18921 22971 18955
rect 27445 18921 27479 18955
rect 16037 18853 16071 18887
rect 17233 18853 17267 18887
rect 5917 18785 5951 18819
rect 6745 18785 6779 18819
rect 13444 18785 13478 18819
rect 21741 18785 21775 18819
rect 21833 18785 21867 18819
rect 23489 18785 23523 18819
rect 25973 18785 26007 18819
rect 3985 18717 4019 18751
rect 4169 18717 4203 18751
rect 9137 18717 9171 18751
rect 9393 18717 9427 18751
rect 13645 18717 13679 18751
rect 13737 18717 13771 18751
rect 15945 18717 15979 18751
rect 16129 18717 16163 18751
rect 16773 18717 16807 18751
rect 16957 18717 16991 18751
rect 17325 18717 17359 18751
rect 18245 18717 18279 18751
rect 18521 18717 18555 18751
rect 19901 18717 19935 18751
rect 20821 18717 20855 18751
rect 23397 18717 23431 18751
rect 24961 18717 24995 18751
rect 25053 18717 25087 18751
rect 25697 18717 25731 18751
rect 4353 18649 4387 18683
rect 13185 18649 13219 18683
rect 13553 18581 13587 18615
rect 18889 18581 18923 18615
rect 21649 18581 21683 18615
rect 23305 18581 23339 18615
rect 4905 18377 4939 18411
rect 14841 18377 14875 18411
rect 17417 18377 17451 18411
rect 20453 18377 20487 18411
rect 26617 18377 26651 18411
rect 2881 18309 2915 18343
rect 7849 18309 7883 18343
rect 9597 18309 9631 18343
rect 17233 18309 17267 18343
rect 4813 18241 4847 18275
rect 6745 18241 6779 18275
rect 13093 18241 13127 18275
rect 13553 18241 13587 18275
rect 13921 18241 13955 18275
rect 14933 18241 14967 18275
rect 24961 18241 24995 18275
rect 25789 18241 25823 18275
rect 26249 18241 26283 18275
rect 2605 18173 2639 18207
rect 4353 18173 4387 18207
rect 14105 18173 14139 18207
rect 18705 18173 18739 18207
rect 18981 18173 19015 18207
rect 13553 18105 13587 18139
rect 16865 18105 16899 18139
rect 6653 18037 6687 18071
rect 17233 18037 17267 18071
rect 24869 18037 24903 18071
rect 2881 17833 2915 17867
rect 4077 17833 4111 17867
rect 9689 17833 9723 17867
rect 19901 17833 19935 17867
rect 9413 17697 9447 17731
rect 11805 17697 11839 17731
rect 15577 17697 15611 17731
rect 22753 17697 22787 17731
rect 2973 17629 3007 17663
rect 4169 17629 4203 17663
rect 5549 17629 5583 17663
rect 6193 17629 6227 17663
rect 9321 17629 9355 17663
rect 14565 17629 14599 17663
rect 19993 17629 20027 17663
rect 24593 17629 24627 17663
rect 24860 17629 24894 17663
rect 27905 17629 27939 17663
rect 7205 17561 7239 17595
rect 12072 17561 12106 17595
rect 14289 17561 14323 17595
rect 14657 17561 14691 17595
rect 15025 17561 15059 17595
rect 15844 17561 15878 17595
rect 22477 17561 22511 17595
rect 28181 17561 28215 17595
rect 5457 17493 5491 17527
rect 13185 17493 13219 17527
rect 14473 17493 14507 17527
rect 16957 17493 16991 17527
rect 22109 17493 22143 17527
rect 22569 17493 22603 17527
rect 25973 17493 26007 17527
rect 16957 17289 16991 17323
rect 27629 17289 27663 17323
rect 13921 17221 13955 17255
rect 14473 17221 14507 17255
rect 22293 17221 22327 17255
rect 24041 17221 24075 17255
rect 26249 17221 26283 17255
rect 27261 17221 27295 17255
rect 2789 17153 2823 17187
rect 4445 17153 4479 17187
rect 5917 17153 5951 17187
rect 7297 17153 7331 17187
rect 11713 17153 11747 17187
rect 11969 17153 12003 17187
rect 13829 17153 13863 17187
rect 14013 17153 14047 17187
rect 15025 17153 15059 17187
rect 15209 17153 15243 17187
rect 17057 17151 17091 17185
rect 24501 17153 24535 17187
rect 24685 17153 24719 17187
rect 24961 17153 24995 17187
rect 25329 17153 25363 17187
rect 26157 17153 26191 17187
rect 26341 17153 26375 17187
rect 27169 17153 27203 17187
rect 27445 17153 27479 17187
rect 4997 17085 5031 17119
rect 14381 17085 14415 17119
rect 15393 17085 15427 17119
rect 22017 17085 22051 17119
rect 24869 17085 24903 17119
rect 2697 16949 2731 16983
rect 4353 16949 4387 16983
rect 9505 16949 9539 16983
rect 13093 16949 13127 16983
rect 8309 16745 8343 16779
rect 12357 16745 12391 16779
rect 16221 16745 16255 16779
rect 25237 16745 25271 16779
rect 27629 16745 27663 16779
rect 24041 16677 24075 16711
rect 24685 16677 24719 16711
rect 6561 16609 6595 16643
rect 6837 16609 6871 16643
rect 9137 16609 9171 16643
rect 11713 16609 11747 16643
rect 11897 16609 11931 16643
rect 13645 16609 13679 16643
rect 14657 16609 14691 16643
rect 18245 16609 18279 16643
rect 18429 16609 18463 16643
rect 22293 16609 22327 16643
rect 27169 16609 27203 16643
rect 2513 16541 2547 16575
rect 3341 16541 3375 16575
rect 13001 16541 13035 16575
rect 13185 16541 13219 16575
rect 14289 16541 14323 16575
rect 14749 16541 14783 16575
rect 16129 16541 16163 16575
rect 16681 16541 16715 16575
rect 24869 16541 24903 16575
rect 25053 16541 25087 16575
rect 27261 16541 27295 16575
rect 9382 16473 9416 16507
rect 13093 16473 13127 16507
rect 13553 16473 13587 16507
rect 18521 16473 18555 16507
rect 22569 16473 22603 16507
rect 24961 16473 24995 16507
rect 2421 16405 2455 16439
rect 3249 16405 3283 16439
rect 10517 16405 10551 16439
rect 11989 16405 12023 16439
rect 18889 16405 18923 16439
rect 9137 16201 9171 16235
rect 9597 16201 9631 16235
rect 11713 16201 11747 16235
rect 12173 16201 12207 16235
rect 13461 16201 13495 16235
rect 22569 16201 22603 16235
rect 23029 16201 23063 16235
rect 23489 16201 23523 16235
rect 2329 16133 2363 16167
rect 4077 16133 4111 16167
rect 9505 16133 9539 16167
rect 15945 16133 15979 16167
rect 19594 16133 19628 16167
rect 2053 16065 2087 16099
rect 10701 16065 10735 16099
rect 12081 16065 12115 16099
rect 14749 16065 14783 16099
rect 17776 16065 17810 16099
rect 19349 16065 19383 16099
rect 22385 16065 22419 16099
rect 22569 16065 22603 16099
rect 23397 16065 23431 16099
rect 6561 15997 6595 16031
rect 7389 15997 7423 16031
rect 9689 15997 9723 16031
rect 10977 15997 11011 16031
rect 12265 15997 12299 16031
rect 15761 15997 15795 16031
rect 15853 15997 15887 16031
rect 17509 15997 17543 16031
rect 23673 15997 23707 16031
rect 20729 15929 20763 15963
rect 11069 15861 11103 15895
rect 16313 15861 16347 15895
rect 18889 15861 18923 15895
rect 7297 15657 7331 15691
rect 17877 15657 17911 15691
rect 22845 15657 22879 15691
rect 11345 15521 11379 15555
rect 12449 15521 12483 15555
rect 20361 15521 20395 15555
rect 20637 15521 20671 15555
rect 1961 15453 1995 15487
rect 2605 15453 2639 15487
rect 3341 15453 3375 15487
rect 5549 15453 5583 15487
rect 9689 15453 9723 15487
rect 14289 15453 14323 15487
rect 16497 15453 16531 15487
rect 16753 15453 16787 15487
rect 20269 15453 20303 15487
rect 22753 15453 22787 15487
rect 22937 15453 22971 15487
rect 26157 15453 26191 15487
rect 5825 15385 5859 15419
rect 9965 15385 9999 15419
rect 12633 15385 12667 15419
rect 12817 15385 12851 15419
rect 13185 15385 13219 15419
rect 1869 15317 1903 15351
rect 2513 15317 2547 15351
rect 3249 15317 3283 15351
rect 10793 15317 10827 15351
rect 11161 15317 11195 15351
rect 11253 15317 11287 15351
rect 12725 15317 12759 15351
rect 15577 15317 15611 15351
rect 26065 15317 26099 15351
rect 17877 15113 17911 15147
rect 18245 15113 18279 15147
rect 24961 15113 24995 15147
rect 2237 15045 2271 15079
rect 14933 15045 14967 15079
rect 1961 14977 1995 15011
rect 5089 14977 5123 15011
rect 6561 14977 6595 15011
rect 7481 14977 7515 15011
rect 9956 14977 9990 15011
rect 13369 14977 13403 15011
rect 13461 14977 13495 15011
rect 13921 14977 13955 15011
rect 15025 14977 15059 15011
rect 15117 14977 15151 15011
rect 15577 14977 15611 15011
rect 18337 14977 18371 15011
rect 19257 14977 19291 15011
rect 20729 14977 20763 15011
rect 21373 14977 21407 15011
rect 24861 14977 24895 15011
rect 27353 14977 27387 15011
rect 3985 14909 4019 14943
rect 4813 14909 4847 14943
rect 9689 14909 9723 14943
rect 13645 14909 13679 14943
rect 15485 14909 15519 14943
rect 18429 14909 18463 14943
rect 19165 14909 19199 14943
rect 25789 14909 25823 14943
rect 26525 14909 26559 14943
rect 14289 14841 14323 14875
rect 6653 14773 6687 14807
rect 7573 14773 7607 14807
rect 11069 14773 11103 14807
rect 19625 14773 19659 14807
rect 20637 14773 20671 14807
rect 21281 14773 21315 14807
rect 27261 14773 27295 14807
rect 11621 14569 11655 14603
rect 12449 14569 12483 14603
rect 27445 14569 27479 14603
rect 10517 14433 10551 14467
rect 13001 14433 13035 14467
rect 13737 14433 13771 14467
rect 20361 14433 20395 14467
rect 20637 14433 20671 14467
rect 22385 14433 22419 14467
rect 25697 14433 25731 14467
rect 25973 14433 26007 14467
rect 2145 14365 2179 14399
rect 2789 14365 2823 14399
rect 3433 14365 3467 14399
rect 5181 14365 5215 14399
rect 5641 14365 5675 14399
rect 8309 14365 8343 14399
rect 10241 14365 10275 14399
rect 12357 14365 12391 14399
rect 14473 14365 14507 14399
rect 14749 14365 14783 14399
rect 14841 14365 14875 14399
rect 15485 14365 15519 14399
rect 15669 14365 15703 14399
rect 5917 14297 5951 14331
rect 7665 14297 7699 14331
rect 13185 14297 13219 14331
rect 13369 14297 13403 14331
rect 14657 14297 14691 14331
rect 15853 14297 15887 14331
rect 2053 14229 2087 14263
rect 2697 14229 2731 14263
rect 3341 14229 3375 14263
rect 5089 14229 5123 14263
rect 8217 14229 8251 14263
rect 13277 14229 13311 14263
rect 15025 14229 15059 14263
rect 5549 14025 5583 14059
rect 6653 14025 6687 14059
rect 9689 14025 9723 14059
rect 10425 14025 10459 14059
rect 10885 14025 10919 14059
rect 14749 14025 14783 14059
rect 2329 13957 2363 13991
rect 8217 13957 8251 13991
rect 15761 13957 15795 13991
rect 16054 13957 16088 13991
rect 21189 13957 21223 13991
rect 27997 13957 28031 13991
rect 4813 13889 4847 13923
rect 5457 13889 5491 13923
rect 6745 13889 6779 13923
rect 7941 13889 7975 13923
rect 10793 13889 10827 13923
rect 12173 13889 12207 13923
rect 12909 13889 12943 13923
rect 13636 13889 13670 13923
rect 15485 13889 15519 13923
rect 15669 13889 15703 13923
rect 15905 13889 15939 13923
rect 17325 13889 17359 13923
rect 17509 13889 17543 13923
rect 18153 13889 18187 13923
rect 18337 13889 18371 13923
rect 22845 13889 22879 13923
rect 23112 13889 23146 13923
rect 26433 13889 26467 13923
rect 2053 13821 2087 13855
rect 4077 13821 4111 13855
rect 4905 13821 4939 13855
rect 10977 13821 11011 13855
rect 12541 13821 12575 13855
rect 13369 13821 13403 13855
rect 17693 13821 17727 13855
rect 20637 13821 20671 13855
rect 27445 13821 27479 13855
rect 18245 13685 18279 13719
rect 24225 13685 24259 13719
rect 26341 13685 26375 13719
rect 2329 13481 2363 13515
rect 10885 13481 10919 13515
rect 23121 13481 23155 13515
rect 27997 13481 28031 13515
rect 9873 13413 9907 13447
rect 4077 13345 4111 13379
rect 5825 13345 5859 13379
rect 6101 13345 6135 13379
rect 12633 13345 12667 13379
rect 23581 13345 23615 13379
rect 23765 13345 23799 13379
rect 24593 13345 24627 13379
rect 24869 13345 24903 13379
rect 26249 13345 26283 13379
rect 26525 13345 26559 13379
rect 1777 13277 1811 13311
rect 2421 13277 2455 13311
rect 3065 13277 3099 13311
rect 6561 13277 6595 13311
rect 9781 13277 9815 13311
rect 10977 13277 11011 13311
rect 11713 13277 11747 13311
rect 12173 13277 12207 13311
rect 12725 13277 12759 13311
rect 13001 13277 13035 13311
rect 14657 13277 14691 13311
rect 14933 13277 14967 13311
rect 15761 13277 15795 13311
rect 17601 13277 17635 13311
rect 17694 13277 17728 13311
rect 17969 13277 18003 13311
rect 18107 13277 18141 13311
rect 19533 13277 19567 13311
rect 19717 13277 19751 13311
rect 19901 13277 19935 13311
rect 23489 13277 23523 13311
rect 24961 13277 24995 13311
rect 6806 13209 6840 13243
rect 12081 13209 12115 13243
rect 14565 13209 14599 13243
rect 16028 13209 16062 13243
rect 17877 13209 17911 13243
rect 22293 13209 22327 13243
rect 1685 13141 1719 13175
rect 2973 13141 3007 13175
rect 7941 13141 7975 13175
rect 11989 13141 12023 13175
rect 17141 13141 17175 13175
rect 18245 13141 18279 13175
rect 19533 13141 19567 13175
rect 22385 13141 22419 13175
rect 6561 12937 6595 12971
rect 7021 12937 7055 12971
rect 13461 12937 13495 12971
rect 16865 12937 16899 12971
rect 17325 12937 17359 12971
rect 21005 12937 21039 12971
rect 1869 12869 1903 12903
rect 3617 12869 3651 12903
rect 14749 12869 14783 12903
rect 15393 12869 15427 12903
rect 15761 12869 15795 12903
rect 21465 12869 21499 12903
rect 28181 12869 28215 12903
rect 1593 12801 1627 12835
rect 4629 12801 4663 12835
rect 5273 12801 5307 12835
rect 6929 12801 6963 12835
rect 9617 12801 9651 12835
rect 10885 12801 10919 12835
rect 12541 12801 12575 12835
rect 15577 12801 15611 12835
rect 17233 12801 17267 12835
rect 18889 12801 18923 12835
rect 19156 12801 19190 12835
rect 21189 12801 21223 12835
rect 22293 12801 22327 12835
rect 22560 12801 22594 12835
rect 26341 12801 26375 12835
rect 27353 12801 27387 12835
rect 27905 12801 27939 12835
rect 7205 12733 7239 12767
rect 9873 12733 9907 12767
rect 12357 12733 12391 12767
rect 17509 12733 17543 12767
rect 21281 12733 21315 12767
rect 5181 12597 5215 12631
rect 8493 12597 8527 12631
rect 10793 12597 10827 12631
rect 20269 12597 20303 12631
rect 21189 12597 21223 12631
rect 23673 12597 23707 12631
rect 26433 12597 26467 12631
rect 27261 12597 27295 12631
rect 9873 12393 9907 12427
rect 14289 12393 14323 12427
rect 15577 12393 15611 12427
rect 17233 12393 17267 12427
rect 19441 12393 19475 12427
rect 21189 12393 21223 12427
rect 22661 12393 22695 12427
rect 28181 12393 28215 12427
rect 5733 12257 5767 12291
rect 9321 12257 9355 12291
rect 10977 12257 11011 12291
rect 14841 12257 14875 12291
rect 16957 12257 16991 12291
rect 19901 12257 19935 12291
rect 19993 12257 20027 12291
rect 20729 12257 20763 12291
rect 23305 12257 23339 12291
rect 26433 12257 26467 12291
rect 26709 12257 26743 12291
rect 4077 12189 4111 12223
rect 9413 12189 9447 12223
rect 11253 12189 11287 12223
rect 11989 12189 12023 12223
rect 12817 12189 12851 12223
rect 14657 12189 14691 12223
rect 14749 12189 14783 12223
rect 15485 12189 15519 12223
rect 15669 12189 15703 12223
rect 16865 12189 16899 12223
rect 20821 12189 20855 12223
rect 23029 12189 23063 12223
rect 23121 12189 23155 12223
rect 25697 12189 25731 12223
rect 4629 12121 4663 12155
rect 6000 12121 6034 12155
rect 7113 12053 7147 12087
rect 9505 12053 9539 12087
rect 12081 12053 12115 12087
rect 12725 12053 12759 12087
rect 19809 12053 19843 12087
rect 25605 12053 25639 12087
rect 6561 11849 6595 11883
rect 7021 11849 7055 11883
rect 18245 11849 18279 11883
rect 26525 11849 26559 11883
rect 13737 11781 13771 11815
rect 25053 11781 25087 11815
rect 27997 11781 28031 11815
rect 3065 11713 3099 11747
rect 3249 11713 3283 11747
rect 5365 11713 5399 11747
rect 6929 11713 6963 11747
rect 10701 11713 10735 11747
rect 10977 11713 11011 11747
rect 11161 11713 11195 11747
rect 11713 11713 11747 11747
rect 15025 11713 15059 11747
rect 16865 11713 16899 11747
rect 17132 11713 17166 11747
rect 19717 11713 19751 11747
rect 23213 11713 23247 11747
rect 24041 11713 24075 11747
rect 2329 11645 2363 11679
rect 4261 11645 4295 11679
rect 7205 11645 7239 11679
rect 10793 11645 10827 11679
rect 10885 11645 10919 11679
rect 11989 11645 12023 11679
rect 14933 11645 14967 11679
rect 19809 11645 19843 11679
rect 20637 11645 20671 11679
rect 21373 11645 21407 11679
rect 22845 11645 22879 11679
rect 23305 11645 23339 11679
rect 24777 11645 24811 11679
rect 27445 11645 27479 11679
rect 10517 11509 10551 11543
rect 15393 11509 15427 11543
rect 19349 11509 19383 11543
rect 23949 11509 23983 11543
rect 10793 11305 10827 11339
rect 17141 11305 17175 11339
rect 19625 11305 19659 11339
rect 19901 11305 19935 11339
rect 24777 11305 24811 11339
rect 3341 11237 3375 11271
rect 22385 11237 22419 11271
rect 5089 11169 5123 11203
rect 6653 11169 6687 11203
rect 6929 11169 6963 11203
rect 9229 11169 9263 11203
rect 9689 11169 9723 11203
rect 14749 11169 14783 11203
rect 14933 11169 14967 11203
rect 16589 11169 16623 11203
rect 19533 11169 19567 11203
rect 25697 11169 25731 11203
rect 1593 11101 1627 11135
rect 5457 11101 5491 11135
rect 6561 11101 6595 11135
rect 7389 11101 7423 11135
rect 8309 11101 8343 11135
rect 9321 11101 9355 11135
rect 10885 11101 10919 11135
rect 11805 11101 11839 11135
rect 14657 11101 14691 11135
rect 16681 11101 16715 11135
rect 19717 11101 19751 11135
rect 20637 11101 20671 11135
rect 21097 11101 21131 11135
rect 23305 11101 23339 11135
rect 24685 11101 24719 11135
rect 26617 11101 26651 11135
rect 1869 11033 1903 11067
rect 11529 11033 11563 11067
rect 19441 11033 19475 11067
rect 7481 10965 7515 10999
rect 8217 10965 8251 10999
rect 14289 10965 14323 10999
rect 16773 10965 16807 10999
rect 20545 10965 20579 10999
rect 23397 10965 23431 10999
rect 2421 10761 2455 10795
rect 14657 10761 14691 10795
rect 24593 10761 24627 10795
rect 7389 10693 7423 10727
rect 9137 10693 9171 10727
rect 13544 10693 13578 10727
rect 19717 10693 19751 10727
rect 23121 10693 23155 10727
rect 2513 10625 2547 10659
rect 2973 10625 3007 10659
rect 7113 10625 7147 10659
rect 13277 10625 13311 10659
rect 17233 10625 17267 10659
rect 19257 10625 19291 10659
rect 22845 10625 22879 10659
rect 27905 10625 27939 10659
rect 3065 10557 3099 10591
rect 3617 10557 3651 10591
rect 3893 10557 3927 10591
rect 17325 10557 17359 10591
rect 17417 10557 17451 10591
rect 21465 10557 21499 10591
rect 28181 10557 28215 10591
rect 5365 10421 5399 10455
rect 16865 10421 16899 10455
rect 19165 10421 19199 10455
rect 2329 10217 2363 10251
rect 9965 10217 9999 10251
rect 17877 10217 17911 10251
rect 18889 10217 18923 10251
rect 22017 10217 22051 10251
rect 6377 10149 6411 10183
rect 27629 10149 27663 10183
rect 4169 10081 4203 10115
rect 4997 10081 5031 10115
rect 6101 10081 6135 10115
rect 8217 10081 8251 10115
rect 12357 10081 12391 10115
rect 18429 10081 18463 10115
rect 20269 10081 20303 10115
rect 20545 10081 20579 10115
rect 24041 10081 24075 10115
rect 27169 10081 27203 10115
rect 2421 10013 2455 10047
rect 4261 10013 4295 10047
rect 6009 10013 6043 10047
rect 7297 10013 7331 10047
rect 7481 10013 7515 10047
rect 11345 10013 11379 10047
rect 16497 10013 16531 10047
rect 16764 10013 16798 10047
rect 18521 10013 18555 10047
rect 19809 10013 19843 10047
rect 23029 10013 23063 10047
rect 27261 10013 27295 10047
rect 11100 9945 11134 9979
rect 12265 9945 12299 9979
rect 11805 9877 11839 9911
rect 12173 9877 12207 9911
rect 19717 9877 19751 9911
rect 26525 9673 26559 9707
rect 27629 9673 27663 9707
rect 4629 9605 4663 9639
rect 9689 9605 9723 9639
rect 10609 9605 10643 9639
rect 19257 9605 19291 9639
rect 2789 9537 2823 9571
rect 4721 9537 4755 9571
rect 9597 9537 9631 9571
rect 9781 9537 9815 9571
rect 10241 9537 10275 9571
rect 10334 9537 10368 9571
rect 10517 9537 10551 9571
rect 10747 9537 10781 9571
rect 14933 9537 14967 9571
rect 17509 9537 17543 9571
rect 26433 9537 26467 9571
rect 26617 9537 26651 9571
rect 18981 9469 19015 9503
rect 20729 9469 20763 9503
rect 27169 9469 27203 9503
rect 10885 9401 10919 9435
rect 27537 9401 27571 9435
rect 2697 9333 2731 9367
rect 14841 9333 14875 9367
rect 17417 9333 17451 9367
rect 10517 9129 10551 9163
rect 18797 9129 18831 9163
rect 26893 9129 26927 9163
rect 9597 9061 9631 9095
rect 27997 9061 28031 9095
rect 2697 8993 2731 9027
rect 7021 8993 7055 9027
rect 7297 8993 7331 9027
rect 11713 8993 11747 9027
rect 17785 8993 17819 9027
rect 19717 8993 19751 9027
rect 20453 8993 20487 9027
rect 23857 8993 23891 9027
rect 27905 8993 27939 9027
rect 2605 8925 2639 8959
rect 6929 8925 6963 8959
rect 9505 8925 9539 8959
rect 9689 8925 9723 8959
rect 10149 8925 10183 8959
rect 11437 8925 11471 8959
rect 14381 8925 14415 8959
rect 15945 8925 15979 8959
rect 18245 8925 18279 8959
rect 18705 8925 18739 8959
rect 22661 8925 22695 8959
rect 22845 8925 22879 8959
rect 23673 8925 23707 8959
rect 27077 8925 27111 8959
rect 27169 8925 27203 8959
rect 27261 8925 27295 8959
rect 27389 8925 27423 8959
rect 10333 8857 10367 8891
rect 15393 8857 15427 8891
rect 28365 8857 28399 8891
rect 3433 8789 3467 8823
rect 11069 8789 11103 8823
rect 11529 8789 11563 8823
rect 16037 8789 16071 8823
rect 22845 8789 22879 8823
rect 23305 8789 23339 8823
rect 23765 8789 23799 8823
rect 4077 8585 4111 8619
rect 8125 8585 8159 8619
rect 10885 8585 10919 8619
rect 15853 8585 15887 8619
rect 18613 8585 18647 8619
rect 24593 8585 24627 8619
rect 27721 8585 27755 8619
rect 2605 8517 2639 8551
rect 10517 8517 10551 8551
rect 14381 8517 14415 8551
rect 17141 8517 17175 8551
rect 23121 8517 23155 8551
rect 6745 8449 6779 8483
rect 7012 8449 7046 8483
rect 10701 8449 10735 8483
rect 11713 8449 11747 8483
rect 11897 8449 11931 8483
rect 13645 8449 13679 8483
rect 16865 8449 16899 8483
rect 22845 8449 22879 8483
rect 27353 8449 27387 8483
rect 2329 8381 2363 8415
rect 13553 8381 13587 8415
rect 14105 8381 14139 8415
rect 27445 8381 27479 8415
rect 11897 8313 11931 8347
rect 2605 8041 2639 8075
rect 5825 8041 5859 8075
rect 9321 8041 9355 8075
rect 12173 8041 12207 8075
rect 16037 8041 16071 8075
rect 26801 8041 26835 8075
rect 27813 8041 27847 8075
rect 9505 7905 9539 7939
rect 17693 7905 17727 7939
rect 20269 7905 20303 7939
rect 22201 7905 22235 7939
rect 2697 7837 2731 7871
rect 3341 7837 3375 7871
rect 8493 7837 8527 7871
rect 9321 7837 9355 7871
rect 10793 7837 10827 7871
rect 11060 7837 11094 7871
rect 13737 7837 13771 7871
rect 14289 7837 14323 7871
rect 16681 7837 16715 7871
rect 24593 7837 24627 7871
rect 24777 7837 24811 7871
rect 27261 7837 27295 7871
rect 27629 7837 27663 7871
rect 4537 7769 4571 7803
rect 6929 7769 6963 7803
rect 9597 7769 9631 7803
rect 13645 7769 13679 7803
rect 14565 7769 14599 7803
rect 20536 7769 20570 7803
rect 22477 7769 22511 7803
rect 24685 7769 24719 7803
rect 26249 7769 26283 7803
rect 26525 7769 26559 7803
rect 27445 7769 27479 7803
rect 27537 7769 27571 7803
rect 3249 7701 3283 7735
rect 9137 7701 9171 7735
rect 21649 7701 21683 7735
rect 23949 7701 23983 7735
rect 26433 7701 26467 7735
rect 26617 7701 26651 7735
rect 3893 7497 3927 7531
rect 7389 7497 7423 7531
rect 7849 7497 7883 7531
rect 10333 7497 10367 7531
rect 18705 7497 18739 7531
rect 21189 7497 21223 7531
rect 23213 7497 23247 7531
rect 23581 7497 23615 7531
rect 23673 7497 23707 7531
rect 26341 7497 26375 7531
rect 26617 7497 26651 7531
rect 27537 7497 27571 7531
rect 2421 7429 2455 7463
rect 4712 7429 4746 7463
rect 15025 7429 15059 7463
rect 19993 7429 20027 7463
rect 25329 7429 25363 7463
rect 27353 7429 27387 7463
rect 4445 7361 4479 7395
rect 7757 7361 7791 7395
rect 21281 7361 21315 7395
rect 25145 7361 25179 7395
rect 25421 7361 25455 7395
rect 25549 7367 25583 7401
rect 26249 7361 26283 7395
rect 26433 7361 26467 7395
rect 27169 7361 27203 7395
rect 27997 7361 28031 7395
rect 2145 7293 2179 7327
rect 8033 7293 8067 7327
rect 10425 7293 10459 7327
rect 10609 7293 10643 7327
rect 14197 7293 14231 7327
rect 23857 7293 23891 7327
rect 25237 7293 25271 7327
rect 26065 7225 26099 7259
rect 5825 7157 5859 7191
rect 9965 7157 9999 7191
rect 28089 7157 28123 7191
rect 4905 6953 4939 6987
rect 7665 6953 7699 6987
rect 27721 6953 27755 6987
rect 2697 6817 2731 6851
rect 3433 6817 3467 6851
rect 5549 6817 5583 6851
rect 6653 6817 6687 6851
rect 7757 6817 7791 6851
rect 10885 6817 10919 6851
rect 12817 6817 12851 6851
rect 17141 6817 17175 6851
rect 2605 6749 2639 6783
rect 5365 6749 5399 6783
rect 7665 6749 7699 6783
rect 7941 6749 7975 6783
rect 10618 6749 10652 6783
rect 16865 6749 16899 6783
rect 19441 6749 19475 6783
rect 19625 6749 19659 6783
rect 22661 6749 22695 6783
rect 22917 6749 22951 6783
rect 25697 6749 25731 6783
rect 25789 6749 25823 6783
rect 26341 6749 26375 6783
rect 26608 6749 26642 6783
rect 5273 6681 5307 6715
rect 6101 6613 6135 6647
rect 6469 6613 6503 6647
rect 6561 6613 6595 6647
rect 8125 6613 8159 6647
rect 9505 6613 9539 6647
rect 12265 6613 12299 6647
rect 12633 6613 12667 6647
rect 12725 6613 12759 6647
rect 18613 6613 18647 6647
rect 19533 6613 19567 6647
rect 24041 6613 24075 6647
rect 2605 6409 2639 6443
rect 13277 6409 13311 6443
rect 17601 6409 17635 6443
rect 24317 6409 24351 6443
rect 6653 6341 6687 6375
rect 12164 6341 12198 6375
rect 2697 6273 2731 6307
rect 3157 6273 3191 6307
rect 5089 6273 5123 6307
rect 6837 6273 6871 6307
rect 7665 6273 7699 6307
rect 10526 6273 10560 6307
rect 10793 6273 10827 6307
rect 11897 6273 11931 6307
rect 17509 6273 17543 6307
rect 17693 6273 17727 6307
rect 18521 6273 18555 6307
rect 20453 6273 20487 6307
rect 20637 6273 20671 6307
rect 23193 6273 23227 6307
rect 27905 6273 27939 6307
rect 5181 6205 5215 6239
rect 7757 6205 7791 6239
rect 8033 6205 8067 6239
rect 18153 6205 18187 6239
rect 22937 6205 22971 6239
rect 28181 6205 28215 6239
rect 5457 6137 5491 6171
rect 3249 6069 3283 6103
rect 7021 6069 7055 6103
rect 9413 6069 9447 6103
rect 19947 6069 19981 6103
rect 20545 6069 20579 6103
rect 6837 5865 6871 5899
rect 7849 5865 7883 5899
rect 9873 5865 9907 5899
rect 11805 5865 11839 5899
rect 17187 5865 17221 5899
rect 21281 5865 21315 5899
rect 5457 5729 5491 5763
rect 10517 5729 10551 5763
rect 12265 5729 12299 5763
rect 19809 5729 19843 5763
rect 2605 5661 2639 5695
rect 3065 5661 3099 5695
rect 3985 5661 4019 5695
rect 5724 5661 5758 5695
rect 7297 5661 7331 5695
rect 7665 5661 7699 5695
rect 8309 5661 8343 5695
rect 8493 5661 8527 5695
rect 10333 5661 10367 5695
rect 12173 5661 12207 5695
rect 14749 5661 14783 5695
rect 14933 5661 14967 5695
rect 15393 5661 15427 5695
rect 15761 5661 15795 5695
rect 19533 5661 19567 5695
rect 21741 5661 21775 5695
rect 21925 5661 21959 5695
rect 27813 5661 27847 5695
rect 7481 5593 7515 5627
rect 7573 5593 7607 5627
rect 10241 5593 10275 5627
rect 27546 5593 27580 5627
rect 3433 5525 3467 5559
rect 4077 5525 4111 5559
rect 8309 5525 8343 5559
rect 14933 5525 14967 5559
rect 21741 5525 21775 5559
rect 26433 5525 26467 5559
rect 2605 5321 2639 5355
rect 7389 5321 7423 5355
rect 15761 5321 15795 5355
rect 16865 5321 16899 5355
rect 26157 5321 26191 5355
rect 27261 5321 27295 5355
rect 27905 5321 27939 5355
rect 4077 5253 4111 5287
rect 6837 5253 6871 5287
rect 7757 5253 7791 5287
rect 4353 5185 4387 5219
rect 6745 5185 6779 5219
rect 6929 5185 6963 5219
rect 7573 5185 7607 5219
rect 16865 5185 16899 5219
rect 17049 5185 17083 5219
rect 22017 5185 22051 5219
rect 22201 5185 22235 5219
rect 22661 5185 22695 5219
rect 22845 5185 22879 5219
rect 26249 5185 26283 5219
rect 26341 5185 26375 5219
rect 27169 5185 27203 5219
rect 27813 5185 27847 5219
rect 14013 5117 14047 5151
rect 14289 5117 14323 5151
rect 25973 5117 26007 5151
rect 22109 4981 22143 5015
rect 22753 4981 22787 5015
rect 26249 4981 26283 5015
rect 24041 4777 24075 4811
rect 27353 4777 27387 4811
rect 27905 4777 27939 4811
rect 6469 4641 6503 4675
rect 20729 4641 20763 4675
rect 28273 4641 28307 4675
rect 4721 4573 4755 4607
rect 6745 4573 6779 4607
rect 7849 4573 7883 4607
rect 9965 4573 9999 4607
rect 10517 4573 10551 4607
rect 10701 4573 10735 4607
rect 20361 4573 20395 4607
rect 22661 4573 22695 4607
rect 25513 4573 25547 4607
rect 27077 4573 27111 4607
rect 27169 4573 27203 4607
rect 28181 4573 28215 4607
rect 22928 4505 22962 4539
rect 25789 4505 25823 4539
rect 26065 4505 26099 4539
rect 4629 4437 4663 4471
rect 7389 4437 7423 4471
rect 7941 4437 7975 4471
rect 9873 4437 9907 4471
rect 11529 4437 11563 4471
rect 22155 4437 22189 4471
rect 25697 4437 25731 4471
rect 25881 4437 25915 4471
rect 26709 4437 26743 4471
rect 11069 4233 11103 4267
rect 27721 4233 27755 4267
rect 28273 4233 28307 4267
rect 27445 4165 27479 4199
rect 3341 4097 3375 4131
rect 3801 4097 3835 4131
rect 6653 4097 6687 4131
rect 7389 4097 7423 4131
rect 7757 4097 7791 4131
rect 11713 4097 11747 4131
rect 17233 4097 17267 4131
rect 19829 4097 19863 4131
rect 23388 4097 23422 4131
rect 25605 4097 25639 4131
rect 25789 4097 25823 4131
rect 25973 4097 26007 4131
rect 26249 4097 26283 4131
rect 27169 4097 27203 4131
rect 27353 4097 27387 4131
rect 27537 4097 27571 4131
rect 28181 4097 28215 4131
rect 28365 4097 28399 4131
rect 4077 4029 4111 4063
rect 8309 4029 8343 4063
rect 9321 4029 9355 4063
rect 9597 4029 9631 4063
rect 12909 4029 12943 4063
rect 13277 4029 13311 4063
rect 14703 4029 14737 4063
rect 17141 4029 17175 4063
rect 20085 4029 20119 4063
rect 23121 4029 23155 4063
rect 3249 3961 3283 3995
rect 5549 3893 5583 3927
rect 6745 3893 6779 3927
rect 11805 3893 11839 3927
rect 16865 3893 16899 3927
rect 18705 3893 18739 3927
rect 24501 3893 24535 3927
rect 26249 3893 26283 3927
rect 10149 3689 10183 3723
rect 10793 3689 10827 3723
rect 16129 3689 16163 3723
rect 19993 3689 20027 3723
rect 22799 3689 22833 3723
rect 24685 3689 24719 3723
rect 25881 3689 25915 3723
rect 8493 3621 8527 3655
rect 4169 3553 4203 3587
rect 5089 3553 5123 3587
rect 7021 3553 7055 3587
rect 12265 3553 12299 3587
rect 16589 3553 16623 3587
rect 19533 3553 19567 3587
rect 21373 3553 21407 3587
rect 4445 3485 4479 3519
rect 6285 3485 6319 3519
rect 6745 3485 6779 3519
rect 10241 3485 10275 3519
rect 12541 3485 12575 3519
rect 14749 3485 14783 3519
rect 16856 3485 16890 3519
rect 19625 3485 19659 3519
rect 21005 3485 21039 3519
rect 24777 3485 24811 3519
rect 27261 3485 27295 3519
rect 27721 3485 27755 3519
rect 14994 3417 15028 3451
rect 27016 3417 27050 3451
rect 27813 3417 27847 3451
rect 6193 3349 6227 3383
rect 17969 3349 18003 3383
rect 10885 3145 10919 3179
rect 14013 3145 14047 3179
rect 14933 3145 14967 3179
rect 18981 3145 19015 3179
rect 23765 3145 23799 3179
rect 25697 3145 25731 3179
rect 26249 3145 26283 3179
rect 4261 3077 4295 3111
rect 8125 3077 8159 3111
rect 17868 3077 17902 3111
rect 24562 3077 24596 3111
rect 6009 3009 6043 3043
rect 8401 3009 8435 3043
rect 9873 3009 9907 3043
rect 10241 3009 10275 3043
rect 12889 3009 12923 3043
rect 16057 3009 16091 3043
rect 19809 3009 19843 3043
rect 22017 3009 22051 3043
rect 26157 3009 26191 3043
rect 27169 3009 27203 3043
rect 27353 3009 27387 3043
rect 12633 2941 12667 2975
rect 16313 2941 16347 2975
rect 17601 2941 17635 2975
rect 19441 2941 19475 2975
rect 19717 2941 19751 2975
rect 22293 2941 22327 2975
rect 24317 2941 24351 2975
rect 6653 2873 6687 2907
rect 27169 2805 27203 2839
rect 7297 2601 7331 2635
rect 12357 2601 12391 2635
rect 13737 2465 13771 2499
rect 7389 2397 7423 2431
rect 27905 2397 27939 2431
rect 13492 2329 13526 2363
rect 28181 2329 28215 2363
<< metal1 >>
rect 1104 27770 28888 27792
rect 1104 27718 4423 27770
rect 4475 27718 4487 27770
rect 4539 27718 4551 27770
rect 4603 27718 4615 27770
rect 4667 27718 4679 27770
rect 4731 27718 11369 27770
rect 11421 27718 11433 27770
rect 11485 27718 11497 27770
rect 11549 27718 11561 27770
rect 11613 27718 11625 27770
rect 11677 27718 18315 27770
rect 18367 27718 18379 27770
rect 18431 27718 18443 27770
rect 18495 27718 18507 27770
rect 18559 27718 18571 27770
rect 18623 27718 25261 27770
rect 25313 27718 25325 27770
rect 25377 27718 25389 27770
rect 25441 27718 25453 27770
rect 25505 27718 25517 27770
rect 25569 27718 28888 27770
rect 1104 27696 28888 27718
rect 17678 27480 17684 27532
rect 17736 27520 17742 27532
rect 27890 27520 27896 27532
rect 17736 27492 27896 27520
rect 17736 27480 17742 27492
rect 27890 27480 27896 27492
rect 27948 27480 27954 27532
rect 3053 27455 3111 27461
rect 3053 27421 3065 27455
rect 3099 27421 3111 27455
rect 3053 27415 3111 27421
rect 3237 27455 3295 27461
rect 3237 27421 3249 27455
rect 3283 27452 3295 27455
rect 3326 27452 3332 27464
rect 3283 27424 3332 27452
rect 3283 27421 3295 27424
rect 3237 27415 3295 27421
rect 3068 27384 3096 27415
rect 3326 27412 3332 27424
rect 3384 27412 3390 27464
rect 5718 27412 5724 27464
rect 5776 27452 5782 27464
rect 6641 27455 6699 27461
rect 6641 27452 6653 27455
rect 5776 27424 6653 27452
rect 5776 27412 5782 27424
rect 6641 27421 6653 27424
rect 6687 27421 6699 27455
rect 9582 27452 9588 27464
rect 9543 27424 9588 27452
rect 6641 27415 6699 27421
rect 9582 27412 9588 27424
rect 9640 27412 9646 27464
rect 13078 27452 13084 27464
rect 13039 27424 13084 27452
rect 13078 27412 13084 27424
rect 13136 27412 13142 27464
rect 17034 27452 17040 27464
rect 16995 27424 17040 27452
rect 17034 27412 17040 27424
rect 17092 27412 17098 27464
rect 20622 27452 20628 27464
rect 20583 27424 20628 27452
rect 20622 27412 20628 27424
rect 20680 27412 20686 27464
rect 22189 27455 22247 27461
rect 22189 27421 22201 27455
rect 22235 27452 22247 27455
rect 22278 27452 22284 27464
rect 22235 27424 22284 27452
rect 22235 27421 22247 27424
rect 22189 27415 22247 27421
rect 22278 27412 22284 27424
rect 22336 27412 22342 27464
rect 24118 27412 24124 27464
rect 24176 27452 24182 27464
rect 24673 27455 24731 27461
rect 24673 27452 24685 27455
rect 24176 27424 24685 27452
rect 24176 27412 24182 27424
rect 24673 27421 24685 27424
rect 24719 27421 24731 27455
rect 27706 27452 27712 27464
rect 27667 27424 27712 27452
rect 24673 27415 24731 27421
rect 27706 27412 27712 27424
rect 27764 27412 27770 27464
rect 4522 27384 4528 27396
rect 3068 27356 4528 27384
rect 4522 27344 4528 27356
rect 4580 27344 4586 27396
rect 10137 27387 10195 27393
rect 10137 27353 10149 27387
rect 10183 27384 10195 27387
rect 12618 27384 12624 27396
rect 10183 27356 12624 27384
rect 10183 27353 10195 27356
rect 10137 27347 10195 27353
rect 12618 27344 12624 27356
rect 12676 27344 12682 27396
rect 13633 27387 13691 27393
rect 13633 27353 13645 27387
rect 13679 27384 13691 27387
rect 13722 27384 13728 27396
rect 13679 27356 13728 27384
rect 13679 27353 13691 27356
rect 13633 27347 13691 27353
rect 13722 27344 13728 27356
rect 13780 27344 13786 27396
rect 28074 27384 28080 27396
rect 28035 27356 28080 27384
rect 28074 27344 28080 27356
rect 28132 27344 28138 27396
rect 3142 27316 3148 27328
rect 3103 27288 3148 27316
rect 3142 27276 3148 27288
rect 3200 27276 3206 27328
rect 6914 27276 6920 27328
rect 6972 27316 6978 27328
rect 16942 27316 16948 27328
rect 6972 27288 7017 27316
rect 16903 27288 16948 27316
rect 6972 27276 6978 27288
rect 16942 27276 16948 27288
rect 17000 27276 17006 27328
rect 20898 27316 20904 27328
rect 20859 27288 20904 27316
rect 20898 27276 20904 27288
rect 20956 27276 20962 27328
rect 22097 27319 22155 27325
rect 22097 27285 22109 27319
rect 22143 27316 22155 27319
rect 22186 27316 22192 27328
rect 22143 27288 22192 27316
rect 22143 27285 22155 27288
rect 22097 27279 22155 27285
rect 22186 27276 22192 27288
rect 22244 27276 22250 27328
rect 24946 27316 24952 27328
rect 24907 27288 24952 27316
rect 24946 27276 24952 27288
rect 25004 27276 25010 27328
rect 1104 27226 29048 27248
rect 1104 27174 7896 27226
rect 7948 27174 7960 27226
rect 8012 27174 8024 27226
rect 8076 27174 8088 27226
rect 8140 27174 8152 27226
rect 8204 27174 14842 27226
rect 14894 27174 14906 27226
rect 14958 27174 14970 27226
rect 15022 27174 15034 27226
rect 15086 27174 15098 27226
rect 15150 27174 21788 27226
rect 21840 27174 21852 27226
rect 21904 27174 21916 27226
rect 21968 27174 21980 27226
rect 22032 27174 22044 27226
rect 22096 27174 28734 27226
rect 28786 27174 28798 27226
rect 28850 27174 28862 27226
rect 28914 27174 28926 27226
rect 28978 27174 28990 27226
rect 29042 27174 29048 27226
rect 1104 27152 29048 27174
rect 3418 27044 3424 27056
rect 2608 27016 3424 27044
rect 2608 26985 2636 27016
rect 3418 27004 3424 27016
rect 3476 27004 3482 27056
rect 4522 27044 4528 27056
rect 4483 27016 4528 27044
rect 4522 27004 4528 27016
rect 4580 27044 4586 27056
rect 5258 27044 5264 27056
rect 4580 27016 5264 27044
rect 4580 27004 4586 27016
rect 5258 27004 5264 27016
rect 5316 27004 5322 27056
rect 16942 27044 16948 27056
rect 16903 27016 16948 27044
rect 16942 27004 16948 27016
rect 17000 27004 17006 27056
rect 22830 27044 22836 27056
rect 22204 27016 22836 27044
rect 2866 26985 2872 26988
rect 2593 26979 2651 26985
rect 2593 26945 2605 26979
rect 2639 26945 2651 26979
rect 2593 26939 2651 26945
rect 2860 26939 2872 26985
rect 2924 26976 2930 26988
rect 5077 26979 5135 26985
rect 2924 26948 2960 26976
rect 2866 26936 2872 26939
rect 2924 26936 2930 26948
rect 5077 26945 5089 26979
rect 5123 26976 5135 26979
rect 6914 26976 6920 26988
rect 5123 26948 6920 26976
rect 5123 26945 5135 26948
rect 5077 26939 5135 26945
rect 6914 26936 6920 26948
rect 6972 26936 6978 26988
rect 7285 26979 7343 26985
rect 7285 26945 7297 26979
rect 7331 26976 7343 26979
rect 7837 26979 7895 26985
rect 7837 26976 7849 26979
rect 7331 26948 7849 26976
rect 7331 26945 7343 26948
rect 7285 26939 7343 26945
rect 7837 26945 7849 26948
rect 7883 26976 7895 26979
rect 8294 26976 8300 26988
rect 7883 26948 8300 26976
rect 7883 26945 7895 26948
rect 7837 26939 7895 26945
rect 8294 26936 8300 26948
rect 8352 26936 8358 26988
rect 9490 26976 9496 26988
rect 9246 26948 9496 26976
rect 9490 26936 9496 26948
rect 9548 26936 9554 26988
rect 10410 26976 10416 26988
rect 10371 26948 10416 26976
rect 10410 26936 10416 26948
rect 10468 26936 10474 26988
rect 11885 26979 11943 26985
rect 11885 26945 11897 26979
rect 11931 26976 11943 26979
rect 12250 26976 12256 26988
rect 11931 26948 12256 26976
rect 11931 26945 11943 26948
rect 11885 26939 11943 26945
rect 12250 26936 12256 26948
rect 12308 26936 12314 26988
rect 15286 26976 15292 26988
rect 13938 26948 15292 26976
rect 15286 26936 15292 26948
rect 15344 26936 15350 26988
rect 19794 26976 19800 26988
rect 19755 26948 19800 26976
rect 19794 26936 19800 26948
rect 19852 26936 19858 26988
rect 19978 26976 19984 26988
rect 19939 26948 19984 26976
rect 19978 26936 19984 26948
rect 20036 26936 20042 26988
rect 22204 26985 22232 27016
rect 22830 27004 22836 27016
rect 22888 27044 22894 27056
rect 22888 27016 26234 27044
rect 22888 27004 22894 27016
rect 22189 26979 22247 26985
rect 22189 26945 22201 26979
rect 22235 26945 22247 26979
rect 22189 26939 22247 26945
rect 22278 26936 22284 26988
rect 22336 26976 22342 26988
rect 23014 26976 23020 26988
rect 22336 26948 23020 26976
rect 22336 26936 22342 26948
rect 23014 26936 23020 26948
rect 23072 26936 23078 26988
rect 25774 26976 25780 26988
rect 25735 26948 25780 26976
rect 25774 26936 25780 26948
rect 25832 26936 25838 26988
rect 26206 26976 26234 27016
rect 27522 27004 27528 27056
rect 27580 27044 27586 27056
rect 28169 27047 28227 27053
rect 28169 27044 28181 27047
rect 27580 27016 28181 27044
rect 27580 27004 27586 27016
rect 28169 27013 28181 27016
rect 28215 27013 28227 27047
rect 28169 27007 28227 27013
rect 27341 26979 27399 26985
rect 27341 26976 27353 26979
rect 26206 26948 27353 26976
rect 27341 26945 27353 26948
rect 27387 26976 27399 26979
rect 27706 26976 27712 26988
rect 27387 26948 27712 26976
rect 27387 26945 27399 26948
rect 27341 26939 27399 26945
rect 27706 26936 27712 26948
rect 27764 26936 27770 26988
rect 27890 26976 27896 26988
rect 27851 26948 27896 26976
rect 27890 26936 27896 26948
rect 27948 26936 27954 26988
rect 8754 26908 8760 26920
rect 8715 26880 8760 26908
rect 8754 26868 8760 26880
rect 8812 26868 8818 26920
rect 9585 26911 9643 26917
rect 9585 26877 9597 26911
rect 9631 26908 9643 26911
rect 9674 26908 9680 26920
rect 9631 26880 9680 26908
rect 9631 26877 9643 26880
rect 9585 26871 9643 26877
rect 9674 26868 9680 26880
rect 9732 26868 9738 26920
rect 12526 26908 12532 26920
rect 12487 26880 12532 26908
rect 12526 26868 12532 26880
rect 12584 26868 12590 26920
rect 12802 26908 12808 26920
rect 12763 26880 12808 26908
rect 12802 26868 12808 26880
rect 12860 26868 12866 26920
rect 20346 26908 20352 26920
rect 20307 26880 20352 26908
rect 20346 26868 20352 26880
rect 20404 26868 20410 26920
rect 20898 26868 20904 26920
rect 20956 26908 20962 26920
rect 22922 26908 22928 26920
rect 20956 26880 22508 26908
rect 22883 26880 22928 26908
rect 20956 26868 20962 26880
rect 16758 26800 16764 26852
rect 16816 26840 16822 26852
rect 17221 26843 17279 26849
rect 17221 26840 17233 26843
rect 16816 26812 17233 26840
rect 16816 26800 16822 26812
rect 17221 26809 17233 26812
rect 17267 26840 17279 26843
rect 22370 26840 22376 26852
rect 17267 26812 22376 26840
rect 17267 26809 17279 26812
rect 17221 26803 17279 26809
rect 22370 26800 22376 26812
rect 22428 26800 22434 26852
rect 22480 26840 22508 26880
rect 22922 26868 22928 26880
rect 22980 26868 22986 26920
rect 26050 26908 26056 26920
rect 26011 26880 26056 26908
rect 26050 26868 26056 26880
rect 26108 26868 26114 26920
rect 26605 26911 26663 26917
rect 26605 26877 26617 26911
rect 26651 26908 26663 26911
rect 26694 26908 26700 26920
rect 26651 26880 26700 26908
rect 26651 26877 26663 26880
rect 26605 26871 26663 26877
rect 26694 26868 26700 26880
rect 26752 26868 26758 26920
rect 23934 26840 23940 26852
rect 22480 26812 23940 26840
rect 23934 26800 23940 26812
rect 23992 26800 23998 26852
rect 3973 26775 4031 26781
rect 3973 26741 3985 26775
rect 4019 26772 4031 26775
rect 4154 26772 4160 26784
rect 4019 26744 4160 26772
rect 4019 26741 4031 26744
rect 3973 26735 4031 26741
rect 4154 26732 4160 26744
rect 4212 26732 4218 26784
rect 6546 26732 6552 26784
rect 6604 26772 6610 26784
rect 7193 26775 7251 26781
rect 7193 26772 7205 26775
rect 6604 26744 7205 26772
rect 6604 26732 6610 26744
rect 7193 26741 7205 26744
rect 7239 26741 7251 26775
rect 7193 26735 7251 26741
rect 7929 26775 7987 26781
rect 7929 26741 7941 26775
rect 7975 26772 7987 26775
rect 8386 26772 8392 26784
rect 7975 26744 8392 26772
rect 7975 26741 7987 26744
rect 7929 26735 7987 26741
rect 8386 26732 8392 26744
rect 8444 26732 8450 26784
rect 10502 26772 10508 26784
rect 10463 26744 10508 26772
rect 10502 26732 10508 26744
rect 10560 26732 10566 26784
rect 10778 26732 10784 26784
rect 10836 26772 10842 26784
rect 11793 26775 11851 26781
rect 11793 26772 11805 26775
rect 10836 26744 11805 26772
rect 10836 26732 10842 26744
rect 11793 26741 11805 26744
rect 11839 26741 11851 26775
rect 11793 26735 11851 26741
rect 13170 26732 13176 26784
rect 13228 26772 13234 26784
rect 14277 26775 14335 26781
rect 14277 26772 14289 26775
rect 13228 26744 14289 26772
rect 13228 26732 13234 26744
rect 14277 26741 14289 26744
rect 14323 26741 14335 26775
rect 14277 26735 14335 26741
rect 21726 26732 21732 26784
rect 21784 26772 21790 26784
rect 22097 26775 22155 26781
rect 22097 26772 22109 26775
rect 21784 26744 22109 26772
rect 21784 26732 21790 26744
rect 22097 26741 22109 26744
rect 22143 26741 22155 26775
rect 23382 26772 23388 26784
rect 23343 26744 23388 26772
rect 22097 26735 22155 26741
rect 23382 26732 23388 26744
rect 23440 26732 23446 26784
rect 27246 26772 27252 26784
rect 27207 26744 27252 26772
rect 27246 26732 27252 26744
rect 27304 26732 27310 26784
rect 1104 26682 28888 26704
rect 1104 26630 4423 26682
rect 4475 26630 4487 26682
rect 4539 26630 4551 26682
rect 4603 26630 4615 26682
rect 4667 26630 4679 26682
rect 4731 26630 11369 26682
rect 11421 26630 11433 26682
rect 11485 26630 11497 26682
rect 11549 26630 11561 26682
rect 11613 26630 11625 26682
rect 11677 26630 18315 26682
rect 18367 26630 18379 26682
rect 18431 26630 18443 26682
rect 18495 26630 18507 26682
rect 18559 26630 18571 26682
rect 18623 26630 25261 26682
rect 25313 26630 25325 26682
rect 25377 26630 25389 26682
rect 25441 26630 25453 26682
rect 25505 26630 25517 26682
rect 25569 26630 28888 26682
rect 1104 26608 28888 26630
rect 4154 26568 4160 26580
rect 4115 26540 4160 26568
rect 4154 26528 4160 26540
rect 4212 26528 4218 26580
rect 8754 26528 8760 26580
rect 8812 26568 8818 26580
rect 9858 26568 9864 26580
rect 8812 26540 9864 26568
rect 8812 26528 8818 26540
rect 9858 26528 9864 26540
rect 9916 26568 9922 26580
rect 9916 26540 11836 26568
rect 9916 26528 9922 26540
rect 4801 26503 4859 26509
rect 4801 26469 4813 26503
rect 4847 26500 4859 26503
rect 4982 26500 4988 26512
rect 4847 26472 4988 26500
rect 4847 26469 4859 26472
rect 4801 26463 4859 26469
rect 4982 26460 4988 26472
rect 5040 26460 5046 26512
rect 3418 26432 3424 26444
rect 3379 26404 3424 26432
rect 3418 26392 3424 26404
rect 3476 26392 3482 26444
rect 6546 26432 6552 26444
rect 6507 26404 6552 26432
rect 6546 26392 6552 26404
rect 6604 26392 6610 26444
rect 8021 26435 8079 26441
rect 8021 26401 8033 26435
rect 8067 26432 8079 26435
rect 8294 26432 8300 26444
rect 8067 26404 8300 26432
rect 8067 26401 8079 26404
rect 8021 26395 8079 26401
rect 8294 26392 8300 26404
rect 8352 26432 8358 26444
rect 9306 26432 9312 26444
rect 8352 26404 9312 26432
rect 8352 26392 8358 26404
rect 9306 26392 9312 26404
rect 9364 26392 9370 26444
rect 10502 26432 10508 26444
rect 10463 26404 10508 26432
rect 10502 26392 10508 26404
rect 10560 26392 10566 26444
rect 10778 26432 10784 26444
rect 10739 26404 10784 26432
rect 10778 26392 10784 26404
rect 10836 26392 10842 26444
rect 11808 26432 11836 26540
rect 12802 26528 12808 26580
rect 12860 26568 12866 26580
rect 12989 26571 13047 26577
rect 12989 26568 13001 26571
rect 12860 26540 13001 26568
rect 12860 26528 12866 26540
rect 12989 26537 13001 26540
rect 13035 26537 13047 26571
rect 17678 26568 17684 26580
rect 17639 26540 17684 26568
rect 12989 26531 13047 26537
rect 17678 26528 17684 26540
rect 17736 26528 17742 26580
rect 19794 26528 19800 26580
rect 19852 26568 19858 26580
rect 22462 26568 22468 26580
rect 19852 26540 22468 26568
rect 19852 26528 19858 26540
rect 22462 26528 22468 26540
rect 22520 26528 22526 26580
rect 23014 26528 23020 26580
rect 23072 26568 23078 26580
rect 23477 26571 23535 26577
rect 23477 26568 23489 26571
rect 23072 26540 23489 26568
rect 23072 26528 23078 26540
rect 23477 26537 23489 26540
rect 23523 26537 23535 26571
rect 27706 26568 27712 26580
rect 27667 26540 27712 26568
rect 23477 26531 23535 26537
rect 27706 26528 27712 26540
rect 27764 26528 27770 26580
rect 15286 26432 15292 26444
rect 11808 26404 14412 26432
rect 15247 26404 15292 26432
rect 2866 26324 2872 26376
rect 2924 26364 2930 26376
rect 3436 26364 3464 26392
rect 14384 26376 14412 26404
rect 15286 26392 15292 26404
rect 15344 26392 15350 26444
rect 21726 26432 21732 26444
rect 21687 26404 21732 26432
rect 21726 26392 21732 26404
rect 21784 26392 21790 26444
rect 22005 26435 22063 26441
rect 22005 26401 22017 26435
rect 22051 26432 22063 26435
rect 22094 26432 22100 26444
rect 22051 26404 22100 26432
rect 22051 26401 22063 26404
rect 22005 26395 22063 26401
rect 22094 26392 22100 26404
rect 22152 26392 22158 26444
rect 26237 26435 26295 26441
rect 26237 26401 26249 26435
rect 26283 26432 26295 26435
rect 27246 26432 27252 26444
rect 26283 26404 27252 26432
rect 26283 26401 26295 26404
rect 26237 26395 26295 26401
rect 27246 26392 27252 26404
rect 27304 26392 27310 26444
rect 5074 26364 5080 26376
rect 2924 26336 3464 26364
rect 3988 26336 4936 26364
rect 5035 26336 5080 26364
rect 2924 26324 2930 26336
rect 3142 26256 3148 26308
rect 3200 26305 3206 26308
rect 3200 26296 3212 26305
rect 3200 26268 3245 26296
rect 3200 26259 3212 26268
rect 3200 26256 3206 26259
rect 3326 26256 3332 26308
rect 3384 26296 3390 26308
rect 3988 26305 4016 26336
rect 3973 26299 4031 26305
rect 3973 26296 3985 26299
rect 3384 26268 3985 26296
rect 3384 26256 3390 26268
rect 3973 26265 3985 26268
rect 4019 26265 4031 26299
rect 3973 26259 4031 26265
rect 4189 26299 4247 26305
rect 4189 26265 4201 26299
rect 4235 26296 4247 26299
rect 4430 26296 4436 26308
rect 4235 26268 4436 26296
rect 4235 26265 4247 26268
rect 4189 26259 4247 26265
rect 4430 26256 4436 26268
rect 4488 26296 4494 26308
rect 4801 26299 4859 26305
rect 4801 26296 4813 26299
rect 4488 26268 4813 26296
rect 4488 26256 4494 26268
rect 4801 26265 4813 26268
rect 4847 26265 4859 26299
rect 4801 26259 4859 26265
rect 2041 26231 2099 26237
rect 2041 26197 2053 26231
rect 2087 26228 2099 26231
rect 2130 26228 2136 26240
rect 2087 26200 2136 26228
rect 2087 26197 2099 26200
rect 2041 26191 2099 26197
rect 2130 26188 2136 26200
rect 2188 26228 2194 26240
rect 3344 26228 3372 26256
rect 4908 26240 4936 26336
rect 5074 26324 5080 26336
rect 5132 26324 5138 26376
rect 6270 26364 6276 26376
rect 6231 26336 6276 26364
rect 6270 26324 6276 26336
rect 6328 26324 6334 26376
rect 7650 26324 7656 26376
rect 7708 26324 7714 26376
rect 9585 26367 9643 26373
rect 9585 26333 9597 26367
rect 9631 26364 9643 26367
rect 10134 26364 10140 26376
rect 9631 26336 10140 26364
rect 9631 26333 9643 26336
rect 9585 26327 9643 26333
rect 10134 26324 10140 26336
rect 10192 26364 10198 26376
rect 10410 26364 10416 26376
rect 10192 26336 10416 26364
rect 10192 26324 10198 26336
rect 10410 26324 10416 26336
rect 10468 26324 10474 26376
rect 13081 26367 13139 26373
rect 13081 26333 13093 26367
rect 13127 26364 13139 26367
rect 13170 26364 13176 26376
rect 13127 26336 13176 26364
rect 13127 26333 13139 26336
rect 13081 26327 13139 26333
rect 13170 26324 13176 26336
rect 13228 26324 13234 26376
rect 14366 26364 14372 26376
rect 14327 26336 14372 26364
rect 14366 26324 14372 26336
rect 14424 26324 14430 26376
rect 14550 26324 14556 26376
rect 14608 26324 14614 26376
rect 16298 26364 16304 26376
rect 16259 26336 16304 26364
rect 16298 26324 16304 26336
rect 16356 26324 16362 26376
rect 18138 26364 18144 26376
rect 18099 26336 18144 26364
rect 18138 26324 18144 26336
rect 18196 26324 18202 26376
rect 21266 26324 21272 26376
rect 21324 26364 21330 26376
rect 21324 26336 21369 26364
rect 21324 26324 21330 26336
rect 23106 26324 23112 26376
rect 23164 26324 23170 26376
rect 25317 26367 25375 26373
rect 25317 26333 25329 26367
rect 25363 26333 25375 26367
rect 25317 26327 25375 26333
rect 25409 26367 25467 26373
rect 25409 26333 25421 26367
rect 25455 26364 25467 26367
rect 25961 26367 26019 26373
rect 25961 26364 25973 26367
rect 25455 26336 25973 26364
rect 25455 26333 25467 26336
rect 25409 26327 25467 26333
rect 25961 26333 25973 26336
rect 26007 26333 26019 26367
rect 25961 26327 26019 26333
rect 11790 26256 11796 26308
rect 11848 26256 11854 26308
rect 16568 26299 16626 26305
rect 16568 26265 16580 26299
rect 16614 26296 16626 26299
rect 16758 26296 16764 26308
rect 16614 26268 16764 26296
rect 16614 26265 16626 26268
rect 16568 26259 16626 26265
rect 16758 26256 16764 26268
rect 16816 26256 16822 26308
rect 20346 26256 20352 26308
rect 20404 26256 20410 26308
rect 20714 26256 20720 26308
rect 20772 26296 20778 26308
rect 20993 26299 21051 26305
rect 20993 26296 21005 26299
rect 20772 26268 21005 26296
rect 20772 26256 20778 26268
rect 20993 26265 21005 26268
rect 21039 26265 21051 26299
rect 25332 26296 25360 26327
rect 26142 26296 26148 26308
rect 25332 26268 26148 26296
rect 20993 26259 21051 26265
rect 26142 26256 26148 26268
rect 26200 26256 26206 26308
rect 26694 26256 26700 26308
rect 26752 26256 26758 26308
rect 4338 26228 4344 26240
rect 2188 26200 3372 26228
rect 4299 26200 4344 26228
rect 2188 26188 2194 26200
rect 4338 26188 4344 26200
rect 4396 26188 4402 26240
rect 4890 26188 4896 26240
rect 4948 26228 4954 26240
rect 4985 26231 5043 26237
rect 4985 26228 4997 26231
rect 4948 26200 4997 26228
rect 4948 26188 4954 26200
rect 4985 26197 4997 26200
rect 5031 26197 5043 26231
rect 4985 26191 5043 26197
rect 8662 26188 8668 26240
rect 8720 26228 8726 26240
rect 9493 26231 9551 26237
rect 9493 26228 9505 26231
rect 8720 26200 9505 26228
rect 8720 26188 8726 26200
rect 9493 26197 9505 26200
rect 9539 26197 9551 26231
rect 9493 26191 9551 26197
rect 12066 26188 12072 26240
rect 12124 26228 12130 26240
rect 12250 26228 12256 26240
rect 12124 26200 12256 26228
rect 12124 26188 12130 26200
rect 12250 26188 12256 26200
rect 12308 26188 12314 26240
rect 18233 26231 18291 26237
rect 18233 26197 18245 26231
rect 18279 26228 18291 26231
rect 18782 26228 18788 26240
rect 18279 26200 18788 26228
rect 18279 26197 18291 26200
rect 18233 26191 18291 26197
rect 18782 26188 18788 26200
rect 18840 26188 18846 26240
rect 19521 26231 19579 26237
rect 19521 26197 19533 26231
rect 19567 26228 19579 26231
rect 19702 26228 19708 26240
rect 19567 26200 19708 26228
rect 19567 26197 19579 26200
rect 19521 26191 19579 26197
rect 19702 26188 19708 26200
rect 19760 26188 19766 26240
rect 1104 26138 29048 26160
rect 1104 26086 7896 26138
rect 7948 26086 7960 26138
rect 8012 26086 8024 26138
rect 8076 26086 8088 26138
rect 8140 26086 8152 26138
rect 8204 26086 14842 26138
rect 14894 26086 14906 26138
rect 14958 26086 14970 26138
rect 15022 26086 15034 26138
rect 15086 26086 15098 26138
rect 15150 26086 21788 26138
rect 21840 26086 21852 26138
rect 21904 26086 21916 26138
rect 21968 26086 21980 26138
rect 22032 26086 22044 26138
rect 22096 26086 28734 26138
rect 28786 26086 28798 26138
rect 28850 26086 28862 26138
rect 28914 26086 28926 26138
rect 28978 26086 28990 26138
rect 29042 26086 29048 26138
rect 1104 26064 29048 26086
rect 2593 26027 2651 26033
rect 2593 25993 2605 26027
rect 2639 26024 2651 26027
rect 2774 26024 2780 26036
rect 2639 25996 2780 26024
rect 2639 25993 2651 25996
rect 2593 25987 2651 25993
rect 2774 25984 2780 25996
rect 2832 25984 2838 26036
rect 4430 26024 4436 26036
rect 4391 25996 4436 26024
rect 4430 25984 4436 25996
rect 4488 25984 4494 26036
rect 4893 26027 4951 26033
rect 4893 25993 4905 26027
rect 4939 25993 4951 26027
rect 9490 26024 9496 26036
rect 4893 25987 4951 25993
rect 7300 25996 9496 26024
rect 3320 25959 3378 25965
rect 3320 25925 3332 25959
rect 3366 25956 3378 25959
rect 4908 25956 4936 25987
rect 3366 25928 4936 25956
rect 3366 25925 3378 25928
rect 3320 25919 3378 25925
rect 2130 25888 2136 25900
rect 2091 25860 2136 25888
rect 2130 25848 2136 25860
rect 2188 25848 2194 25900
rect 2409 25891 2467 25897
rect 2409 25857 2421 25891
rect 2455 25888 2467 25891
rect 2455 25860 4108 25888
rect 2455 25857 2467 25860
rect 2409 25851 2467 25857
rect 2866 25780 2872 25832
rect 2924 25820 2930 25832
rect 3053 25823 3111 25829
rect 3053 25820 3065 25823
rect 2924 25792 3065 25820
rect 2924 25780 2930 25792
rect 3053 25789 3065 25792
rect 3099 25789 3111 25823
rect 4080 25820 4108 25860
rect 4338 25848 4344 25900
rect 4396 25888 4402 25900
rect 4893 25891 4951 25897
rect 4893 25888 4905 25891
rect 4396 25860 4905 25888
rect 4396 25848 4402 25860
rect 4893 25857 4905 25860
rect 4939 25857 4951 25891
rect 4893 25851 4951 25857
rect 4982 25848 4988 25900
rect 5040 25888 5046 25900
rect 5040 25860 5085 25888
rect 7300 25874 7328 25996
rect 9490 25984 9496 25996
rect 9548 25984 9554 26036
rect 10134 26024 10140 26036
rect 10095 25996 10140 26024
rect 10134 25984 10140 25996
rect 10192 25984 10198 26036
rect 12253 26027 12311 26033
rect 12253 25993 12265 26027
rect 12299 26024 12311 26027
rect 12526 26024 12532 26036
rect 12299 25996 12532 26024
rect 12299 25993 12311 25996
rect 12253 25987 12311 25993
rect 12526 25984 12532 25996
rect 12584 25984 12590 26036
rect 17313 26027 17371 26033
rect 17313 25993 17325 26027
rect 17359 26024 17371 26027
rect 18138 26024 18144 26036
rect 17359 25996 18144 26024
rect 17359 25993 17371 25996
rect 17313 25987 17371 25993
rect 18138 25984 18144 25996
rect 18196 25984 18202 26036
rect 20257 26027 20315 26033
rect 20257 25993 20269 26027
rect 20303 26024 20315 26027
rect 20714 26024 20720 26036
rect 20303 25996 20720 26024
rect 20303 25993 20315 25996
rect 20257 25987 20315 25993
rect 20714 25984 20720 25996
rect 20772 25984 20778 26036
rect 20901 26027 20959 26033
rect 20901 25993 20913 26027
rect 20947 26024 20959 26027
rect 21266 26024 21272 26036
rect 20947 25996 21272 26024
rect 20947 25993 20959 25996
rect 20901 25987 20959 25993
rect 21266 25984 21272 25996
rect 21324 25984 21330 26036
rect 22278 25984 22284 26036
rect 22336 25984 22342 26036
rect 23106 26024 23112 26036
rect 23067 25996 23112 26024
rect 23106 25984 23112 25996
rect 23164 25984 23170 26036
rect 23934 26024 23940 26036
rect 23895 25996 23940 26024
rect 23934 25984 23940 25996
rect 23992 25984 23998 26036
rect 7650 25956 7656 25968
rect 7611 25928 7656 25956
rect 7650 25916 7656 25928
rect 7708 25916 7714 25968
rect 8662 25956 8668 25968
rect 8623 25928 8668 25956
rect 8662 25916 8668 25928
rect 8720 25916 8726 25968
rect 9674 25916 9680 25968
rect 9732 25916 9738 25968
rect 13541 25959 13599 25965
rect 13541 25925 13553 25959
rect 13587 25956 13599 25959
rect 14369 25959 14427 25965
rect 14369 25956 14381 25959
rect 13587 25928 14381 25956
rect 13587 25925 13599 25928
rect 13541 25919 13599 25925
rect 14369 25925 14381 25928
rect 14415 25925 14427 25959
rect 14369 25919 14427 25925
rect 15378 25916 15384 25968
rect 15436 25916 15442 25968
rect 18230 25916 18236 25968
rect 18288 25916 18294 25968
rect 18782 25956 18788 25968
rect 18743 25928 18788 25956
rect 18782 25916 18788 25928
rect 18840 25916 18846 25968
rect 22296 25956 22324 25984
rect 21008 25928 22324 25956
rect 8386 25888 8392 25900
rect 8347 25860 8392 25888
rect 5040 25848 5046 25860
rect 8386 25848 8392 25860
rect 8444 25848 8450 25900
rect 12066 25848 12072 25900
rect 12124 25888 12130 25900
rect 12161 25891 12219 25897
rect 12161 25888 12173 25891
rect 12124 25860 12173 25888
rect 12124 25848 12130 25860
rect 12161 25857 12173 25860
rect 12207 25857 12219 25891
rect 12161 25851 12219 25857
rect 13633 25891 13691 25897
rect 13633 25857 13645 25891
rect 13679 25888 13691 25891
rect 19702 25888 19708 25900
rect 13679 25860 13952 25888
rect 19663 25860 19708 25888
rect 13679 25857 13691 25860
rect 13633 25851 13691 25857
rect 4798 25820 4804 25832
rect 4080 25792 4804 25820
rect 3053 25783 3111 25789
rect 4798 25780 4804 25792
rect 4856 25780 4862 25832
rect 5169 25823 5227 25829
rect 5169 25789 5181 25823
rect 5215 25820 5227 25823
rect 5258 25820 5264 25832
rect 5215 25792 5264 25820
rect 5215 25789 5227 25792
rect 5169 25783 5227 25789
rect 5258 25780 5264 25792
rect 5316 25780 5322 25832
rect 6638 25780 6644 25832
rect 6696 25820 6702 25832
rect 6825 25823 6883 25829
rect 6825 25820 6837 25823
rect 6696 25792 6837 25820
rect 6696 25780 6702 25792
rect 6825 25789 6837 25792
rect 6871 25820 6883 25823
rect 8754 25820 8760 25832
rect 6871 25792 8760 25820
rect 6871 25789 6883 25792
rect 6825 25783 6883 25789
rect 8754 25780 8760 25792
rect 8812 25780 8818 25832
rect 2225 25687 2283 25693
rect 2225 25653 2237 25687
rect 2271 25684 2283 25687
rect 4154 25684 4160 25696
rect 2271 25656 4160 25684
rect 2271 25653 2283 25656
rect 2225 25647 2283 25653
rect 4154 25644 4160 25656
rect 4212 25644 4218 25696
rect 13924 25684 13952 25860
rect 19702 25848 19708 25860
rect 19760 25888 19766 25900
rect 21008 25897 21036 25928
rect 20165 25891 20223 25897
rect 20165 25888 20177 25891
rect 19760 25860 20177 25888
rect 19760 25848 19766 25860
rect 20165 25857 20177 25860
rect 20211 25857 20223 25891
rect 20165 25851 20223 25857
rect 20993 25891 21051 25897
rect 20993 25857 21005 25891
rect 21039 25857 21051 25891
rect 22462 25888 22468 25900
rect 22423 25860 22468 25888
rect 20993 25851 21051 25857
rect 22462 25848 22468 25860
rect 22520 25888 22526 25900
rect 25774 25888 25780 25900
rect 22520 25860 25780 25888
rect 22520 25848 22526 25860
rect 25774 25848 25780 25860
rect 25832 25848 25838 25900
rect 26142 25848 26148 25900
rect 26200 25888 26206 25900
rect 27157 25891 27215 25897
rect 27157 25888 27169 25891
rect 26200 25860 27169 25888
rect 26200 25848 26206 25860
rect 27157 25857 27169 25860
rect 27203 25857 27215 25891
rect 27157 25851 27215 25857
rect 14090 25820 14096 25832
rect 14051 25792 14096 25820
rect 14090 25780 14096 25792
rect 14148 25780 14154 25832
rect 19061 25823 19119 25829
rect 19061 25789 19073 25823
rect 19107 25820 19119 25823
rect 19613 25823 19671 25829
rect 19613 25820 19625 25823
rect 19107 25792 19625 25820
rect 19107 25789 19119 25792
rect 19061 25783 19119 25789
rect 19613 25789 19625 25792
rect 19659 25789 19671 25823
rect 19613 25783 19671 25789
rect 19978 25780 19984 25832
rect 20036 25820 20042 25832
rect 22189 25823 22247 25829
rect 22189 25820 22201 25823
rect 20036 25792 22201 25820
rect 20036 25780 20042 25792
rect 22189 25789 22201 25792
rect 22235 25789 22247 25823
rect 24026 25820 24032 25832
rect 23987 25792 24032 25820
rect 22189 25783 22247 25789
rect 24026 25780 24032 25792
rect 24084 25780 24090 25832
rect 24121 25823 24179 25829
rect 24121 25789 24133 25823
rect 24167 25789 24179 25823
rect 24121 25783 24179 25789
rect 23658 25712 23664 25764
rect 23716 25752 23722 25764
rect 24136 25752 24164 25783
rect 23716 25724 24164 25752
rect 25792 25752 25820 25848
rect 26050 25820 26056 25832
rect 26011 25792 26056 25820
rect 26050 25780 26056 25792
rect 26108 25780 26114 25832
rect 26510 25820 26516 25832
rect 26471 25792 26516 25820
rect 26510 25780 26516 25792
rect 26568 25780 26574 25832
rect 27430 25752 27436 25764
rect 25792 25724 27436 25752
rect 23716 25712 23722 25724
rect 27430 25712 27436 25724
rect 27488 25712 27494 25764
rect 15654 25684 15660 25696
rect 13924 25656 15660 25684
rect 15654 25644 15660 25656
rect 15712 25684 15718 25696
rect 15841 25687 15899 25693
rect 15841 25684 15853 25687
rect 15712 25656 15853 25684
rect 15712 25644 15718 25656
rect 15841 25653 15853 25656
rect 15887 25653 15899 25687
rect 23566 25684 23572 25696
rect 23527 25656 23572 25684
rect 15841 25647 15899 25653
rect 23566 25644 23572 25656
rect 23624 25644 23630 25696
rect 27249 25687 27307 25693
rect 27249 25653 27261 25687
rect 27295 25684 27307 25687
rect 27522 25684 27528 25696
rect 27295 25656 27528 25684
rect 27295 25653 27307 25656
rect 27249 25647 27307 25653
rect 27522 25644 27528 25656
rect 27580 25644 27586 25696
rect 1104 25594 28888 25616
rect 1104 25542 4423 25594
rect 4475 25542 4487 25594
rect 4539 25542 4551 25594
rect 4603 25542 4615 25594
rect 4667 25542 4679 25594
rect 4731 25542 11369 25594
rect 11421 25542 11433 25594
rect 11485 25542 11497 25594
rect 11549 25542 11561 25594
rect 11613 25542 11625 25594
rect 11677 25542 18315 25594
rect 18367 25542 18379 25594
rect 18431 25542 18443 25594
rect 18495 25542 18507 25594
rect 18559 25542 18571 25594
rect 18623 25542 25261 25594
rect 25313 25542 25325 25594
rect 25377 25542 25389 25594
rect 25441 25542 25453 25594
rect 25505 25542 25517 25594
rect 25569 25542 28888 25594
rect 1104 25520 28888 25542
rect 3329 25483 3387 25489
rect 3329 25449 3341 25483
rect 3375 25480 3387 25483
rect 4246 25480 4252 25492
rect 3375 25452 4252 25480
rect 3375 25449 3387 25452
rect 3329 25443 3387 25449
rect 4246 25440 4252 25452
rect 4304 25440 4310 25492
rect 4798 25440 4804 25492
rect 4856 25480 4862 25492
rect 5261 25483 5319 25489
rect 5261 25480 5273 25483
rect 4856 25452 5273 25480
rect 4856 25440 4862 25452
rect 5261 25449 5273 25452
rect 5307 25449 5319 25483
rect 5261 25443 5319 25449
rect 6181 25483 6239 25489
rect 6181 25449 6193 25483
rect 6227 25480 6239 25483
rect 6270 25480 6276 25492
rect 6227 25452 6276 25480
rect 6227 25449 6239 25452
rect 6181 25443 6239 25449
rect 6270 25440 6276 25452
rect 6328 25440 6334 25492
rect 13633 25483 13691 25489
rect 13633 25449 13645 25483
rect 13679 25480 13691 25483
rect 14090 25480 14096 25492
rect 13679 25452 14096 25480
rect 13679 25449 13691 25452
rect 13633 25443 13691 25449
rect 14090 25440 14096 25452
rect 14148 25440 14154 25492
rect 22649 25483 22707 25489
rect 22649 25449 22661 25483
rect 22695 25480 22707 25483
rect 22922 25480 22928 25492
rect 22695 25452 22928 25480
rect 22695 25449 22707 25452
rect 22649 25443 22707 25449
rect 22922 25440 22928 25452
rect 22980 25440 22986 25492
rect 8113 25415 8171 25421
rect 8113 25381 8125 25415
rect 8159 25381 8171 25415
rect 19794 25412 19800 25424
rect 8113 25375 8171 25381
rect 17880 25384 19800 25412
rect 5074 25304 5080 25356
rect 5132 25304 5138 25356
rect 7742 25304 7748 25356
rect 7800 25344 7806 25356
rect 8128 25344 8156 25375
rect 9217 25347 9275 25353
rect 9217 25344 9229 25347
rect 7800 25316 9229 25344
rect 7800 25304 7806 25316
rect 9217 25313 9229 25316
rect 9263 25313 9275 25347
rect 9217 25307 9275 25313
rect 9677 25347 9735 25353
rect 9677 25313 9689 25347
rect 9723 25344 9735 25347
rect 11238 25344 11244 25356
rect 9723 25316 11244 25344
rect 9723 25313 9735 25316
rect 9677 25307 9735 25313
rect 11238 25304 11244 25316
rect 11296 25304 11302 25356
rect 11790 25344 11796 25356
rect 11751 25316 11796 25344
rect 11790 25304 11796 25316
rect 11848 25304 11854 25356
rect 14550 25344 14556 25356
rect 13648 25316 14556 25344
rect 3142 25276 3148 25288
rect 3103 25248 3148 25276
rect 3142 25236 3148 25248
rect 3200 25236 3206 25288
rect 3421 25279 3479 25285
rect 3421 25245 3433 25279
rect 3467 25276 3479 25279
rect 4154 25276 4160 25288
rect 3467 25248 4160 25276
rect 3467 25245 3479 25248
rect 3421 25239 3479 25245
rect 4154 25236 4160 25248
rect 4212 25236 4218 25288
rect 4249 25279 4307 25285
rect 4249 25245 4261 25279
rect 4295 25276 4307 25279
rect 4338 25276 4344 25288
rect 4295 25248 4344 25276
rect 4295 25245 4307 25248
rect 4249 25239 4307 25245
rect 4338 25236 4344 25248
rect 4396 25236 4402 25288
rect 4985 25279 5043 25285
rect 4985 25276 4997 25279
rect 4448 25248 4997 25276
rect 4448 25208 4476 25248
rect 4985 25245 4997 25248
rect 5031 25276 5043 25279
rect 5092 25276 5120 25304
rect 5031 25248 5120 25276
rect 6273 25279 6331 25285
rect 5031 25245 5043 25248
rect 4985 25239 5043 25245
rect 6273 25245 6285 25279
rect 6319 25276 6331 25279
rect 6362 25276 6368 25288
rect 6319 25248 6368 25276
rect 6319 25245 6331 25248
rect 6273 25239 6331 25245
rect 6362 25236 6368 25248
rect 6420 25236 6426 25288
rect 6733 25279 6791 25285
rect 6733 25245 6745 25279
rect 6779 25276 6791 25279
rect 9306 25276 9312 25288
rect 6779 25248 6914 25276
rect 9267 25248 9312 25276
rect 6779 25245 6791 25248
rect 6733 25239 6791 25245
rect 4356 25180 4476 25208
rect 4525 25211 4583 25217
rect 2958 25140 2964 25152
rect 2919 25112 2964 25140
rect 2958 25100 2964 25112
rect 3016 25100 3022 25152
rect 3973 25143 4031 25149
rect 3973 25109 3985 25143
rect 4019 25140 4031 25143
rect 4062 25140 4068 25152
rect 4019 25112 4068 25140
rect 4019 25109 4031 25112
rect 3973 25103 4031 25109
rect 4062 25100 4068 25112
rect 4120 25100 4126 25152
rect 4246 25100 4252 25152
rect 4304 25140 4310 25152
rect 4356 25149 4384 25180
rect 4525 25177 4537 25211
rect 4571 25208 4583 25211
rect 4890 25208 4896 25220
rect 4571 25180 4896 25208
rect 4571 25177 4583 25180
rect 4525 25171 4583 25177
rect 4890 25168 4896 25180
rect 4948 25208 4954 25220
rect 5077 25211 5135 25217
rect 5077 25208 5089 25211
rect 4948 25180 5089 25208
rect 4948 25168 4954 25180
rect 5077 25177 5089 25180
rect 5123 25177 5135 25211
rect 5258 25208 5264 25220
rect 5219 25180 5264 25208
rect 5077 25171 5135 25177
rect 5258 25168 5264 25180
rect 5316 25168 5322 25220
rect 4341 25143 4399 25149
rect 4341 25140 4353 25143
rect 4304 25112 4353 25140
rect 4304 25100 4310 25112
rect 4341 25109 4353 25112
rect 4387 25109 4399 25143
rect 6886 25140 6914 25248
rect 9306 25236 9312 25248
rect 9364 25236 9370 25288
rect 9950 25236 9956 25288
rect 10008 25276 10014 25288
rect 10873 25279 10931 25285
rect 10873 25276 10885 25279
rect 10008 25248 10885 25276
rect 10008 25236 10014 25248
rect 10873 25245 10885 25248
rect 10919 25245 10931 25279
rect 10873 25239 10931 25245
rect 7000 25211 7058 25217
rect 7000 25177 7012 25211
rect 7046 25208 7058 25211
rect 7466 25208 7472 25220
rect 7046 25180 7472 25208
rect 7046 25177 7058 25180
rect 7000 25171 7058 25177
rect 7466 25168 7472 25180
rect 7524 25168 7530 25220
rect 9490 25168 9496 25220
rect 9548 25208 9554 25220
rect 10980 25208 11008 25262
rect 13170 25236 13176 25288
rect 13228 25276 13234 25288
rect 13541 25279 13599 25285
rect 13541 25276 13553 25279
rect 13228 25248 13553 25276
rect 13228 25236 13234 25248
rect 13541 25245 13553 25248
rect 13587 25245 13599 25279
rect 13541 25239 13599 25245
rect 13648 25208 13676 25316
rect 14366 25276 14372 25288
rect 14327 25248 14372 25276
rect 14366 25236 14372 25248
rect 14424 25236 14430 25288
rect 14476 25262 14504 25316
rect 14550 25304 14556 25316
rect 14608 25304 14614 25356
rect 15378 25344 15384 25356
rect 15339 25316 15384 25344
rect 15378 25304 15384 25316
rect 15436 25304 15442 25356
rect 17880 25344 17908 25384
rect 19794 25372 19800 25384
rect 19852 25372 19858 25424
rect 17788 25316 17908 25344
rect 17788 25285 17816 25316
rect 18230 25304 18236 25356
rect 18288 25344 18294 25356
rect 18325 25347 18383 25353
rect 18325 25344 18337 25347
rect 18288 25316 18337 25344
rect 18288 25304 18294 25316
rect 18325 25313 18337 25316
rect 18371 25313 18383 25347
rect 22940 25344 22968 25440
rect 23569 25347 23627 25353
rect 23569 25344 23581 25347
rect 22940 25316 23581 25344
rect 18325 25307 18383 25313
rect 23569 25313 23581 25316
rect 23615 25313 23627 25347
rect 23569 25307 23627 25313
rect 23658 25304 23664 25356
rect 23716 25344 23722 25356
rect 23716 25316 23761 25344
rect 23716 25304 23722 25316
rect 24026 25304 24032 25356
rect 24084 25344 24090 25356
rect 24673 25347 24731 25353
rect 24673 25344 24685 25347
rect 24084 25316 24685 25344
rect 24084 25304 24090 25316
rect 24673 25313 24685 25316
rect 24719 25313 24731 25347
rect 24673 25307 24731 25313
rect 25038 25304 25044 25356
rect 25096 25344 25102 25356
rect 25133 25347 25191 25353
rect 25133 25344 25145 25347
rect 25096 25316 25145 25344
rect 25096 25304 25102 25316
rect 25133 25313 25145 25316
rect 25179 25313 25191 25347
rect 25133 25307 25191 25313
rect 26053 25347 26111 25353
rect 26053 25313 26065 25347
rect 26099 25344 26111 25347
rect 26142 25344 26148 25356
rect 26099 25316 26148 25344
rect 26099 25313 26111 25316
rect 26053 25307 26111 25313
rect 17773 25279 17831 25285
rect 17773 25245 17785 25279
rect 17819 25245 17831 25279
rect 17773 25239 17831 25245
rect 17865 25279 17923 25285
rect 17865 25245 17877 25279
rect 17911 25276 17923 25279
rect 19794 25276 19800 25288
rect 17911 25248 19800 25276
rect 17911 25245 17923 25248
rect 17865 25239 17923 25245
rect 19794 25236 19800 25248
rect 19852 25276 19858 25288
rect 19978 25276 19984 25288
rect 19852 25248 19984 25276
rect 19852 25236 19858 25248
rect 19978 25236 19984 25248
rect 20036 25236 20042 25288
rect 21269 25279 21327 25285
rect 21269 25245 21281 25279
rect 21315 25276 21327 25279
rect 22738 25276 22744 25288
rect 21315 25248 22744 25276
rect 21315 25245 21327 25248
rect 21269 25239 21327 25245
rect 22738 25236 22744 25248
rect 22796 25236 22802 25288
rect 24765 25279 24823 25285
rect 24765 25245 24777 25279
rect 24811 25276 24823 25279
rect 26068 25276 26096 25307
rect 26142 25304 26148 25316
rect 26200 25304 26206 25356
rect 27522 25344 27528 25356
rect 27483 25316 27528 25344
rect 27522 25304 27528 25316
rect 27580 25304 27586 25356
rect 24811 25248 26096 25276
rect 27801 25279 27859 25285
rect 24811 25245 24823 25248
rect 24765 25239 24823 25245
rect 27801 25245 27813 25279
rect 27847 25245 27859 25279
rect 27801 25239 27859 25245
rect 9548 25180 13676 25208
rect 21536 25211 21594 25217
rect 9548 25168 9554 25180
rect 21536 25177 21548 25211
rect 21582 25208 21594 25211
rect 21582 25180 23152 25208
rect 21582 25177 21594 25180
rect 21536 25171 21594 25177
rect 7098 25140 7104 25152
rect 6886 25112 7104 25140
rect 4341 25103 4399 25109
rect 7098 25100 7104 25112
rect 7156 25100 7162 25152
rect 23124 25149 23152 25180
rect 26510 25168 26516 25220
rect 26568 25168 26574 25220
rect 27246 25168 27252 25220
rect 27304 25208 27310 25220
rect 27816 25208 27844 25239
rect 27304 25180 27844 25208
rect 27304 25168 27310 25180
rect 23109 25143 23167 25149
rect 23109 25109 23121 25143
rect 23155 25109 23167 25143
rect 23474 25140 23480 25152
rect 23435 25112 23480 25140
rect 23109 25103 23167 25109
rect 23474 25100 23480 25112
rect 23532 25140 23538 25152
rect 23750 25140 23756 25152
rect 23532 25112 23756 25140
rect 23532 25100 23538 25112
rect 23750 25100 23756 25112
rect 23808 25140 23814 25152
rect 28074 25140 28080 25152
rect 23808 25112 28080 25140
rect 23808 25100 23814 25112
rect 28074 25100 28080 25112
rect 28132 25100 28138 25152
rect 1104 25050 29048 25072
rect 1104 24998 7896 25050
rect 7948 24998 7960 25050
rect 8012 24998 8024 25050
rect 8076 24998 8088 25050
rect 8140 24998 8152 25050
rect 8204 24998 14842 25050
rect 14894 24998 14906 25050
rect 14958 24998 14970 25050
rect 15022 24998 15034 25050
rect 15086 24998 15098 25050
rect 15150 24998 21788 25050
rect 21840 24998 21852 25050
rect 21904 24998 21916 25050
rect 21968 24998 21980 25050
rect 22032 24998 22044 25050
rect 22096 24998 28734 25050
rect 28786 24998 28798 25050
rect 28850 24998 28862 25050
rect 28914 24998 28926 25050
rect 28978 24998 28990 25050
rect 29042 24998 29048 25050
rect 1104 24976 29048 24998
rect 4154 24896 4160 24948
rect 4212 24936 4218 24948
rect 4249 24939 4307 24945
rect 4249 24936 4261 24939
rect 4212 24908 4261 24936
rect 4212 24896 4218 24908
rect 4249 24905 4261 24908
rect 4295 24905 4307 24939
rect 7466 24936 7472 24948
rect 7427 24908 7472 24936
rect 4249 24899 4307 24905
rect 7466 24896 7472 24908
rect 7524 24896 7530 24948
rect 7742 24896 7748 24948
rect 7800 24936 7806 24948
rect 7929 24939 7987 24945
rect 7929 24936 7941 24939
rect 7800 24908 7941 24936
rect 7800 24896 7806 24908
rect 7929 24905 7941 24908
rect 7975 24905 7987 24939
rect 7929 24899 7987 24905
rect 12069 24939 12127 24945
rect 12069 24905 12081 24939
rect 12115 24936 12127 24939
rect 23474 24936 23480 24948
rect 12115 24908 23480 24936
rect 12115 24905 12127 24908
rect 12069 24899 12127 24905
rect 23474 24896 23480 24908
rect 23532 24896 23538 24948
rect 24026 24896 24032 24948
rect 24084 24936 24090 24948
rect 24213 24939 24271 24945
rect 24213 24936 24225 24939
rect 24084 24908 24225 24936
rect 24084 24896 24090 24908
rect 24213 24905 24225 24908
rect 24259 24905 24271 24939
rect 24213 24899 24271 24905
rect 2038 24828 2044 24880
rect 2096 24868 2102 24880
rect 3970 24868 3976 24880
rect 2096 24840 3976 24868
rect 2096 24828 2102 24840
rect 3970 24828 3976 24840
rect 4028 24828 4034 24880
rect 7837 24871 7895 24877
rect 7837 24837 7849 24871
rect 7883 24868 7895 24871
rect 9490 24868 9496 24880
rect 7883 24840 9496 24868
rect 7883 24837 7895 24840
rect 7837 24831 7895 24837
rect 9490 24828 9496 24840
rect 9548 24868 9554 24880
rect 14274 24868 14280 24880
rect 9548 24840 14280 24868
rect 9548 24828 9554 24840
rect 14274 24828 14280 24840
rect 14332 24828 14338 24880
rect 23382 24828 23388 24880
rect 23440 24868 23446 24880
rect 23440 24840 23704 24868
rect 23440 24828 23446 24840
rect 2958 24760 2964 24812
rect 3016 24800 3022 24812
rect 3125 24803 3183 24809
rect 3125 24800 3137 24803
rect 3016 24772 3137 24800
rect 3016 24760 3022 24772
rect 3125 24769 3137 24772
rect 3171 24769 3183 24803
rect 3125 24763 3183 24769
rect 10781 24803 10839 24809
rect 10781 24769 10793 24803
rect 10827 24800 10839 24803
rect 12066 24800 12072 24812
rect 10827 24772 12072 24800
rect 10827 24769 10839 24772
rect 10781 24763 10839 24769
rect 12066 24760 12072 24772
rect 12124 24760 12130 24812
rect 14645 24803 14703 24809
rect 14645 24769 14657 24803
rect 14691 24800 14703 24803
rect 15654 24800 15660 24812
rect 14691 24772 15660 24800
rect 14691 24769 14703 24772
rect 14645 24763 14703 24769
rect 15654 24760 15660 24772
rect 15712 24760 15718 24812
rect 17126 24809 17132 24812
rect 17120 24763 17132 24809
rect 17184 24800 17190 24812
rect 17184 24772 17220 24800
rect 17126 24760 17132 24763
rect 17184 24760 17190 24772
rect 18138 24760 18144 24812
rect 18196 24800 18202 24812
rect 18877 24803 18935 24809
rect 18877 24800 18889 24803
rect 18196 24772 18889 24800
rect 18196 24760 18202 24772
rect 18877 24769 18889 24772
rect 18923 24769 18935 24803
rect 18877 24763 18935 24769
rect 23100 24803 23158 24809
rect 23100 24769 23112 24803
rect 23146 24800 23158 24803
rect 23566 24800 23572 24812
rect 23146 24772 23572 24800
rect 23146 24769 23158 24772
rect 23100 24763 23158 24769
rect 23566 24760 23572 24772
rect 23624 24760 23630 24812
rect 23676 24800 23704 24840
rect 24780 24840 24992 24868
rect 24780 24800 24808 24840
rect 24964 24809 24992 24840
rect 23676 24772 24808 24800
rect 24857 24803 24915 24809
rect 24857 24769 24869 24803
rect 24903 24769 24915 24803
rect 24857 24763 24915 24769
rect 24949 24803 25007 24809
rect 24949 24769 24961 24803
rect 24995 24769 25007 24803
rect 25130 24800 25136 24812
rect 25091 24772 25136 24800
rect 24949 24763 25007 24769
rect 2866 24732 2872 24744
rect 2827 24704 2872 24732
rect 2866 24692 2872 24704
rect 2924 24692 2930 24744
rect 7742 24692 7748 24744
rect 7800 24732 7806 24744
rect 8021 24735 8079 24741
rect 8021 24732 8033 24735
rect 7800 24704 8033 24732
rect 7800 24692 7806 24704
rect 8021 24701 8033 24704
rect 8067 24701 8079 24735
rect 8021 24695 8079 24701
rect 10873 24735 10931 24741
rect 10873 24701 10885 24735
rect 10919 24732 10931 24735
rect 11790 24732 11796 24744
rect 10919 24704 11796 24732
rect 10919 24701 10931 24704
rect 10873 24695 10931 24701
rect 11790 24692 11796 24704
rect 11848 24732 11854 24744
rect 12161 24735 12219 24741
rect 12161 24732 12173 24735
rect 11848 24704 12173 24732
rect 11848 24692 11854 24704
rect 12161 24701 12173 24704
rect 12207 24701 12219 24735
rect 12342 24732 12348 24744
rect 12303 24704 12348 24732
rect 12161 24695 12219 24701
rect 12342 24692 12348 24704
rect 12400 24692 12406 24744
rect 14734 24732 14740 24744
rect 14647 24704 14740 24732
rect 14734 24692 14740 24704
rect 14792 24732 14798 24744
rect 15010 24732 15016 24744
rect 14792 24704 15016 24732
rect 14792 24692 14798 24704
rect 15010 24692 15016 24704
rect 15068 24692 15074 24744
rect 16850 24732 16856 24744
rect 16811 24704 16856 24732
rect 16850 24692 16856 24704
rect 16908 24692 16914 24744
rect 18785 24735 18843 24741
rect 18785 24732 18797 24735
rect 18248 24704 18797 24732
rect 11149 24667 11207 24673
rect 11149 24633 11161 24667
rect 11195 24664 11207 24667
rect 12434 24664 12440 24676
rect 11195 24636 12440 24664
rect 11195 24633 11207 24636
rect 11149 24627 11207 24633
rect 12434 24624 12440 24636
rect 12492 24624 12498 24676
rect 11698 24596 11704 24608
rect 11659 24568 11704 24596
rect 11698 24556 11704 24568
rect 11756 24556 11762 24608
rect 12710 24556 12716 24608
rect 12768 24596 12774 24608
rect 14277 24599 14335 24605
rect 14277 24596 14289 24599
rect 12768 24568 14289 24596
rect 12768 24556 12774 24568
rect 14277 24565 14289 24568
rect 14323 24565 14335 24599
rect 14277 24559 14335 24565
rect 17494 24556 17500 24608
rect 17552 24596 17558 24608
rect 18248 24605 18276 24704
rect 18785 24701 18797 24704
rect 18831 24701 18843 24735
rect 18785 24695 18843 24701
rect 22738 24692 22744 24744
rect 22796 24732 22802 24744
rect 22833 24735 22891 24741
rect 22833 24732 22845 24735
rect 22796 24704 22845 24732
rect 22796 24692 22802 24704
rect 22833 24701 22845 24704
rect 22879 24701 22891 24735
rect 22833 24695 22891 24701
rect 24872 24664 24900 24763
rect 25130 24760 25136 24772
rect 25188 24760 25194 24812
rect 26142 24800 26148 24812
rect 26103 24772 26148 24800
rect 26142 24760 26148 24772
rect 26200 24760 26206 24812
rect 26053 24735 26111 24741
rect 26053 24701 26065 24735
rect 26099 24732 26111 24735
rect 27246 24732 27252 24744
rect 26099 24704 27252 24732
rect 26099 24701 26111 24704
rect 26053 24695 26111 24701
rect 27246 24692 27252 24704
rect 27304 24692 27310 24744
rect 23768 24636 24900 24664
rect 18233 24599 18291 24605
rect 18233 24596 18245 24599
rect 17552 24568 18245 24596
rect 17552 24556 17558 24568
rect 18233 24565 18245 24568
rect 18279 24565 18291 24599
rect 18233 24559 18291 24565
rect 19245 24599 19303 24605
rect 19245 24565 19257 24599
rect 19291 24596 19303 24599
rect 23768 24596 23796 24636
rect 24670 24596 24676 24608
rect 19291 24568 23796 24596
rect 24631 24568 24676 24596
rect 19291 24565 19303 24568
rect 19245 24559 19303 24565
rect 24670 24556 24676 24568
rect 24728 24556 24734 24608
rect 25038 24596 25044 24608
rect 24999 24568 25044 24596
rect 25038 24556 25044 24568
rect 25096 24556 25102 24608
rect 1104 24506 28888 24528
rect 1104 24454 4423 24506
rect 4475 24454 4487 24506
rect 4539 24454 4551 24506
rect 4603 24454 4615 24506
rect 4667 24454 4679 24506
rect 4731 24454 11369 24506
rect 11421 24454 11433 24506
rect 11485 24454 11497 24506
rect 11549 24454 11561 24506
rect 11613 24454 11625 24506
rect 11677 24454 18315 24506
rect 18367 24454 18379 24506
rect 18431 24454 18443 24506
rect 18495 24454 18507 24506
rect 18559 24454 18571 24506
rect 18623 24454 25261 24506
rect 25313 24454 25325 24506
rect 25377 24454 25389 24506
rect 25441 24454 25453 24506
rect 25505 24454 25517 24506
rect 25569 24454 28888 24506
rect 1104 24432 28888 24454
rect 3142 24352 3148 24404
rect 3200 24392 3206 24404
rect 3973 24395 4031 24401
rect 3973 24392 3985 24395
rect 3200 24364 3985 24392
rect 3200 24352 3206 24364
rect 3973 24361 3985 24364
rect 4019 24361 4031 24395
rect 11790 24392 11796 24404
rect 11751 24364 11796 24392
rect 3973 24355 4031 24361
rect 11790 24352 11796 24364
rect 11848 24352 11854 24404
rect 12710 24392 12716 24404
rect 12671 24364 12716 24392
rect 12710 24352 12716 24364
rect 12768 24352 12774 24404
rect 15010 24352 15016 24404
rect 15068 24392 15074 24404
rect 15657 24395 15715 24401
rect 15657 24392 15669 24395
rect 15068 24364 15669 24392
rect 15068 24352 15074 24364
rect 15657 24361 15669 24364
rect 15703 24361 15715 24395
rect 15657 24355 15715 24361
rect 17037 24395 17095 24401
rect 17037 24361 17049 24395
rect 17083 24392 17095 24395
rect 17126 24392 17132 24404
rect 17083 24364 17132 24392
rect 17083 24361 17095 24364
rect 17037 24355 17095 24361
rect 17126 24352 17132 24364
rect 17184 24352 17190 24404
rect 5258 24256 5264 24268
rect 2884 24228 5264 24256
rect 2774 24148 2780 24200
rect 2832 24188 2838 24200
rect 2884 24197 2912 24228
rect 2869 24191 2927 24197
rect 2869 24188 2881 24191
rect 2832 24160 2881 24188
rect 2832 24148 2838 24160
rect 2869 24157 2881 24160
rect 2915 24157 2927 24191
rect 2869 24151 2927 24157
rect 3053 24191 3111 24197
rect 3053 24157 3065 24191
rect 3099 24157 3111 24191
rect 3053 24151 3111 24157
rect 3973 24191 4031 24197
rect 3973 24157 3985 24191
rect 4019 24188 4031 24191
rect 4062 24188 4068 24200
rect 4019 24160 4068 24188
rect 4019 24157 4031 24160
rect 3973 24151 4031 24157
rect 3068 24120 3096 24151
rect 4062 24148 4068 24160
rect 4120 24148 4126 24200
rect 4172 24197 4200 24228
rect 5258 24216 5264 24228
rect 5316 24216 5322 24268
rect 17494 24256 17500 24268
rect 17455 24228 17500 24256
rect 17494 24216 17500 24228
rect 17552 24216 17558 24268
rect 17678 24256 17684 24268
rect 17639 24228 17684 24256
rect 17678 24216 17684 24228
rect 17736 24216 17742 24268
rect 22462 24216 22468 24268
rect 22520 24256 22526 24268
rect 22557 24259 22615 24265
rect 22557 24256 22569 24259
rect 22520 24228 22569 24256
rect 22520 24216 22526 24228
rect 22557 24225 22569 24228
rect 22603 24256 22615 24259
rect 23658 24256 23664 24268
rect 22603 24228 23664 24256
rect 22603 24225 22615 24228
rect 22557 24219 22615 24225
rect 23658 24216 23664 24228
rect 23716 24216 23722 24268
rect 4157 24191 4215 24197
rect 4157 24157 4169 24191
rect 4203 24157 4215 24191
rect 6362 24188 6368 24200
rect 6323 24160 6368 24188
rect 4157 24151 4215 24157
rect 6362 24148 6368 24160
rect 6420 24148 6426 24200
rect 9398 24148 9404 24200
rect 9456 24188 9462 24200
rect 10413 24191 10471 24197
rect 10413 24188 10425 24191
rect 9456 24160 10425 24188
rect 9456 24148 9462 24160
rect 10413 24157 10425 24160
rect 10459 24157 10471 24191
rect 10413 24151 10471 24157
rect 10680 24191 10738 24197
rect 10680 24157 10692 24191
rect 10726 24188 10738 24191
rect 11698 24188 11704 24200
rect 10726 24160 11704 24188
rect 10726 24157 10738 24160
rect 10680 24151 10738 24157
rect 11698 24148 11704 24160
rect 11756 24148 11762 24200
rect 12434 24188 12440 24200
rect 12395 24160 12440 24188
rect 12434 24148 12440 24160
rect 12492 24148 12498 24200
rect 12526 24148 12532 24200
rect 12584 24188 12590 24200
rect 14277 24191 14335 24197
rect 12584 24160 12629 24188
rect 12584 24148 12590 24160
rect 14277 24157 14289 24191
rect 14323 24188 14335 24191
rect 16850 24188 16856 24200
rect 14323 24160 16856 24188
rect 14323 24157 14335 24160
rect 14277 24151 14335 24157
rect 16850 24148 16856 24160
rect 16908 24148 16914 24200
rect 18138 24148 18144 24200
rect 18196 24188 18202 24200
rect 18509 24191 18567 24197
rect 18509 24188 18521 24191
rect 18196 24160 18521 24188
rect 18196 24148 18202 24160
rect 18509 24157 18521 24160
rect 18555 24157 18567 24191
rect 19610 24188 19616 24200
rect 19571 24160 19616 24188
rect 18509 24151 18567 24157
rect 19610 24148 19616 24160
rect 19668 24148 19674 24200
rect 22370 24188 22376 24200
rect 22331 24160 22376 24188
rect 22370 24148 22376 24160
rect 22428 24148 22434 24200
rect 27614 24148 27620 24200
rect 27672 24188 27678 24200
rect 27893 24191 27951 24197
rect 27893 24188 27905 24191
rect 27672 24160 27905 24188
rect 27672 24148 27678 24160
rect 27893 24157 27905 24160
rect 27939 24157 27951 24191
rect 27893 24151 27951 24157
rect 4246 24120 4252 24132
rect 3068 24092 4252 24120
rect 4246 24080 4252 24092
rect 4304 24080 4310 24132
rect 11238 24080 11244 24132
rect 11296 24120 11302 24132
rect 12713 24123 12771 24129
rect 12713 24120 12725 24123
rect 11296 24092 12725 24120
rect 11296 24080 11302 24092
rect 12713 24089 12725 24092
rect 12759 24089 12771 24123
rect 12713 24083 12771 24089
rect 14366 24080 14372 24132
rect 14424 24120 14430 24132
rect 14522 24123 14580 24129
rect 14522 24120 14534 24123
rect 14424 24092 14534 24120
rect 14424 24080 14430 24092
rect 14522 24089 14534 24092
rect 14568 24089 14580 24123
rect 17405 24123 17463 24129
rect 17405 24120 17417 24123
rect 14522 24083 14580 24089
rect 16546 24092 17417 24120
rect 2961 24055 3019 24061
rect 2961 24021 2973 24055
rect 3007 24052 3019 24055
rect 3878 24052 3884 24064
rect 3007 24024 3884 24052
rect 3007 24021 3019 24024
rect 2961 24015 3019 24021
rect 3878 24012 3884 24024
rect 3936 24012 3942 24064
rect 6457 24055 6515 24061
rect 6457 24021 6469 24055
rect 6503 24052 6515 24055
rect 6822 24052 6828 24064
rect 6503 24024 6828 24052
rect 6503 24021 6515 24024
rect 6457 24015 6515 24021
rect 6822 24012 6828 24024
rect 6880 24012 6886 24064
rect 12158 24012 12164 24064
rect 12216 24052 12222 24064
rect 12253 24055 12311 24061
rect 12253 24052 12265 24055
rect 12216 24024 12265 24052
rect 12216 24012 12222 24024
rect 12253 24021 12265 24024
rect 12299 24021 12311 24055
rect 12253 24015 12311 24021
rect 14274 24012 14280 24064
rect 14332 24052 14338 24064
rect 16546 24052 16574 24092
rect 17405 24089 17417 24092
rect 17451 24120 17463 24123
rect 20898 24120 20904 24132
rect 17451 24092 20904 24120
rect 17451 24089 17463 24092
rect 17405 24083 17463 24089
rect 20898 24080 20904 24092
rect 20956 24080 20962 24132
rect 28166 24120 28172 24132
rect 28127 24092 28172 24120
rect 28166 24080 28172 24092
rect 28224 24080 28230 24132
rect 18598 24052 18604 24064
rect 14332 24024 16574 24052
rect 18559 24024 18604 24052
rect 14332 24012 14338 24024
rect 18598 24012 18604 24024
rect 18656 24012 18662 24064
rect 18874 24012 18880 24064
rect 18932 24052 18938 24064
rect 19521 24055 19579 24061
rect 19521 24052 19533 24055
rect 18932 24024 19533 24052
rect 18932 24012 18938 24024
rect 19521 24021 19533 24024
rect 19567 24021 19579 24055
rect 19521 24015 19579 24021
rect 22005 24055 22063 24061
rect 22005 24021 22017 24055
rect 22051 24052 22063 24055
rect 22278 24052 22284 24064
rect 22051 24024 22284 24052
rect 22051 24021 22063 24024
rect 22005 24015 22063 24021
rect 22278 24012 22284 24024
rect 22336 24012 22342 24064
rect 22465 24055 22523 24061
rect 22465 24021 22477 24055
rect 22511 24052 22523 24055
rect 23474 24052 23480 24064
rect 22511 24024 23480 24052
rect 22511 24021 22523 24024
rect 22465 24015 22523 24021
rect 23474 24012 23480 24024
rect 23532 24012 23538 24064
rect 1104 23962 29048 23984
rect 1104 23910 7896 23962
rect 7948 23910 7960 23962
rect 8012 23910 8024 23962
rect 8076 23910 8088 23962
rect 8140 23910 8152 23962
rect 8204 23910 14842 23962
rect 14894 23910 14906 23962
rect 14958 23910 14970 23962
rect 15022 23910 15034 23962
rect 15086 23910 15098 23962
rect 15150 23910 21788 23962
rect 21840 23910 21852 23962
rect 21904 23910 21916 23962
rect 21968 23910 21980 23962
rect 22032 23910 22044 23962
rect 22096 23910 28734 23962
rect 28786 23910 28798 23962
rect 28850 23910 28862 23962
rect 28914 23910 28926 23962
rect 28978 23910 28990 23962
rect 29042 23910 29048 23962
rect 1104 23888 29048 23910
rect 2866 23848 2872 23860
rect 2827 23820 2872 23848
rect 2866 23808 2872 23820
rect 2924 23808 2930 23860
rect 6362 23808 6368 23860
rect 6420 23848 6426 23860
rect 7834 23848 7840 23860
rect 6420 23820 7840 23848
rect 6420 23808 6426 23820
rect 7834 23808 7840 23820
rect 7892 23848 7898 23860
rect 8297 23851 8355 23857
rect 8297 23848 8309 23851
rect 7892 23820 8309 23848
rect 7892 23808 7898 23820
rect 8297 23817 8309 23820
rect 8343 23817 8355 23851
rect 8297 23811 8355 23817
rect 23385 23851 23443 23857
rect 23385 23817 23397 23851
rect 23431 23848 23443 23851
rect 23474 23848 23480 23860
rect 23431 23820 23480 23848
rect 23431 23817 23443 23820
rect 23385 23811 23443 23817
rect 23474 23808 23480 23820
rect 23532 23808 23538 23860
rect 6822 23780 6828 23792
rect 6783 23752 6828 23780
rect 6822 23740 6828 23752
rect 6880 23740 6886 23792
rect 7282 23740 7288 23792
rect 7340 23740 7346 23792
rect 18874 23780 18880 23792
rect 18835 23752 18880 23780
rect 18874 23740 18880 23752
rect 18932 23740 18938 23792
rect 19426 23740 19432 23792
rect 19484 23740 19490 23792
rect 22278 23789 22284 23792
rect 22272 23780 22284 23789
rect 22239 23752 22284 23780
rect 22272 23743 22284 23752
rect 22278 23740 22284 23743
rect 22336 23740 22342 23792
rect 26050 23740 26056 23792
rect 26108 23780 26114 23792
rect 26108 23752 27384 23780
rect 26108 23740 26114 23752
rect 4338 23712 4344 23724
rect 4299 23684 4344 23712
rect 4338 23672 4344 23684
rect 4396 23672 4402 23724
rect 14274 23672 14280 23724
rect 14332 23712 14338 23724
rect 15105 23715 15163 23721
rect 15105 23712 15117 23715
rect 14332 23684 15117 23712
rect 14332 23672 14338 23684
rect 15105 23681 15117 23684
rect 15151 23681 15163 23715
rect 18598 23712 18604 23724
rect 18559 23684 18604 23712
rect 15105 23675 15163 23681
rect 18598 23672 18604 23684
rect 18656 23672 18662 23724
rect 20530 23672 20536 23724
rect 20588 23712 20594 23724
rect 22005 23715 22063 23721
rect 22005 23712 22017 23715
rect 20588 23684 22017 23712
rect 20588 23672 20594 23684
rect 22005 23681 22017 23684
rect 22051 23681 22063 23715
rect 22005 23675 22063 23681
rect 26142 23672 26148 23724
rect 26200 23712 26206 23724
rect 26421 23715 26479 23721
rect 26421 23712 26433 23715
rect 26200 23684 26433 23712
rect 26200 23672 26206 23684
rect 26421 23681 26433 23684
rect 26467 23681 26479 23715
rect 26421 23675 26479 23681
rect 27356 23656 27384 23752
rect 27430 23672 27436 23724
rect 27488 23712 27494 23724
rect 27488 23684 27533 23712
rect 27488 23672 27494 23684
rect 6546 23644 6552 23656
rect 6507 23616 6552 23644
rect 6546 23604 6552 23616
rect 6604 23604 6610 23656
rect 14550 23644 14556 23656
rect 14511 23616 14556 23644
rect 14550 23604 14556 23616
rect 14608 23604 14614 23656
rect 19610 23604 19616 23656
rect 19668 23644 19674 23656
rect 20625 23647 20683 23653
rect 20625 23644 20637 23647
rect 19668 23616 20637 23644
rect 19668 23604 19674 23616
rect 20625 23613 20637 23616
rect 20671 23613 20683 23647
rect 27338 23644 27344 23656
rect 27299 23616 27344 23644
rect 20625 23607 20683 23613
rect 27338 23604 27344 23616
rect 27396 23604 27402 23656
rect 27982 23604 27988 23656
rect 28040 23644 28046 23656
rect 28169 23647 28227 23653
rect 28169 23644 28181 23647
rect 28040 23616 28181 23644
rect 28040 23604 28046 23616
rect 28169 23613 28181 23616
rect 28215 23613 28227 23647
rect 28169 23607 28227 23613
rect 26513 23511 26571 23517
rect 26513 23477 26525 23511
rect 26559 23508 26571 23511
rect 26694 23508 26700 23520
rect 26559 23480 26700 23508
rect 26559 23477 26571 23480
rect 26513 23471 26571 23477
rect 26694 23468 26700 23480
rect 26752 23468 26758 23520
rect 1104 23418 28888 23440
rect 1104 23366 4423 23418
rect 4475 23366 4487 23418
rect 4539 23366 4551 23418
rect 4603 23366 4615 23418
rect 4667 23366 4679 23418
rect 4731 23366 11369 23418
rect 11421 23366 11433 23418
rect 11485 23366 11497 23418
rect 11549 23366 11561 23418
rect 11613 23366 11625 23418
rect 11677 23366 18315 23418
rect 18367 23366 18379 23418
rect 18431 23366 18443 23418
rect 18495 23366 18507 23418
rect 18559 23366 18571 23418
rect 18623 23366 25261 23418
rect 25313 23366 25325 23418
rect 25377 23366 25389 23418
rect 25441 23366 25453 23418
rect 25505 23366 25517 23418
rect 25569 23366 28888 23418
rect 1104 23344 28888 23366
rect 3329 23307 3387 23313
rect 3329 23273 3341 23307
rect 3375 23304 3387 23307
rect 4062 23304 4068 23316
rect 3375 23276 4068 23304
rect 3375 23273 3387 23276
rect 3329 23267 3387 23273
rect 4062 23264 4068 23276
rect 4120 23264 4126 23316
rect 11149 23307 11207 23313
rect 11149 23273 11161 23307
rect 11195 23304 11207 23307
rect 12526 23304 12532 23316
rect 11195 23276 12532 23304
rect 11195 23273 11207 23276
rect 11149 23267 11207 23273
rect 12526 23264 12532 23276
rect 12584 23264 12590 23316
rect 14277 23307 14335 23313
rect 14277 23273 14289 23307
rect 14323 23304 14335 23307
rect 14366 23304 14372 23316
rect 14323 23276 14372 23304
rect 14323 23273 14335 23276
rect 14277 23267 14335 23273
rect 14366 23264 14372 23276
rect 14424 23264 14430 23316
rect 25130 23304 25136 23316
rect 25091 23276 25136 23304
rect 25130 23264 25136 23276
rect 25188 23264 25194 23316
rect 26142 23264 26148 23316
rect 26200 23304 26206 23316
rect 28169 23307 28227 23313
rect 28169 23304 28181 23307
rect 26200 23276 28181 23304
rect 26200 23264 26234 23276
rect 28169 23273 28181 23276
rect 28215 23273 28227 23307
rect 28169 23267 28227 23273
rect 2774 23236 2780 23248
rect 2332 23208 2780 23236
rect 2222 23060 2228 23112
rect 2280 23100 2286 23112
rect 2332 23109 2360 23208
rect 2774 23196 2780 23208
rect 2832 23196 2838 23248
rect 23477 23239 23535 23245
rect 23477 23205 23489 23239
rect 23523 23236 23535 23239
rect 23658 23236 23664 23248
rect 23523 23208 23664 23236
rect 23523 23205 23535 23208
rect 23477 23199 23535 23205
rect 23658 23196 23664 23208
rect 23716 23196 23722 23248
rect 26206 23236 26234 23264
rect 23860 23208 26234 23236
rect 2409 23171 2467 23177
rect 2409 23137 2421 23171
rect 2455 23168 2467 23171
rect 6638 23168 6644 23180
rect 2455 23140 3188 23168
rect 2455 23137 2467 23140
rect 2409 23131 2467 23137
rect 2317 23103 2375 23109
rect 2317 23100 2329 23103
rect 2280 23072 2329 23100
rect 2280 23060 2286 23072
rect 2317 23069 2329 23072
rect 2363 23069 2375 23103
rect 2317 23063 2375 23069
rect 2501 23103 2559 23109
rect 2501 23069 2513 23103
rect 2547 23100 2559 23103
rect 3050 23100 3056 23112
rect 2547 23072 3056 23100
rect 2547 23069 2559 23072
rect 2501 23063 2559 23069
rect 3050 23060 3056 23072
rect 3108 23060 3114 23112
rect 3160 23109 3188 23140
rect 6288 23140 6644 23168
rect 3145 23103 3203 23109
rect 3145 23069 3157 23103
rect 3191 23069 3203 23103
rect 3145 23063 3203 23069
rect 3418 23060 3424 23112
rect 3476 23100 3482 23112
rect 3970 23100 3976 23112
rect 3476 23072 3521 23100
rect 3931 23072 3976 23100
rect 3476 23060 3482 23072
rect 3970 23060 3976 23072
rect 4028 23060 4034 23112
rect 5810 23060 5816 23112
rect 5868 23100 5874 23112
rect 6288 23109 6316 23140
rect 6638 23128 6644 23140
rect 6696 23128 6702 23180
rect 7282 23168 7288 23180
rect 7243 23140 7288 23168
rect 7282 23128 7288 23140
rect 7340 23128 7346 23180
rect 8113 23171 8171 23177
rect 8113 23137 8125 23171
rect 8159 23168 8171 23171
rect 8202 23168 8208 23180
rect 8159 23140 8208 23168
rect 8159 23137 8171 23140
rect 8113 23131 8171 23137
rect 8202 23128 8208 23140
rect 8260 23128 8266 23180
rect 8389 23171 8447 23177
rect 8389 23137 8401 23171
rect 8435 23168 8447 23171
rect 9766 23168 9772 23180
rect 8435 23140 9772 23168
rect 8435 23137 8447 23140
rect 8389 23131 8447 23137
rect 9766 23128 9772 23140
rect 9824 23128 9830 23180
rect 10502 23128 10508 23180
rect 10560 23168 10566 23180
rect 10689 23171 10747 23177
rect 10689 23168 10701 23171
rect 10560 23140 10701 23168
rect 10560 23128 10566 23140
rect 10689 23137 10701 23140
rect 10735 23137 10747 23171
rect 12618 23168 12624 23180
rect 10689 23131 10747 23137
rect 12268 23140 12624 23168
rect 6273 23103 6331 23109
rect 6273 23100 6285 23103
rect 5868 23072 6285 23100
rect 5868 23060 5874 23072
rect 6273 23069 6285 23072
rect 6319 23069 6331 23103
rect 6273 23063 6331 23069
rect 6454 23060 6460 23112
rect 6512 23060 6518 23112
rect 7834 23060 7840 23112
rect 7892 23100 7898 23112
rect 12268 23109 12296 23140
rect 12618 23128 12624 23140
rect 12676 23168 12682 23180
rect 13170 23168 13176 23180
rect 12676 23140 13176 23168
rect 12676 23128 12682 23140
rect 13170 23128 13176 23140
rect 13228 23128 13234 23180
rect 14734 23168 14740 23180
rect 14695 23140 14740 23168
rect 14734 23128 14740 23140
rect 14792 23128 14798 23180
rect 14829 23171 14887 23177
rect 14829 23137 14841 23171
rect 14875 23137 14887 23171
rect 14829 23131 14887 23137
rect 8021 23103 8079 23109
rect 8021 23100 8033 23103
rect 7892 23072 8033 23100
rect 7892 23060 7898 23072
rect 8021 23069 8033 23072
rect 8067 23069 8079 23103
rect 8021 23063 8079 23069
rect 10781 23103 10839 23109
rect 10781 23069 10793 23103
rect 10827 23069 10839 23103
rect 10781 23063 10839 23069
rect 12253 23103 12311 23109
rect 12253 23069 12265 23103
rect 12299 23069 12311 23103
rect 12253 23063 12311 23069
rect 12437 23103 12495 23109
rect 12437 23069 12449 23103
rect 12483 23100 12495 23103
rect 12802 23100 12808 23112
rect 12483 23072 12808 23100
rect 12483 23069 12495 23072
rect 12437 23063 12495 23069
rect 2774 22924 2780 22976
rect 2832 22964 2838 22976
rect 2961 22967 3019 22973
rect 2961 22964 2973 22967
rect 2832 22936 2973 22964
rect 2832 22924 2838 22936
rect 2961 22933 2973 22936
rect 3007 22933 3019 22967
rect 2961 22927 3019 22933
rect 4338 22924 4344 22976
rect 4396 22964 4402 22976
rect 5261 22967 5319 22973
rect 5261 22964 5273 22967
rect 4396 22936 5273 22964
rect 4396 22924 4402 22936
rect 5261 22933 5273 22936
rect 5307 22933 5319 22967
rect 5261 22927 5319 22933
rect 6362 22924 6368 22976
rect 6420 22964 6426 22976
rect 6730 22964 6736 22976
rect 6420 22936 6736 22964
rect 6420 22924 6426 22936
rect 6730 22924 6736 22936
rect 6788 22964 6794 22976
rect 10796 22964 10824 23063
rect 12802 23060 12808 23072
rect 12860 23060 12866 23112
rect 14642 23060 14648 23112
rect 14700 23100 14706 23112
rect 14844 23100 14872 23131
rect 23566 23128 23572 23180
rect 23624 23168 23630 23180
rect 23753 23171 23811 23177
rect 23753 23168 23765 23171
rect 23624 23140 23765 23168
rect 23624 23128 23630 23140
rect 23753 23137 23765 23140
rect 23799 23137 23811 23171
rect 23753 23131 23811 23137
rect 15654 23100 15660 23112
rect 14700 23072 14872 23100
rect 15615 23072 15660 23100
rect 14700 23060 14706 23072
rect 15654 23060 15660 23072
rect 15712 23060 15718 23112
rect 23860 23109 23888 23208
rect 24026 23128 24032 23180
rect 24084 23168 24090 23180
rect 24673 23171 24731 23177
rect 24673 23168 24685 23171
rect 24084 23140 24685 23168
rect 24084 23128 24090 23140
rect 24673 23137 24685 23140
rect 24719 23137 24731 23171
rect 26694 23168 26700 23180
rect 26655 23140 26700 23168
rect 24673 23131 24731 23137
rect 26694 23128 26700 23140
rect 26752 23128 26758 23180
rect 23845 23103 23903 23109
rect 23845 23069 23857 23103
rect 23891 23069 23903 23103
rect 23845 23063 23903 23069
rect 24765 23103 24823 23109
rect 24765 23069 24777 23103
rect 24811 23100 24823 23103
rect 26234 23100 26240 23112
rect 24811 23072 26240 23100
rect 24811 23069 24823 23072
rect 24765 23063 24823 23069
rect 26234 23060 26240 23072
rect 26292 23060 26298 23112
rect 26418 23100 26424 23112
rect 26379 23072 26424 23100
rect 26418 23060 26424 23072
rect 26476 23060 26482 23112
rect 19794 22992 19800 23044
rect 19852 23032 19858 23044
rect 20809 23035 20867 23041
rect 20809 23032 20821 23035
rect 19852 23004 20821 23032
rect 19852 22992 19858 23004
rect 20809 23001 20821 23004
rect 20855 23001 20867 23035
rect 22554 23032 22560 23044
rect 22515 23004 22560 23032
rect 20809 22995 20867 23001
rect 22554 22992 22560 23004
rect 22612 22992 22618 23044
rect 27982 23032 27988 23044
rect 27922 23004 27988 23032
rect 27982 22992 27988 23004
rect 28040 22992 28046 23044
rect 12250 22964 12256 22976
rect 6788 22936 10824 22964
rect 12211 22936 12256 22964
rect 6788 22924 6794 22936
rect 12250 22924 12256 22936
rect 12308 22924 12314 22976
rect 14090 22924 14096 22976
rect 14148 22964 14154 22976
rect 14550 22964 14556 22976
rect 14148 22936 14556 22964
rect 14148 22924 14154 22936
rect 14550 22924 14556 22936
rect 14608 22964 14614 22976
rect 14645 22967 14703 22973
rect 14645 22964 14657 22967
rect 14608 22936 14657 22964
rect 14608 22924 14614 22936
rect 14645 22933 14657 22936
rect 14691 22933 14703 22967
rect 14645 22927 14703 22933
rect 15565 22967 15623 22973
rect 15565 22933 15577 22967
rect 15611 22964 15623 22967
rect 16206 22964 16212 22976
rect 15611 22936 16212 22964
rect 15611 22933 15623 22936
rect 15565 22927 15623 22933
rect 16206 22924 16212 22936
rect 16264 22924 16270 22976
rect 1104 22874 29048 22896
rect 1104 22822 7896 22874
rect 7948 22822 7960 22874
rect 8012 22822 8024 22874
rect 8076 22822 8088 22874
rect 8140 22822 8152 22874
rect 8204 22822 14842 22874
rect 14894 22822 14906 22874
rect 14958 22822 14970 22874
rect 15022 22822 15034 22874
rect 15086 22822 15098 22874
rect 15150 22822 21788 22874
rect 21840 22822 21852 22874
rect 21904 22822 21916 22874
rect 21968 22822 21980 22874
rect 22032 22822 22044 22874
rect 22096 22822 28734 22874
rect 28786 22822 28798 22874
rect 28850 22822 28862 22874
rect 28914 22822 28926 22874
rect 28978 22822 28990 22874
rect 29042 22822 29048 22874
rect 1104 22800 29048 22822
rect 4154 22720 4160 22772
rect 4212 22760 4218 22772
rect 4265 22763 4323 22769
rect 4265 22760 4277 22763
rect 4212 22732 4277 22760
rect 4212 22720 4218 22732
rect 4265 22729 4277 22732
rect 4311 22729 4323 22763
rect 4265 22723 4323 22729
rect 5353 22763 5411 22769
rect 5353 22729 5365 22763
rect 5399 22760 5411 22763
rect 6546 22760 6552 22772
rect 5399 22732 6552 22760
rect 5399 22729 5411 22732
rect 5353 22723 5411 22729
rect 6546 22720 6552 22732
rect 6604 22720 6610 22772
rect 8294 22720 8300 22772
rect 8352 22760 8358 22772
rect 8481 22763 8539 22769
rect 8481 22760 8493 22763
rect 8352 22732 8493 22760
rect 8352 22720 8358 22732
rect 8481 22729 8493 22732
rect 8527 22729 8539 22763
rect 16942 22760 16948 22772
rect 8481 22723 8539 22729
rect 13648 22732 16948 22760
rect 3418 22652 3424 22704
rect 3476 22692 3482 22704
rect 4065 22695 4123 22701
rect 4065 22692 4077 22695
rect 3476 22664 4077 22692
rect 3476 22652 3482 22664
rect 4065 22661 4077 22664
rect 4111 22661 4123 22695
rect 4065 22655 4123 22661
rect 7300 22664 9444 22692
rect 2492 22627 2550 22633
rect 2492 22593 2504 22627
rect 2538 22624 2550 22627
rect 3694 22624 3700 22636
rect 2538 22596 3700 22624
rect 2538 22593 2550 22596
rect 2492 22587 2550 22593
rect 3694 22584 3700 22596
rect 3752 22584 3758 22636
rect 4246 22584 4252 22636
rect 4304 22584 4310 22636
rect 5445 22627 5503 22633
rect 5445 22593 5457 22627
rect 5491 22624 5503 22627
rect 6362 22624 6368 22636
rect 5491 22596 6368 22624
rect 5491 22593 5503 22596
rect 5445 22587 5503 22593
rect 6362 22584 6368 22596
rect 6420 22584 6426 22636
rect 7098 22624 7104 22636
rect 7011 22596 7104 22624
rect 7098 22584 7104 22596
rect 7156 22624 7162 22636
rect 7300 22624 7328 22664
rect 9416 22636 9444 22664
rect 11054 22652 11060 22704
rect 11112 22692 11118 22704
rect 11977 22695 12035 22701
rect 11977 22692 11989 22695
rect 11112 22664 11989 22692
rect 11112 22652 11118 22664
rect 11977 22661 11989 22664
rect 12023 22661 12035 22695
rect 11977 22655 12035 22661
rect 12069 22695 12127 22701
rect 12069 22661 12081 22695
rect 12115 22692 12127 22695
rect 12434 22692 12440 22704
rect 12115 22664 12440 22692
rect 12115 22661 12127 22664
rect 12069 22655 12127 22661
rect 12434 22652 12440 22664
rect 12492 22652 12498 22704
rect 7156 22596 7328 22624
rect 7368 22627 7426 22633
rect 7156 22584 7162 22596
rect 7368 22593 7380 22627
rect 7414 22624 7426 22627
rect 7650 22624 7656 22636
rect 7414 22596 7656 22624
rect 7414 22593 7426 22596
rect 7368 22587 7426 22593
rect 7650 22584 7656 22596
rect 7708 22584 7714 22636
rect 9398 22624 9404 22636
rect 9359 22596 9404 22624
rect 9398 22584 9404 22596
rect 9456 22584 9462 22636
rect 9674 22633 9680 22636
rect 9668 22587 9680 22633
rect 9732 22624 9738 22636
rect 9732 22596 9768 22624
rect 9674 22584 9680 22587
rect 9732 22584 9738 22596
rect 11146 22584 11152 22636
rect 11204 22624 11210 22636
rect 11839 22627 11897 22633
rect 11839 22624 11851 22627
rect 11204 22596 11851 22624
rect 11204 22584 11210 22596
rect 11839 22593 11851 22596
rect 11885 22593 11897 22627
rect 12250 22624 12256 22636
rect 12211 22596 12256 22624
rect 11839 22587 11897 22593
rect 12250 22584 12256 22596
rect 12308 22584 12314 22636
rect 13648 22633 13676 22732
rect 16942 22720 16948 22732
rect 17000 22720 17006 22772
rect 19426 22760 19432 22772
rect 19387 22732 19432 22760
rect 19426 22720 19432 22732
rect 19484 22720 19490 22772
rect 22554 22720 22560 22772
rect 22612 22760 22618 22772
rect 23382 22760 23388 22772
rect 22612 22732 23388 22760
rect 22612 22720 22618 22732
rect 23382 22720 23388 22732
rect 23440 22760 23446 22772
rect 23937 22763 23995 22769
rect 23937 22760 23949 22763
rect 23440 22732 23949 22760
rect 23440 22720 23446 22732
rect 23937 22729 23949 22732
rect 23983 22729 23995 22763
rect 23937 22723 23995 22729
rect 26418 22720 26424 22772
rect 26476 22760 26482 22772
rect 26513 22763 26571 22769
rect 26513 22760 26525 22763
rect 26476 22732 26525 22760
rect 26476 22720 26482 22732
rect 26513 22729 26525 22732
rect 26559 22729 26571 22763
rect 26513 22723 26571 22729
rect 15286 22652 15292 22704
rect 15344 22652 15350 22704
rect 12345 22627 12403 22633
rect 12345 22593 12357 22627
rect 12391 22593 12403 22627
rect 12345 22587 12403 22593
rect 13633 22627 13691 22633
rect 13633 22593 13645 22627
rect 13679 22593 13691 22627
rect 13633 22587 13691 22593
rect 2038 22516 2044 22568
rect 2096 22556 2102 22568
rect 2225 22559 2283 22565
rect 2225 22556 2237 22559
rect 2096 22528 2237 22556
rect 2096 22516 2102 22528
rect 2225 22525 2237 22528
rect 2271 22525 2283 22559
rect 2225 22519 2283 22525
rect 4264 22488 4292 22584
rect 11238 22516 11244 22568
rect 11296 22556 11302 22568
rect 12360 22556 12388 22587
rect 16206 22584 16212 22636
rect 16264 22624 16270 22636
rect 16264 22596 16309 22624
rect 16264 22584 16270 22596
rect 17770 22584 17776 22636
rect 17828 22624 17834 22636
rect 17865 22627 17923 22633
rect 17865 22624 17877 22627
rect 17828 22596 17877 22624
rect 17828 22584 17834 22596
rect 17865 22593 17877 22596
rect 17911 22593 17923 22627
rect 19794 22624 19800 22636
rect 19755 22596 19800 22624
rect 17865 22587 17923 22593
rect 19794 22584 19800 22596
rect 19852 22584 19858 22636
rect 19886 22584 19892 22636
rect 19944 22624 19950 22636
rect 20073 22627 20131 22633
rect 20073 22624 20085 22627
rect 19944 22596 20085 22624
rect 19944 22584 19950 22596
rect 20073 22593 20085 22596
rect 20119 22593 20131 22627
rect 22646 22624 22652 22636
rect 22607 22596 22652 22624
rect 20073 22587 20131 22593
rect 22646 22584 22652 22596
rect 22704 22584 22710 22636
rect 26234 22584 26240 22636
rect 26292 22624 26298 22636
rect 26605 22627 26663 22633
rect 26605 22624 26617 22627
rect 26292 22596 26617 22624
rect 26292 22584 26298 22596
rect 26605 22593 26617 22596
rect 26651 22624 26663 22627
rect 27341 22627 27399 22633
rect 27341 22624 27353 22627
rect 26651 22596 27353 22624
rect 26651 22593 26663 22596
rect 26605 22587 26663 22593
rect 27341 22593 27353 22596
rect 27387 22624 27399 22627
rect 27522 22624 27528 22636
rect 27387 22596 27528 22624
rect 27387 22593 27399 22596
rect 27341 22587 27399 22593
rect 27522 22584 27528 22596
rect 27580 22584 27586 22636
rect 13354 22556 13360 22568
rect 11296 22528 12388 22556
rect 13315 22528 13360 22556
rect 11296 22516 11302 22528
rect 13354 22516 13360 22528
rect 13412 22516 13418 22568
rect 14182 22556 14188 22568
rect 14143 22528 14188 22556
rect 14182 22516 14188 22528
rect 14240 22516 14246 22568
rect 15930 22556 15936 22568
rect 15891 22528 15936 22556
rect 15930 22516 15936 22528
rect 15988 22516 15994 22568
rect 17954 22556 17960 22568
rect 17915 22528 17960 22556
rect 17954 22516 17960 22528
rect 18012 22516 18018 22568
rect 18049 22559 18107 22565
rect 18049 22525 18061 22559
rect 18095 22525 18107 22559
rect 18049 22519 18107 22525
rect 4433 22491 4491 22497
rect 4433 22488 4445 22491
rect 4264 22460 4445 22488
rect 4433 22457 4445 22460
rect 4479 22488 4491 22491
rect 4798 22488 4804 22500
rect 4479 22460 4804 22488
rect 4479 22457 4491 22460
rect 4433 22451 4491 22457
rect 4798 22448 4804 22460
rect 4856 22448 4862 22500
rect 17678 22448 17684 22500
rect 17736 22488 17742 22500
rect 17862 22488 17868 22500
rect 17736 22460 17868 22488
rect 17736 22448 17742 22460
rect 17862 22448 17868 22460
rect 17920 22488 17926 22500
rect 18064 22488 18092 22519
rect 17920 22460 18092 22488
rect 17920 22448 17926 22460
rect 3605 22423 3663 22429
rect 3605 22389 3617 22423
rect 3651 22420 3663 22423
rect 4154 22420 4160 22432
rect 3651 22392 4160 22420
rect 3651 22389 3663 22392
rect 3605 22383 3663 22389
rect 4154 22380 4160 22392
rect 4212 22420 4218 22432
rect 4249 22423 4307 22429
rect 4249 22420 4261 22423
rect 4212 22392 4261 22420
rect 4212 22380 4218 22392
rect 4249 22389 4261 22392
rect 4295 22389 4307 22423
rect 4249 22383 4307 22389
rect 10781 22423 10839 22429
rect 10781 22389 10793 22423
rect 10827 22420 10839 22423
rect 10962 22420 10968 22432
rect 10827 22392 10968 22420
rect 10827 22389 10839 22392
rect 10781 22383 10839 22389
rect 10962 22380 10968 22392
rect 11020 22380 11026 22432
rect 11701 22423 11759 22429
rect 11701 22389 11713 22423
rect 11747 22420 11759 22423
rect 11974 22420 11980 22432
rect 11747 22392 11980 22420
rect 11747 22389 11759 22392
rect 11701 22383 11759 22389
rect 11974 22380 11980 22392
rect 12032 22380 12038 22432
rect 17494 22420 17500 22432
rect 17455 22392 17500 22420
rect 17494 22380 17500 22392
rect 17552 22380 17558 22432
rect 27246 22420 27252 22432
rect 27207 22392 27252 22420
rect 27246 22380 27252 22392
rect 27304 22380 27310 22432
rect 1104 22330 28888 22352
rect 1104 22278 4423 22330
rect 4475 22278 4487 22330
rect 4539 22278 4551 22330
rect 4603 22278 4615 22330
rect 4667 22278 4679 22330
rect 4731 22278 11369 22330
rect 11421 22278 11433 22330
rect 11485 22278 11497 22330
rect 11549 22278 11561 22330
rect 11613 22278 11625 22330
rect 11677 22278 18315 22330
rect 18367 22278 18379 22330
rect 18431 22278 18443 22330
rect 18495 22278 18507 22330
rect 18559 22278 18571 22330
rect 18623 22278 25261 22330
rect 25313 22278 25325 22330
rect 25377 22278 25389 22330
rect 25441 22278 25453 22330
rect 25505 22278 25517 22330
rect 25569 22278 28888 22330
rect 1104 22256 28888 22278
rect 3418 22216 3424 22228
rect 3379 22188 3424 22216
rect 3418 22176 3424 22188
rect 3476 22176 3482 22228
rect 7650 22216 7656 22228
rect 7611 22188 7656 22216
rect 7650 22176 7656 22188
rect 7708 22176 7714 22228
rect 17954 22176 17960 22228
rect 18012 22216 18018 22228
rect 18601 22219 18659 22225
rect 18601 22216 18613 22219
rect 18012 22188 18613 22216
rect 18012 22176 18018 22188
rect 18601 22185 18613 22188
rect 18647 22185 18659 22219
rect 24026 22216 24032 22228
rect 23987 22188 24032 22216
rect 18601 22179 18659 22185
rect 3436 22080 3464 22176
rect 7742 22108 7748 22160
rect 7800 22148 7806 22160
rect 10410 22148 10416 22160
rect 7800 22120 10416 22148
rect 7800 22108 7806 22120
rect 4341 22083 4399 22089
rect 4341 22080 4353 22083
rect 3436 22052 4353 22080
rect 4341 22049 4353 22052
rect 4387 22049 4399 22083
rect 6454 22080 6460 22092
rect 4341 22043 4399 22049
rect 5828 22052 6460 22080
rect 5828 22024 5856 22052
rect 6454 22040 6460 22052
rect 6512 22040 6518 22092
rect 8113 22083 8171 22089
rect 8113 22049 8125 22083
rect 8159 22080 8171 22083
rect 8202 22080 8208 22092
rect 8159 22052 8208 22080
rect 8159 22049 8171 22052
rect 8113 22043 8171 22049
rect 8202 22040 8208 22052
rect 8260 22040 8266 22092
rect 8312 22089 8340 22120
rect 10410 22108 10416 22120
rect 10468 22108 10474 22160
rect 8297 22083 8355 22089
rect 8297 22049 8309 22083
rect 8343 22080 8355 22083
rect 8343 22052 8377 22080
rect 8343 22049 8355 22052
rect 8297 22043 8355 22049
rect 12434 22040 12440 22092
rect 12492 22080 12498 22092
rect 15286 22080 15292 22092
rect 12492 22052 12537 22080
rect 15247 22052 15292 22080
rect 12492 22040 12498 22052
rect 15286 22040 15292 22052
rect 15344 22040 15350 22092
rect 18616 22080 18644 22179
rect 24026 22176 24032 22188
rect 24084 22176 24090 22228
rect 26500 22219 26558 22225
rect 26500 22185 26512 22219
rect 26546 22216 26558 22219
rect 27246 22216 27252 22228
rect 26546 22188 27252 22216
rect 26546 22185 26558 22188
rect 26500 22179 26558 22185
rect 27246 22176 27252 22188
rect 27304 22176 27310 22228
rect 19521 22083 19579 22089
rect 19521 22080 19533 22083
rect 18616 22052 19533 22080
rect 19521 22049 19533 22052
rect 19567 22049 19579 22083
rect 19978 22080 19984 22092
rect 19939 22052 19984 22080
rect 19521 22043 19579 22049
rect 19978 22040 19984 22052
rect 20036 22040 20042 22092
rect 27522 22040 27528 22092
rect 27580 22080 27586 22092
rect 27985 22083 28043 22089
rect 27985 22080 27997 22083
rect 27580 22052 27997 22080
rect 27580 22040 27586 22052
rect 27985 22049 27997 22052
rect 28031 22049 28043 22083
rect 27985 22043 28043 22049
rect 14464 22024 14516 22030
rect 2038 22012 2044 22024
rect 1999 21984 2044 22012
rect 2038 21972 2044 21984
rect 2096 21972 2102 22024
rect 2308 22015 2366 22021
rect 2308 21981 2320 22015
rect 2354 22012 2366 22015
rect 2774 22012 2780 22024
rect 2354 21984 2780 22012
rect 2354 21981 2366 21984
rect 2308 21975 2366 21981
rect 2774 21972 2780 21984
rect 2832 21972 2838 22024
rect 3050 21972 3056 22024
rect 3108 22012 3114 22024
rect 3973 22015 4031 22021
rect 3973 22012 3985 22015
rect 3108 21984 3985 22012
rect 3108 21972 3114 21984
rect 3973 21981 3985 21984
rect 4019 22012 4031 22015
rect 4062 22012 4068 22024
rect 4019 21984 4068 22012
rect 4019 21981 4031 21984
rect 3973 21975 4031 21981
rect 4062 21972 4068 21984
rect 4120 21972 4126 22024
rect 4157 22015 4215 22021
rect 4157 21981 4169 22015
rect 4203 22012 4215 22015
rect 4246 22012 4252 22024
rect 4203 21984 4252 22012
rect 4203 21981 4215 21984
rect 4157 21975 4215 21981
rect 4246 21972 4252 21984
rect 4304 21972 4310 22024
rect 5534 21972 5540 22024
rect 5592 22012 5598 22024
rect 5629 22015 5687 22021
rect 5629 22012 5641 22015
rect 5592 21984 5641 22012
rect 5592 21972 5598 21984
rect 5629 21981 5641 21984
rect 5675 21981 5687 22015
rect 5629 21975 5687 21981
rect 5810 21972 5816 22024
rect 5868 21972 5874 22024
rect 10410 21972 10416 22024
rect 10468 22012 10474 22024
rect 12250 22012 12256 22024
rect 10468 21984 12256 22012
rect 10468 21972 10474 21984
rect 12250 21972 12256 21984
rect 12308 21972 12314 22024
rect 12618 22012 12624 22024
rect 12579 21984 12624 22012
rect 12618 21972 12624 21984
rect 12676 21972 12682 22024
rect 12802 22012 12808 22024
rect 12763 21984 12808 22012
rect 12802 21972 12808 21984
rect 12860 21972 12866 22024
rect 13262 22012 13268 22024
rect 13223 21984 13268 22012
rect 13262 21972 13268 21984
rect 13320 21972 13326 22024
rect 14369 22015 14427 22021
rect 14369 21981 14381 22015
rect 14415 21981 14427 22015
rect 14369 21975 14427 21981
rect 6362 21944 6368 21956
rect 6323 21916 6368 21944
rect 6362 21904 6368 21916
rect 6420 21904 6426 21956
rect 9582 21904 9588 21956
rect 9640 21944 9646 21956
rect 10229 21947 10287 21953
rect 10229 21944 10241 21947
rect 9640 21916 10241 21944
rect 9640 21904 9646 21916
rect 10229 21913 10241 21916
rect 10275 21913 10287 21947
rect 10229 21907 10287 21913
rect 11977 21947 12035 21953
rect 11977 21913 11989 21947
rect 12023 21944 12035 21947
rect 12526 21944 12532 21956
rect 12023 21916 12532 21944
rect 12023 21913 12035 21916
rect 11977 21907 12035 21913
rect 12526 21904 12532 21916
rect 12584 21904 12590 21956
rect 13538 21944 13544 21956
rect 13499 21916 13544 21944
rect 13538 21904 13544 21916
rect 13596 21904 13602 21956
rect 8021 21879 8079 21885
rect 8021 21845 8033 21879
rect 8067 21876 8079 21879
rect 9398 21876 9404 21888
rect 8067 21848 9404 21876
rect 8067 21845 8079 21848
rect 8021 21839 8079 21845
rect 9398 21836 9404 21848
rect 9456 21836 9462 21888
rect 9858 21836 9864 21888
rect 9916 21876 9922 21888
rect 14384 21876 14412 21975
rect 16850 21972 16856 22024
rect 16908 22012 16914 22024
rect 17221 22015 17279 22021
rect 17221 22012 17233 22015
rect 16908 21984 17233 22012
rect 16908 21972 16914 21984
rect 17221 21981 17233 21984
rect 17267 22012 17279 22015
rect 17310 22012 17316 22024
rect 17267 21984 17316 22012
rect 17267 21981 17279 21984
rect 17221 21975 17279 21981
rect 17310 21972 17316 21984
rect 17368 21972 17374 22024
rect 17494 22021 17500 22024
rect 17488 21975 17500 22021
rect 17552 22012 17558 22024
rect 19610 22012 19616 22024
rect 17552 21984 17588 22012
rect 19571 21984 19616 22012
rect 17494 21972 17500 21975
rect 17552 21972 17558 21984
rect 19610 21972 19616 21984
rect 19668 21972 19674 22024
rect 22649 22015 22707 22021
rect 22649 21981 22661 22015
rect 22695 22012 22707 22015
rect 22738 22012 22744 22024
rect 22695 21984 22744 22012
rect 22695 21981 22707 21984
rect 22649 21975 22707 21981
rect 22738 21972 22744 21984
rect 22796 21972 22802 22024
rect 26234 22012 26240 22024
rect 26195 21984 26240 22012
rect 26234 21972 26240 21984
rect 26292 21972 26298 22024
rect 14464 21966 14516 21972
rect 22916 21947 22974 21953
rect 22916 21913 22928 21947
rect 22962 21944 22974 21947
rect 23198 21944 23204 21956
rect 22962 21916 23204 21944
rect 22962 21913 22974 21916
rect 22916 21907 22974 21913
rect 23198 21904 23204 21916
rect 23256 21904 23262 21956
rect 28258 21944 28264 21956
rect 27738 21916 28264 21944
rect 28258 21904 28264 21916
rect 28316 21904 28322 21956
rect 9916 21848 14412 21876
rect 9916 21836 9922 21848
rect 1104 21786 29048 21808
rect 1104 21734 7896 21786
rect 7948 21734 7960 21786
rect 8012 21734 8024 21786
rect 8076 21734 8088 21786
rect 8140 21734 8152 21786
rect 8204 21734 14842 21786
rect 14894 21734 14906 21786
rect 14958 21734 14970 21786
rect 15022 21734 15034 21786
rect 15086 21734 15098 21786
rect 15150 21734 21788 21786
rect 21840 21734 21852 21786
rect 21904 21734 21916 21786
rect 21968 21734 21980 21786
rect 22032 21734 22044 21786
rect 22096 21734 28734 21786
rect 28786 21734 28798 21786
rect 28850 21734 28862 21786
rect 28914 21734 28926 21786
rect 28978 21734 28990 21786
rect 29042 21734 29048 21786
rect 1104 21712 29048 21734
rect 3694 21672 3700 21684
rect 2746 21644 3280 21672
rect 3655 21644 3700 21672
rect 2222 21604 2228 21616
rect 2135 21576 2228 21604
rect 2148 21545 2176 21576
rect 2222 21564 2228 21576
rect 2280 21604 2286 21616
rect 2746 21604 2774 21644
rect 3142 21604 3148 21616
rect 2280 21576 2774 21604
rect 2884 21576 3148 21604
rect 2280 21564 2286 21576
rect 2133 21539 2191 21545
rect 2133 21505 2145 21539
rect 2179 21505 2191 21539
rect 2133 21499 2191 21505
rect 2317 21539 2375 21545
rect 2317 21505 2329 21539
rect 2363 21536 2375 21539
rect 2884 21536 2912 21576
rect 3142 21564 3148 21576
rect 3200 21564 3206 21616
rect 3252 21604 3280 21644
rect 3694 21632 3700 21644
rect 3752 21632 3758 21684
rect 9674 21632 9680 21684
rect 9732 21672 9738 21684
rect 9769 21675 9827 21681
rect 9769 21672 9781 21675
rect 9732 21644 9781 21672
rect 9732 21632 9738 21644
rect 9769 21641 9781 21644
rect 9815 21641 9827 21675
rect 9769 21635 9827 21641
rect 10134 21632 10140 21684
rect 10192 21632 10198 21684
rect 11146 21672 11152 21684
rect 11107 21644 11152 21672
rect 11146 21632 11152 21644
rect 11204 21632 11210 21684
rect 12802 21632 12808 21684
rect 12860 21672 12866 21684
rect 13446 21672 13452 21684
rect 12860 21644 13452 21672
rect 12860 21632 12866 21644
rect 13446 21632 13452 21644
rect 13504 21672 13510 21684
rect 13725 21675 13783 21681
rect 13725 21672 13737 21675
rect 13504 21644 13737 21672
rect 13504 21632 13510 21644
rect 13725 21641 13737 21644
rect 13771 21641 13783 21675
rect 13725 21635 13783 21641
rect 15381 21675 15439 21681
rect 15381 21641 15393 21675
rect 15427 21672 15439 21675
rect 15930 21672 15936 21684
rect 15427 21644 15936 21672
rect 15427 21641 15439 21644
rect 15381 21635 15439 21641
rect 15930 21632 15936 21644
rect 15988 21632 15994 21684
rect 21542 21672 21548 21684
rect 16040 21644 21548 21672
rect 4798 21604 4804 21616
rect 3252 21576 4804 21604
rect 4798 21564 4804 21576
rect 4856 21564 4862 21616
rect 10152 21604 10180 21632
rect 10870 21604 10876 21616
rect 10152 21576 10876 21604
rect 10870 21564 10876 21576
rect 10928 21604 10934 21616
rect 10928 21576 11192 21604
rect 10928 21564 10934 21576
rect 2363 21508 2912 21536
rect 2961 21539 3019 21545
rect 2363 21505 2375 21508
rect 2317 21499 2375 21505
rect 2961 21505 2973 21539
rect 3007 21505 3019 21539
rect 3878 21536 3884 21548
rect 3839 21508 3884 21536
rect 2961 21499 3019 21505
rect 2225 21471 2283 21477
rect 2225 21437 2237 21471
rect 2271 21468 2283 21471
rect 2976 21468 3004 21499
rect 3878 21496 3884 21508
rect 3936 21496 3942 21548
rect 4154 21536 4160 21548
rect 4115 21508 4160 21536
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 6730 21536 6736 21548
rect 6691 21508 6736 21536
rect 6730 21496 6736 21508
rect 6788 21496 6794 21548
rect 10134 21536 10140 21548
rect 10095 21508 10140 21536
rect 10134 21496 10140 21508
rect 10192 21496 10198 21548
rect 10229 21539 10287 21545
rect 10229 21505 10241 21539
rect 10275 21536 10287 21539
rect 10686 21536 10692 21548
rect 10275 21508 10692 21536
rect 10275 21505 10287 21508
rect 10229 21499 10287 21505
rect 10686 21496 10692 21508
rect 10744 21536 10750 21548
rect 10962 21536 10968 21548
rect 10744 21508 10968 21536
rect 10744 21496 10750 21508
rect 10962 21496 10968 21508
rect 11020 21496 11026 21548
rect 11164 21545 11192 21576
rect 13538 21564 13544 21616
rect 13596 21604 13602 21616
rect 16040 21604 16068 21644
rect 21542 21632 21548 21644
rect 21600 21672 21606 21684
rect 22738 21672 22744 21684
rect 21600 21644 22744 21672
rect 21600 21632 21606 21644
rect 22738 21632 22744 21644
rect 22796 21632 22802 21684
rect 23198 21672 23204 21684
rect 23159 21644 23204 21672
rect 23198 21632 23204 21644
rect 23256 21632 23262 21684
rect 23661 21675 23719 21681
rect 23661 21641 23673 21675
rect 23707 21672 23719 21675
rect 24026 21672 24032 21684
rect 23707 21644 24032 21672
rect 23707 21641 23719 21644
rect 23661 21635 23719 21641
rect 24026 21632 24032 21644
rect 24084 21632 24090 21684
rect 26234 21632 26240 21684
rect 26292 21672 26298 21684
rect 26329 21675 26387 21681
rect 26329 21672 26341 21675
rect 26292 21644 26341 21672
rect 26292 21632 26298 21644
rect 26329 21641 26341 21644
rect 26375 21641 26387 21675
rect 28258 21672 28264 21684
rect 28219 21644 28264 21672
rect 26329 21635 26387 21641
rect 28258 21632 28264 21644
rect 28316 21632 28322 21684
rect 17310 21604 17316 21616
rect 13596 21576 16068 21604
rect 16960 21576 17316 21604
rect 13596 21564 13602 21576
rect 11149 21539 11207 21545
rect 11149 21505 11161 21539
rect 11195 21505 11207 21539
rect 11149 21499 11207 21505
rect 12612 21539 12670 21545
rect 12612 21505 12624 21539
rect 12658 21536 12670 21539
rect 12986 21536 12992 21548
rect 12658 21508 12992 21536
rect 12658 21505 12670 21508
rect 12612 21499 12670 21505
rect 12986 21496 12992 21508
rect 13044 21496 13050 21548
rect 14182 21496 14188 21548
rect 14240 21536 14246 21548
rect 16960 21545 16988 21576
rect 17310 21564 17316 21576
rect 17368 21604 17374 21616
rect 17494 21604 17500 21616
rect 17368 21576 17500 21604
rect 17368 21564 17374 21576
rect 17494 21564 17500 21576
rect 17552 21564 17558 21616
rect 23474 21564 23480 21616
rect 23532 21604 23538 21616
rect 23569 21607 23627 21613
rect 23569 21604 23581 21607
rect 23532 21576 23581 21604
rect 23532 21564 23538 21576
rect 23569 21573 23581 21576
rect 23615 21604 23627 21607
rect 23750 21604 23756 21616
rect 23615 21576 23756 21604
rect 23615 21573 23627 21576
rect 23569 21567 23627 21573
rect 23750 21564 23756 21576
rect 23808 21564 23814 21616
rect 17218 21545 17224 21548
rect 14645 21539 14703 21545
rect 14645 21536 14657 21539
rect 14240 21508 14657 21536
rect 14240 21496 14246 21508
rect 14645 21505 14657 21508
rect 14691 21536 14703 21539
rect 15289 21539 15347 21545
rect 15289 21536 15301 21539
rect 14691 21508 15301 21536
rect 14691 21505 14703 21508
rect 14645 21499 14703 21505
rect 15289 21505 15301 21508
rect 15335 21505 15347 21539
rect 15289 21499 15347 21505
rect 16945 21539 17003 21545
rect 16945 21505 16957 21539
rect 16991 21505 17003 21539
rect 16945 21499 17003 21505
rect 17212 21499 17224 21545
rect 17276 21536 17282 21548
rect 19245 21539 19303 21545
rect 17276 21508 17312 21536
rect 17218 21496 17224 21499
rect 17276 21496 17282 21508
rect 19245 21505 19257 21539
rect 19291 21536 19303 21539
rect 19702 21536 19708 21548
rect 19291 21508 19708 21536
rect 19291 21505 19303 21508
rect 19245 21499 19303 21505
rect 19702 21496 19708 21508
rect 19760 21496 19766 21548
rect 21634 21496 21640 21548
rect 21692 21536 21698 21548
rect 22005 21539 22063 21545
rect 22005 21536 22017 21539
rect 21692 21508 22017 21536
rect 21692 21496 21698 21508
rect 22005 21505 22017 21508
rect 22051 21505 22063 21539
rect 22005 21499 22063 21505
rect 22189 21539 22247 21545
rect 22189 21505 22201 21539
rect 22235 21536 22247 21539
rect 22830 21536 22836 21548
rect 22235 21508 22836 21536
rect 22235 21505 22247 21508
rect 22189 21499 22247 21505
rect 22830 21496 22836 21508
rect 22888 21496 22894 21548
rect 24765 21539 24823 21545
rect 24765 21505 24777 21539
rect 24811 21536 24823 21539
rect 26418 21536 26424 21548
rect 24811 21508 26424 21536
rect 24811 21505 24823 21508
rect 24765 21499 24823 21505
rect 26418 21496 26424 21508
rect 26476 21496 26482 21548
rect 27430 21536 27436 21548
rect 27391 21508 27436 21536
rect 27430 21496 27436 21508
rect 27488 21496 27494 21548
rect 3234 21468 3240 21480
rect 2271 21440 3004 21468
rect 3195 21440 3240 21468
rect 2271 21437 2283 21440
rect 2225 21431 2283 21437
rect 3234 21428 3240 21440
rect 3292 21428 3298 21480
rect 4062 21468 4068 21480
rect 4023 21440 4068 21468
rect 4062 21428 4068 21440
rect 4120 21428 4126 21480
rect 10410 21468 10416 21480
rect 10371 21440 10416 21468
rect 10410 21428 10416 21440
rect 10468 21428 10474 21480
rect 12342 21468 12348 21480
rect 12303 21440 12348 21468
rect 12342 21428 12348 21440
rect 12400 21428 12406 21480
rect 14734 21468 14740 21480
rect 14695 21440 14740 21468
rect 14734 21428 14740 21440
rect 14792 21428 14798 21480
rect 19153 21471 19211 21477
rect 19153 21468 19165 21471
rect 18340 21440 19165 21468
rect 17954 21360 17960 21412
rect 18012 21400 18018 21412
rect 18340 21409 18368 21440
rect 19153 21437 19165 21440
rect 19199 21437 19211 21471
rect 19153 21431 19211 21437
rect 23845 21471 23903 21477
rect 23845 21437 23857 21471
rect 23891 21468 23903 21471
rect 24673 21471 24731 21477
rect 23891 21440 24532 21468
rect 23891 21437 23903 21440
rect 23845 21431 23903 21437
rect 18325 21403 18383 21409
rect 18325 21400 18337 21403
rect 18012 21372 18337 21400
rect 18012 21360 18018 21372
rect 18325 21369 18337 21372
rect 18371 21369 18383 21403
rect 18325 21363 18383 21369
rect 2774 21292 2780 21344
rect 2832 21332 2838 21344
rect 3145 21335 3203 21341
rect 2832 21304 2877 21332
rect 2832 21292 2838 21304
rect 3145 21301 3157 21335
rect 3191 21332 3203 21335
rect 4890 21332 4896 21344
rect 3191 21304 4896 21332
rect 3191 21301 3203 21304
rect 3145 21295 3203 21301
rect 4890 21292 4896 21304
rect 4948 21292 4954 21344
rect 5626 21292 5632 21344
rect 5684 21332 5690 21344
rect 6641 21335 6699 21341
rect 6641 21332 6653 21335
rect 5684 21304 6653 21332
rect 5684 21292 5690 21304
rect 6641 21301 6653 21304
rect 6687 21301 6699 21335
rect 6641 21295 6699 21301
rect 12250 21292 12256 21344
rect 12308 21332 12314 21344
rect 12710 21332 12716 21344
rect 12308 21304 12716 21332
rect 12308 21292 12314 21304
rect 12710 21292 12716 21304
rect 12768 21292 12774 21344
rect 13814 21292 13820 21344
rect 13872 21332 13878 21344
rect 14277 21335 14335 21341
rect 14277 21332 14289 21335
rect 13872 21304 14289 21332
rect 13872 21292 13878 21304
rect 14277 21301 14289 21304
rect 14323 21301 14335 21335
rect 14277 21295 14335 21301
rect 19613 21335 19671 21341
rect 19613 21301 19625 21335
rect 19659 21332 19671 21335
rect 21818 21332 21824 21344
rect 19659 21304 21824 21332
rect 19659 21301 19671 21304
rect 19613 21295 19671 21301
rect 21818 21292 21824 21304
rect 21876 21292 21882 21344
rect 22097 21335 22155 21341
rect 22097 21301 22109 21335
rect 22143 21332 22155 21335
rect 22278 21332 22284 21344
rect 22143 21304 22284 21332
rect 22143 21301 22155 21304
rect 22097 21295 22155 21301
rect 22278 21292 22284 21304
rect 22336 21292 22342 21344
rect 23566 21292 23572 21344
rect 23624 21332 23630 21344
rect 24397 21335 24455 21341
rect 24397 21332 24409 21335
rect 23624 21304 24409 21332
rect 23624 21292 23630 21304
rect 24397 21301 24409 21304
rect 24443 21301 24455 21335
rect 24504 21332 24532 21440
rect 24673 21437 24685 21471
rect 24719 21437 24731 21471
rect 24673 21431 24731 21437
rect 24688 21400 24716 21431
rect 26234 21428 26240 21480
rect 26292 21468 26298 21480
rect 27338 21468 27344 21480
rect 26292 21440 27344 21468
rect 26292 21428 26298 21440
rect 27338 21428 27344 21440
rect 27396 21428 27402 21480
rect 24762 21400 24768 21412
rect 24688 21372 24768 21400
rect 24762 21360 24768 21372
rect 24820 21360 24826 21412
rect 25130 21332 25136 21344
rect 24504 21304 25136 21332
rect 24397 21295 24455 21301
rect 25130 21292 25136 21304
rect 25188 21292 25194 21344
rect 1104 21242 28888 21264
rect 1104 21190 4423 21242
rect 4475 21190 4487 21242
rect 4539 21190 4551 21242
rect 4603 21190 4615 21242
rect 4667 21190 4679 21242
rect 4731 21190 11369 21242
rect 11421 21190 11433 21242
rect 11485 21190 11497 21242
rect 11549 21190 11561 21242
rect 11613 21190 11625 21242
rect 11677 21190 18315 21242
rect 18367 21190 18379 21242
rect 18431 21190 18443 21242
rect 18495 21190 18507 21242
rect 18559 21190 18571 21242
rect 18623 21190 25261 21242
rect 25313 21190 25325 21242
rect 25377 21190 25389 21242
rect 25441 21190 25453 21242
rect 25505 21190 25517 21242
rect 25569 21190 28888 21242
rect 1104 21168 28888 21190
rect 6730 21088 6736 21140
rect 6788 21128 6794 21140
rect 7101 21131 7159 21137
rect 7101 21128 7113 21131
rect 6788 21100 7113 21128
rect 6788 21088 6794 21100
rect 7101 21097 7113 21100
rect 7147 21097 7159 21131
rect 7101 21091 7159 21097
rect 9398 21088 9404 21140
rect 9456 21128 9462 21140
rect 12986 21128 12992 21140
rect 9456 21100 12848 21128
rect 12947 21100 12992 21128
rect 9456 21088 9462 21100
rect 12820 21060 12848 21100
rect 12986 21088 12992 21100
rect 13044 21088 13050 21140
rect 13354 21088 13360 21140
rect 13412 21128 13418 21140
rect 15930 21128 15936 21140
rect 13412 21100 15936 21128
rect 13412 21088 13418 21100
rect 15930 21088 15936 21100
rect 15988 21088 15994 21140
rect 17218 21088 17224 21140
rect 17276 21128 17282 21140
rect 17313 21131 17371 21137
rect 17313 21128 17325 21131
rect 17276 21100 17325 21128
rect 17276 21088 17282 21100
rect 17313 21097 17325 21100
rect 17359 21097 17371 21131
rect 17313 21091 17371 21097
rect 19978 21088 19984 21140
rect 20036 21128 20042 21140
rect 23569 21131 23627 21137
rect 23569 21128 23581 21131
rect 20036 21100 23581 21128
rect 20036 21088 20042 21100
rect 23569 21097 23581 21100
rect 23615 21097 23627 21131
rect 23569 21091 23627 21097
rect 16758 21060 16764 21072
rect 12820 21032 16764 21060
rect 16758 21020 16764 21032
rect 16816 21060 16822 21072
rect 17126 21060 17132 21072
rect 16816 21032 17132 21060
rect 16816 21020 16822 21032
rect 17126 21020 17132 21032
rect 17184 21020 17190 21072
rect 24029 21063 24087 21069
rect 24029 21029 24041 21063
rect 24075 21029 24087 21063
rect 24029 21023 24087 21029
rect 5353 20995 5411 21001
rect 5353 20961 5365 20995
rect 5399 20992 5411 20995
rect 5718 20992 5724 21004
rect 5399 20964 5724 20992
rect 5399 20961 5411 20964
rect 5353 20955 5411 20961
rect 5718 20952 5724 20964
rect 5776 20952 5782 21004
rect 7742 20952 7748 21004
rect 7800 20992 7806 21004
rect 7929 20995 7987 21001
rect 7929 20992 7941 20995
rect 7800 20964 7941 20992
rect 7800 20952 7806 20964
rect 7929 20961 7941 20964
rect 7975 20961 7987 20995
rect 7929 20955 7987 20961
rect 8389 20995 8447 21001
rect 8389 20961 8401 20995
rect 8435 20992 8447 20995
rect 9674 20992 9680 21004
rect 8435 20964 9680 20992
rect 8435 20961 8447 20964
rect 8389 20955 8447 20961
rect 9674 20952 9680 20964
rect 9732 20952 9738 21004
rect 12161 20995 12219 21001
rect 12161 20961 12173 20995
rect 12207 20992 12219 20995
rect 13446 20992 13452 21004
rect 12207 20964 13308 20992
rect 13407 20964 13452 20992
rect 12207 20961 12219 20964
rect 12161 20955 12219 20961
rect 3329 20927 3387 20933
rect 3329 20893 3341 20927
rect 3375 20924 3387 20927
rect 4338 20924 4344 20936
rect 3375 20896 4344 20924
rect 3375 20893 3387 20896
rect 3329 20887 3387 20893
rect 4338 20884 4344 20896
rect 4396 20884 4402 20936
rect 7650 20884 7656 20936
rect 7708 20924 7714 20936
rect 8021 20927 8079 20933
rect 8021 20924 8033 20927
rect 7708 20896 8033 20924
rect 7708 20884 7714 20896
rect 8021 20893 8033 20896
rect 8067 20893 8079 20927
rect 8021 20887 8079 20893
rect 10134 20884 10140 20936
rect 10192 20924 10198 20936
rect 13280 20924 13308 20964
rect 13446 20952 13452 20964
rect 13504 20952 13510 21004
rect 13633 20995 13691 21001
rect 13633 20961 13645 20995
rect 13679 20992 13691 20995
rect 14642 20992 14648 21004
rect 13679 20964 14648 20992
rect 13679 20961 13691 20964
rect 13633 20955 13691 20961
rect 14642 20952 14648 20964
rect 14700 20992 14706 21004
rect 14829 20995 14887 21001
rect 14829 20992 14841 20995
rect 14700 20964 14841 20992
rect 14700 20952 14706 20964
rect 14829 20961 14841 20964
rect 14875 20961 14887 20995
rect 17862 20992 17868 21004
rect 17823 20964 17868 20992
rect 14829 20955 14887 20961
rect 17862 20952 17868 20964
rect 17920 20952 17926 21004
rect 23658 20992 23664 21004
rect 23619 20964 23664 20992
rect 23658 20952 23664 20964
rect 23716 20952 23722 21004
rect 14458 20924 14464 20936
rect 10192 20896 12756 20924
rect 13280 20896 14464 20924
rect 10192 20884 10198 20896
rect 5626 20856 5632 20868
rect 5587 20828 5632 20856
rect 5626 20816 5632 20828
rect 5684 20816 5690 20868
rect 6362 20816 6368 20868
rect 6420 20816 6426 20868
rect 9582 20816 9588 20868
rect 9640 20856 9646 20868
rect 10413 20859 10471 20865
rect 10413 20856 10425 20859
rect 9640 20828 10425 20856
rect 9640 20816 9646 20828
rect 10413 20825 10425 20828
rect 10459 20825 10471 20859
rect 12728 20856 12756 20896
rect 14458 20884 14464 20896
rect 14516 20884 14522 20936
rect 17126 20884 17132 20936
rect 17184 20924 17190 20936
rect 17681 20927 17739 20933
rect 17681 20924 17693 20927
rect 17184 20896 17693 20924
rect 17184 20884 17190 20896
rect 17681 20893 17693 20896
rect 17727 20893 17739 20927
rect 17681 20887 17739 20893
rect 17773 20927 17831 20933
rect 17773 20893 17785 20927
rect 17819 20924 17831 20927
rect 17954 20924 17960 20936
rect 17819 20896 17960 20924
rect 17819 20893 17831 20896
rect 17773 20887 17831 20893
rect 17954 20884 17960 20896
rect 18012 20884 18018 20936
rect 19981 20927 20039 20933
rect 19981 20893 19993 20927
rect 20027 20924 20039 20927
rect 20070 20924 20076 20936
rect 20027 20896 20076 20924
rect 20027 20893 20039 20896
rect 19981 20887 20039 20893
rect 20070 20884 20076 20896
rect 20128 20924 20134 20936
rect 20530 20924 20536 20936
rect 20128 20896 20536 20924
rect 20128 20884 20134 20896
rect 20530 20884 20536 20896
rect 20588 20884 20594 20936
rect 21818 20924 21824 20936
rect 21779 20896 21824 20924
rect 21818 20884 21824 20896
rect 21876 20884 21882 20936
rect 21914 20927 21972 20933
rect 21914 20893 21926 20927
rect 21960 20893 21972 20927
rect 21914 20887 21972 20893
rect 14550 20856 14556 20868
rect 12728 20828 14556 20856
rect 10413 20819 10471 20825
rect 14550 20816 14556 20828
rect 14608 20856 14614 20868
rect 14645 20859 14703 20865
rect 14645 20856 14657 20859
rect 14608 20828 14657 20856
rect 14608 20816 14614 20828
rect 14645 20825 14657 20828
rect 14691 20825 14703 20859
rect 14645 20819 14703 20825
rect 20248 20859 20306 20865
rect 20248 20825 20260 20859
rect 20294 20856 20306 20859
rect 20438 20856 20444 20868
rect 20294 20828 20444 20856
rect 20294 20825 20306 20828
rect 20248 20819 20306 20825
rect 20438 20816 20444 20828
rect 20496 20816 20502 20868
rect 21266 20816 21272 20868
rect 21324 20856 21330 20868
rect 21928 20856 21956 20887
rect 22094 20884 22100 20936
rect 22152 20924 22158 20936
rect 22152 20896 22197 20924
rect 22152 20884 22158 20896
rect 22278 20884 22284 20936
rect 22336 20933 22342 20936
rect 22336 20924 22344 20933
rect 23566 20924 23572 20936
rect 22336 20896 22381 20924
rect 23527 20896 23572 20924
rect 22336 20887 22344 20896
rect 22336 20884 22342 20887
rect 23566 20884 23572 20896
rect 23624 20884 23630 20936
rect 23842 20924 23848 20936
rect 23803 20896 23848 20924
rect 23842 20884 23848 20896
rect 23900 20884 23906 20936
rect 24044 20924 24072 21023
rect 24670 20952 24676 21004
rect 24728 20992 24734 21004
rect 25041 20995 25099 21001
rect 25041 20992 25053 20995
rect 24728 20964 25053 20992
rect 24728 20952 24734 20964
rect 25041 20961 25053 20964
rect 25087 20961 25099 20995
rect 25041 20955 25099 20961
rect 24581 20927 24639 20933
rect 24581 20924 24593 20927
rect 24044 20896 24593 20924
rect 24581 20893 24593 20896
rect 24627 20893 24639 20927
rect 24581 20887 24639 20893
rect 24857 20927 24915 20933
rect 24857 20893 24869 20927
rect 24903 20893 24915 20927
rect 27890 20924 27896 20936
rect 27851 20896 27896 20924
rect 24857 20887 24915 20893
rect 21324 20828 21956 20856
rect 22189 20859 22247 20865
rect 21324 20816 21330 20828
rect 22189 20825 22201 20859
rect 22235 20856 22247 20859
rect 22370 20856 22376 20868
rect 22235 20828 22376 20856
rect 22235 20825 22247 20828
rect 22189 20819 22247 20825
rect 22370 20816 22376 20828
rect 22428 20816 22434 20868
rect 24872 20856 24900 20887
rect 27890 20884 27896 20896
rect 27948 20884 27954 20936
rect 28166 20856 28172 20868
rect 22480 20828 24900 20856
rect 28127 20828 28172 20856
rect 2038 20788 2044 20800
rect 1999 20760 2044 20788
rect 2038 20748 2044 20760
rect 2096 20748 2102 20800
rect 13354 20788 13360 20800
rect 13315 20760 13360 20788
rect 13354 20748 13360 20760
rect 13412 20748 13418 20800
rect 14274 20788 14280 20800
rect 14235 20760 14280 20788
rect 14274 20748 14280 20760
rect 14332 20748 14338 20800
rect 14734 20748 14740 20800
rect 14792 20788 14798 20800
rect 21361 20791 21419 20797
rect 14792 20760 14837 20788
rect 14792 20748 14798 20760
rect 21361 20757 21373 20791
rect 21407 20788 21419 20791
rect 21634 20788 21640 20800
rect 21407 20760 21640 20788
rect 21407 20757 21419 20760
rect 21361 20751 21419 20757
rect 21634 20748 21640 20760
rect 21692 20748 21698 20800
rect 22480 20797 22508 20828
rect 28166 20816 28172 20828
rect 28224 20816 28230 20868
rect 22465 20791 22523 20797
rect 22465 20757 22477 20791
rect 22511 20757 22523 20791
rect 24854 20788 24860 20800
rect 24815 20760 24860 20788
rect 22465 20751 22523 20757
rect 24854 20748 24860 20760
rect 24912 20748 24918 20800
rect 1104 20698 29048 20720
rect 1104 20646 7896 20698
rect 7948 20646 7960 20698
rect 8012 20646 8024 20698
rect 8076 20646 8088 20698
rect 8140 20646 8152 20698
rect 8204 20646 14842 20698
rect 14894 20646 14906 20698
rect 14958 20646 14970 20698
rect 15022 20646 15034 20698
rect 15086 20646 15098 20698
rect 15150 20646 21788 20698
rect 21840 20646 21852 20698
rect 21904 20646 21916 20698
rect 21968 20646 21980 20698
rect 22032 20646 22044 20698
rect 22096 20646 28734 20698
rect 28786 20646 28798 20698
rect 28850 20646 28862 20698
rect 28914 20646 28926 20698
rect 28978 20646 28990 20698
rect 29042 20646 29048 20698
rect 1104 20624 29048 20646
rect 3234 20544 3240 20596
rect 3292 20584 3298 20596
rect 3421 20587 3479 20593
rect 3421 20584 3433 20587
rect 3292 20556 3433 20584
rect 3292 20544 3298 20556
rect 3421 20553 3433 20556
rect 3467 20553 3479 20587
rect 3421 20547 3479 20553
rect 2308 20519 2366 20525
rect 2308 20485 2320 20519
rect 2354 20516 2366 20519
rect 2774 20516 2780 20528
rect 2354 20488 2780 20516
rect 2354 20485 2366 20488
rect 2308 20479 2366 20485
rect 2774 20476 2780 20488
rect 2832 20476 2838 20528
rect 3436 20516 3464 20547
rect 5718 20544 5724 20596
rect 5776 20584 5782 20596
rect 5813 20587 5871 20593
rect 5813 20584 5825 20587
rect 5776 20556 5825 20584
rect 5776 20544 5782 20556
rect 5813 20553 5825 20556
rect 5859 20553 5871 20587
rect 5813 20547 5871 20553
rect 8205 20587 8263 20593
rect 8205 20553 8217 20587
rect 8251 20584 8263 20587
rect 10134 20584 10140 20596
rect 8251 20556 10140 20584
rect 8251 20553 8263 20556
rect 8205 20547 8263 20553
rect 10134 20544 10140 20556
rect 10192 20544 10198 20596
rect 11054 20584 11060 20596
rect 11015 20556 11060 20584
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 14734 20544 14740 20596
rect 14792 20584 14798 20596
rect 15105 20587 15163 20593
rect 15105 20584 15117 20587
rect 14792 20556 15117 20584
rect 14792 20544 14798 20556
rect 15105 20553 15117 20556
rect 15151 20553 15163 20587
rect 20438 20584 20444 20596
rect 20399 20556 20444 20584
rect 15105 20547 15163 20553
rect 20438 20544 20444 20556
rect 20496 20544 20502 20596
rect 22370 20584 22376 20596
rect 22331 20556 22376 20584
rect 22370 20544 22376 20556
rect 22428 20544 22434 20596
rect 9585 20519 9643 20525
rect 3436 20488 4844 20516
rect 4246 20408 4252 20460
rect 4304 20448 4310 20460
rect 4816 20457 4844 20488
rect 9585 20485 9597 20519
rect 9631 20516 9643 20519
rect 13814 20516 13820 20528
rect 9631 20488 13820 20516
rect 9631 20485 9643 20488
rect 9585 20479 9643 20485
rect 13814 20476 13820 20488
rect 13872 20476 13878 20528
rect 13992 20519 14050 20525
rect 13992 20485 14004 20519
rect 14038 20516 14050 20519
rect 14274 20516 14280 20528
rect 14038 20488 14280 20516
rect 14038 20485 14050 20488
rect 13992 20479 14050 20485
rect 14274 20476 14280 20488
rect 14332 20476 14338 20528
rect 17126 20525 17132 20528
rect 17120 20516 17132 20525
rect 17087 20488 17132 20516
rect 17120 20479 17132 20488
rect 17126 20476 17132 20479
rect 17184 20476 17190 20528
rect 17770 20476 17776 20528
rect 17828 20516 17834 20528
rect 20809 20519 20867 20525
rect 20809 20516 20821 20519
rect 17828 20488 20821 20516
rect 17828 20476 17834 20488
rect 20809 20485 20821 20488
rect 20855 20485 20867 20519
rect 20809 20479 20867 20485
rect 20901 20519 20959 20525
rect 20901 20485 20913 20519
rect 20947 20516 20959 20519
rect 21634 20516 21640 20528
rect 20947 20488 21640 20516
rect 20947 20485 20959 20488
rect 20901 20479 20959 20485
rect 4341 20451 4399 20457
rect 4341 20448 4353 20451
rect 4304 20420 4353 20448
rect 4304 20408 4310 20420
rect 4341 20417 4353 20420
rect 4387 20417 4399 20451
rect 4341 20411 4399 20417
rect 4801 20451 4859 20457
rect 4801 20417 4813 20451
rect 4847 20417 4859 20451
rect 4801 20411 4859 20417
rect 4890 20408 4896 20460
rect 4948 20448 4954 20460
rect 4985 20451 5043 20457
rect 4985 20448 4997 20451
rect 4948 20420 4997 20448
rect 4948 20408 4954 20420
rect 4985 20417 4997 20420
rect 5031 20417 5043 20451
rect 4985 20411 5043 20417
rect 5905 20451 5963 20457
rect 5905 20417 5917 20451
rect 5951 20448 5963 20451
rect 5994 20448 6000 20460
rect 5951 20420 6000 20448
rect 5951 20417 5963 20420
rect 5905 20411 5963 20417
rect 5994 20408 6000 20420
rect 6052 20448 6058 20460
rect 7650 20448 7656 20460
rect 6052 20420 7656 20448
rect 6052 20408 6058 20420
rect 7650 20408 7656 20420
rect 7708 20408 7714 20460
rect 9858 20448 9864 20460
rect 9819 20420 9864 20448
rect 9858 20408 9864 20420
rect 9916 20408 9922 20460
rect 10686 20448 10692 20460
rect 10647 20420 10692 20448
rect 10686 20408 10692 20420
rect 10744 20408 10750 20460
rect 10870 20448 10876 20460
rect 10831 20420 10876 20448
rect 10870 20408 10876 20420
rect 10928 20408 10934 20460
rect 11701 20451 11759 20457
rect 11701 20417 11713 20451
rect 11747 20417 11759 20451
rect 11974 20448 11980 20460
rect 11935 20420 11980 20448
rect 11701 20411 11759 20417
rect 2038 20380 2044 20392
rect 1999 20352 2044 20380
rect 2038 20340 2044 20352
rect 2096 20340 2102 20392
rect 3234 20340 3240 20392
rect 3292 20380 3298 20392
rect 4157 20383 4215 20389
rect 4157 20380 4169 20383
rect 3292 20352 4169 20380
rect 3292 20340 3298 20352
rect 4157 20349 4169 20352
rect 4203 20380 4215 20383
rect 7098 20380 7104 20392
rect 4203 20352 7104 20380
rect 4203 20349 4215 20352
rect 4157 20343 4215 20349
rect 7098 20340 7104 20352
rect 7156 20340 7162 20392
rect 7742 20340 7748 20392
rect 7800 20380 7806 20392
rect 8297 20383 8355 20389
rect 8297 20380 8309 20383
rect 7800 20352 8309 20380
rect 7800 20340 7806 20352
rect 8297 20349 8309 20352
rect 8343 20349 8355 20383
rect 8297 20343 8355 20349
rect 8481 20383 8539 20389
rect 8481 20349 8493 20383
rect 8527 20380 8539 20383
rect 9398 20380 9404 20392
rect 8527 20352 9404 20380
rect 8527 20349 8539 20352
rect 8481 20343 8539 20349
rect 9398 20340 9404 20352
rect 9456 20340 9462 20392
rect 9766 20380 9772 20392
rect 9727 20352 9772 20380
rect 9766 20340 9772 20352
rect 9824 20340 9830 20392
rect 11716 20380 11744 20411
rect 11974 20408 11980 20420
rect 12032 20408 12038 20460
rect 12158 20448 12164 20460
rect 12119 20420 12164 20448
rect 12158 20408 12164 20420
rect 12216 20408 12222 20460
rect 12805 20451 12863 20457
rect 12805 20417 12817 20451
rect 12851 20448 12863 20451
rect 13538 20448 13544 20460
rect 12851 20420 13544 20448
rect 12851 20417 12863 20420
rect 12805 20411 12863 20417
rect 13538 20408 13544 20420
rect 13596 20408 13602 20460
rect 20824 20448 20852 20479
rect 21634 20476 21640 20488
rect 21692 20516 21698 20528
rect 22005 20519 22063 20525
rect 22005 20516 22017 20519
rect 21692 20488 22017 20516
rect 21692 20476 21698 20488
rect 22005 20485 22017 20488
rect 22051 20485 22063 20519
rect 22005 20479 22063 20485
rect 22189 20519 22247 20525
rect 22189 20485 22201 20519
rect 22235 20516 22247 20519
rect 22830 20516 22836 20528
rect 22235 20488 22836 20516
rect 22235 20485 22247 20488
rect 22189 20479 22247 20485
rect 22830 20476 22836 20488
rect 22888 20476 22894 20528
rect 23382 20516 23388 20528
rect 23343 20488 23388 20516
rect 23382 20476 23388 20488
rect 23440 20476 23446 20528
rect 24946 20448 24952 20460
rect 20824 20420 24952 20448
rect 24946 20408 24952 20420
rect 25004 20408 25010 20460
rect 26418 20408 26424 20460
rect 26476 20448 26482 20460
rect 27338 20448 27344 20460
rect 26476 20420 27344 20448
rect 26476 20408 26482 20420
rect 27338 20408 27344 20420
rect 27396 20408 27402 20460
rect 10060 20352 11744 20380
rect 12345 20383 12403 20389
rect 10060 20321 10088 20352
rect 12345 20349 12357 20383
rect 12391 20349 12403 20383
rect 12345 20343 12403 20349
rect 13081 20383 13139 20389
rect 13081 20349 13093 20383
rect 13127 20380 13139 20383
rect 13630 20380 13636 20392
rect 13127 20352 13636 20380
rect 13127 20349 13139 20352
rect 13081 20343 13139 20349
rect 10045 20315 10103 20321
rect 10045 20281 10057 20315
rect 10091 20281 10103 20315
rect 12360 20312 12388 20343
rect 13630 20340 13636 20352
rect 13688 20380 13694 20392
rect 13725 20383 13783 20389
rect 13725 20380 13737 20383
rect 13688 20352 13737 20380
rect 13688 20340 13694 20352
rect 13725 20349 13737 20352
rect 13771 20349 13783 20383
rect 16850 20380 16856 20392
rect 16811 20352 16856 20380
rect 13725 20343 13783 20349
rect 16850 20340 16856 20352
rect 16908 20340 16914 20392
rect 20993 20383 21051 20389
rect 20993 20380 21005 20383
rect 18156 20352 21005 20380
rect 13170 20312 13176 20324
rect 12360 20284 13176 20312
rect 10045 20275 10103 20281
rect 13170 20272 13176 20284
rect 13228 20272 13234 20324
rect 3142 20204 3148 20256
rect 3200 20244 3206 20256
rect 5169 20247 5227 20253
rect 5169 20244 5181 20247
rect 3200 20216 5181 20244
rect 3200 20204 3206 20216
rect 5169 20213 5181 20216
rect 5215 20213 5227 20247
rect 5169 20207 5227 20213
rect 7558 20204 7564 20256
rect 7616 20244 7622 20256
rect 7837 20247 7895 20253
rect 7837 20244 7849 20247
rect 7616 20216 7849 20244
rect 7616 20204 7622 20216
rect 7837 20213 7849 20216
rect 7883 20213 7895 20247
rect 9674 20244 9680 20256
rect 9635 20216 9680 20244
rect 7837 20207 7895 20213
rect 9674 20204 9680 20216
rect 9732 20204 9738 20256
rect 16758 20204 16764 20256
rect 16816 20244 16822 20256
rect 18156 20244 18184 20352
rect 20993 20349 21005 20352
rect 21039 20380 21051 20383
rect 22462 20380 22468 20392
rect 21039 20352 22468 20380
rect 21039 20349 21051 20352
rect 20993 20343 21051 20349
rect 22462 20340 22468 20352
rect 22520 20340 22526 20392
rect 25133 20383 25191 20389
rect 25133 20349 25145 20383
rect 25179 20380 25191 20383
rect 26234 20380 26240 20392
rect 25179 20352 26240 20380
rect 25179 20349 25191 20352
rect 25133 20343 25191 20349
rect 26234 20340 26240 20352
rect 26292 20340 26298 20392
rect 18233 20315 18291 20321
rect 18233 20281 18245 20315
rect 18279 20312 18291 20315
rect 27614 20312 27620 20324
rect 18279 20284 27620 20312
rect 18279 20281 18291 20284
rect 18233 20275 18291 20281
rect 27614 20272 27620 20284
rect 27672 20272 27678 20324
rect 16816 20216 18184 20244
rect 16816 20204 16822 20216
rect 26786 20204 26792 20256
rect 26844 20244 26850 20256
rect 27249 20247 27307 20253
rect 27249 20244 27261 20247
rect 26844 20216 27261 20244
rect 26844 20204 26850 20216
rect 27249 20213 27261 20216
rect 27295 20213 27307 20247
rect 27249 20207 27307 20213
rect 1104 20154 28888 20176
rect 1104 20102 4423 20154
rect 4475 20102 4487 20154
rect 4539 20102 4551 20154
rect 4603 20102 4615 20154
rect 4667 20102 4679 20154
rect 4731 20102 11369 20154
rect 11421 20102 11433 20154
rect 11485 20102 11497 20154
rect 11549 20102 11561 20154
rect 11613 20102 11625 20154
rect 11677 20102 18315 20154
rect 18367 20102 18379 20154
rect 18431 20102 18443 20154
rect 18495 20102 18507 20154
rect 18559 20102 18571 20154
rect 18623 20102 25261 20154
rect 25313 20102 25325 20154
rect 25377 20102 25389 20154
rect 25441 20102 25453 20154
rect 25505 20102 25517 20154
rect 25569 20102 28888 20154
rect 1104 20080 28888 20102
rect 7650 20000 7656 20052
rect 7708 20040 7714 20052
rect 8481 20043 8539 20049
rect 8481 20040 8493 20043
rect 7708 20012 8493 20040
rect 7708 20000 7714 20012
rect 8481 20009 8493 20012
rect 8527 20009 8539 20043
rect 8481 20003 8539 20009
rect 9677 20043 9735 20049
rect 9677 20009 9689 20043
rect 9723 20040 9735 20043
rect 9858 20040 9864 20052
rect 9723 20012 9864 20040
rect 9723 20009 9735 20012
rect 9677 20003 9735 20009
rect 9858 20000 9864 20012
rect 9916 20000 9922 20052
rect 10502 20040 10508 20052
rect 10463 20012 10508 20040
rect 10502 20000 10508 20012
rect 10560 20040 10566 20052
rect 12158 20040 12164 20052
rect 10560 20012 12164 20040
rect 10560 20000 10566 20012
rect 12158 20000 12164 20012
rect 12216 20000 12222 20052
rect 17681 20043 17739 20049
rect 17681 20009 17693 20043
rect 17727 20040 17739 20043
rect 17862 20040 17868 20052
rect 17727 20012 17868 20040
rect 17727 20009 17739 20012
rect 17681 20003 17739 20009
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 20070 20040 20076 20052
rect 20031 20012 20076 20040
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 21266 20040 21272 20052
rect 21227 20012 21272 20040
rect 21266 20000 21272 20012
rect 21324 20000 21330 20052
rect 27338 20000 27344 20052
rect 27396 20040 27402 20052
rect 28261 20043 28319 20049
rect 28261 20040 28273 20043
rect 27396 20012 28273 20040
rect 27396 20000 27402 20012
rect 28261 20009 28273 20012
rect 28307 20009 28319 20043
rect 28261 20003 28319 20009
rect 20088 19972 20116 20000
rect 24029 19975 24087 19981
rect 16040 19944 17632 19972
rect 20088 19944 22692 19972
rect 9401 19907 9459 19913
rect 9401 19873 9413 19907
rect 9447 19904 9459 19907
rect 9766 19904 9772 19916
rect 9447 19876 9772 19904
rect 9447 19873 9459 19876
rect 9401 19867 9459 19873
rect 9766 19864 9772 19876
rect 9824 19864 9830 19916
rect 11885 19907 11943 19913
rect 11885 19873 11897 19907
rect 11931 19904 11943 19907
rect 12342 19904 12348 19916
rect 11931 19876 12348 19904
rect 11931 19873 11943 19876
rect 11885 19867 11943 19873
rect 2038 19836 2044 19848
rect 1999 19808 2044 19836
rect 2038 19796 2044 19808
rect 2096 19796 2102 19848
rect 3973 19839 4031 19845
rect 3973 19836 3985 19839
rect 3436 19808 3985 19836
rect 2308 19771 2366 19777
rect 2308 19737 2320 19771
rect 2354 19768 2366 19771
rect 2774 19768 2780 19780
rect 2354 19740 2780 19768
rect 2354 19737 2366 19740
rect 2308 19731 2366 19737
rect 2774 19728 2780 19740
rect 2832 19728 2838 19780
rect 3436 19709 3464 19808
rect 3973 19805 3985 19808
rect 4019 19805 4031 19839
rect 3973 19799 4031 19805
rect 6638 19796 6644 19848
rect 6696 19836 6702 19848
rect 6733 19839 6791 19845
rect 6733 19836 6745 19839
rect 6696 19808 6745 19836
rect 6696 19796 6702 19808
rect 6733 19805 6745 19808
rect 6779 19805 6791 19839
rect 9306 19836 9312 19848
rect 9267 19808 9312 19836
rect 6733 19799 6791 19805
rect 9306 19796 9312 19808
rect 9364 19796 9370 19848
rect 10594 19796 10600 19848
rect 10652 19836 10658 19848
rect 11900 19836 11928 19867
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 12710 19864 12716 19916
rect 12768 19904 12774 19916
rect 13173 19907 13231 19913
rect 13173 19904 13185 19907
rect 12768 19876 13185 19904
rect 12768 19864 12774 19876
rect 13173 19873 13185 19876
rect 13219 19873 13231 19907
rect 14550 19904 14556 19916
rect 14511 19876 14556 19904
rect 13173 19867 13231 19873
rect 14550 19864 14556 19876
rect 14608 19864 14614 19916
rect 16040 19848 16068 19944
rect 16758 19904 16764 19916
rect 16719 19876 16764 19904
rect 16758 19864 16764 19876
rect 16816 19864 16822 19916
rect 12986 19836 12992 19848
rect 10652 19808 11928 19836
rect 12947 19808 12992 19836
rect 10652 19796 10658 19808
rect 12986 19796 12992 19808
rect 13044 19796 13050 19848
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19836 13599 19839
rect 16022 19836 16028 19848
rect 13587 19808 16028 19836
rect 13587 19805 13599 19808
rect 13541 19799 13599 19805
rect 16022 19796 16028 19808
rect 16080 19796 16086 19848
rect 16577 19839 16635 19845
rect 16577 19805 16589 19839
rect 16623 19805 16635 19839
rect 16942 19836 16948 19848
rect 16903 19808 16948 19836
rect 16577 19799 16635 19805
rect 5902 19728 5908 19780
rect 5960 19768 5966 19780
rect 7009 19771 7067 19777
rect 7009 19768 7021 19771
rect 5960 19740 7021 19768
rect 5960 19728 5966 19740
rect 7009 19737 7021 19740
rect 7055 19737 7067 19771
rect 7009 19731 7067 19737
rect 7466 19728 7472 19780
rect 7524 19728 7530 19780
rect 11606 19768 11612 19780
rect 11664 19777 11670 19780
rect 11576 19740 11612 19768
rect 11606 19728 11612 19740
rect 11664 19731 11676 19777
rect 15381 19771 15439 19777
rect 15381 19737 15393 19771
rect 15427 19768 15439 19771
rect 16482 19768 16488 19780
rect 15427 19740 16488 19768
rect 15427 19737 15439 19740
rect 15381 19731 15439 19737
rect 11664 19728 11670 19731
rect 16482 19728 16488 19740
rect 16540 19728 16546 19780
rect 3421 19703 3479 19709
rect 3421 19669 3433 19703
rect 3467 19669 3479 19703
rect 3421 19663 3479 19669
rect 4338 19660 4344 19712
rect 4396 19700 4402 19712
rect 5169 19703 5227 19709
rect 5169 19700 5181 19703
rect 4396 19672 5181 19700
rect 4396 19660 4402 19672
rect 5169 19669 5181 19672
rect 5215 19669 5227 19703
rect 5169 19663 5227 19669
rect 13354 19660 13360 19712
rect 13412 19700 13418 19712
rect 16592 19700 16620 19799
rect 16942 19796 16948 19808
rect 17000 19796 17006 19848
rect 17604 19845 17632 19944
rect 22664 19916 22692 19944
rect 24029 19941 24041 19975
rect 24075 19941 24087 19975
rect 24029 19935 24087 19941
rect 22646 19904 22652 19916
rect 22559 19876 22652 19904
rect 22646 19864 22652 19876
rect 22704 19864 22710 19916
rect 24044 19904 24072 19935
rect 24762 19904 24768 19916
rect 24044 19876 24768 19904
rect 24762 19864 24768 19876
rect 24820 19904 24826 19916
rect 25041 19907 25099 19913
rect 25041 19904 25053 19907
rect 24820 19876 25053 19904
rect 24820 19864 24826 19876
rect 25041 19873 25053 19876
rect 25087 19873 25099 19907
rect 25041 19867 25099 19873
rect 25130 19864 25136 19916
rect 25188 19904 25194 19916
rect 26786 19904 26792 19916
rect 25188 19876 25233 19904
rect 26747 19876 26792 19904
rect 25188 19864 25194 19876
rect 26786 19864 26792 19876
rect 26844 19864 26850 19916
rect 17589 19839 17647 19845
rect 17589 19805 17601 19839
rect 17635 19805 17647 19839
rect 17589 19799 17647 19805
rect 17773 19839 17831 19845
rect 17773 19805 17785 19839
rect 17819 19805 17831 19839
rect 24946 19836 24952 19848
rect 24907 19808 24952 19836
rect 17773 19799 17831 19805
rect 16960 19768 16988 19796
rect 17788 19768 17816 19799
rect 24946 19796 24952 19808
rect 25004 19796 25010 19848
rect 25869 19839 25927 19845
rect 25869 19805 25881 19839
rect 25915 19805 25927 19839
rect 25869 19799 25927 19805
rect 25961 19839 26019 19845
rect 25961 19805 25973 19839
rect 26007 19836 26019 19839
rect 26513 19839 26571 19845
rect 26513 19836 26525 19839
rect 26007 19808 26525 19836
rect 26007 19805 26019 19808
rect 25961 19799 26019 19805
rect 26513 19805 26525 19808
rect 26559 19805 26571 19839
rect 26513 19799 26571 19805
rect 16960 19740 17816 19768
rect 19610 19728 19616 19780
rect 19668 19768 19674 19780
rect 19797 19771 19855 19777
rect 19797 19768 19809 19771
rect 19668 19740 19809 19768
rect 19668 19728 19674 19740
rect 19797 19737 19809 19740
rect 19843 19737 19855 19771
rect 20898 19768 20904 19780
rect 20859 19740 20904 19768
rect 19797 19731 19855 19737
rect 20898 19728 20904 19740
rect 20956 19728 20962 19780
rect 21085 19771 21143 19777
rect 21085 19737 21097 19771
rect 21131 19768 21143 19771
rect 22278 19768 22284 19780
rect 21131 19740 22284 19768
rect 21131 19737 21143 19740
rect 21085 19731 21143 19737
rect 22278 19728 22284 19740
rect 22336 19728 22342 19780
rect 22916 19771 22974 19777
rect 22916 19737 22928 19771
rect 22962 19768 22974 19771
rect 25884 19768 25912 19799
rect 26326 19768 26332 19780
rect 22962 19740 24624 19768
rect 25884 19740 26332 19768
rect 22962 19737 22974 19740
rect 22916 19731 22974 19737
rect 17034 19700 17040 19712
rect 13412 19672 17040 19700
rect 13412 19660 13418 19672
rect 17034 19660 17040 19672
rect 17092 19660 17098 19712
rect 24596 19709 24624 19740
rect 26326 19728 26332 19740
rect 26384 19728 26390 19780
rect 28074 19768 28080 19780
rect 28014 19740 28080 19768
rect 28074 19728 28080 19740
rect 28132 19728 28138 19780
rect 24581 19703 24639 19709
rect 24581 19669 24593 19703
rect 24627 19669 24639 19703
rect 24581 19663 24639 19669
rect 1104 19610 29048 19632
rect 1104 19558 7896 19610
rect 7948 19558 7960 19610
rect 8012 19558 8024 19610
rect 8076 19558 8088 19610
rect 8140 19558 8152 19610
rect 8204 19558 14842 19610
rect 14894 19558 14906 19610
rect 14958 19558 14970 19610
rect 15022 19558 15034 19610
rect 15086 19558 15098 19610
rect 15150 19558 21788 19610
rect 21840 19558 21852 19610
rect 21904 19558 21916 19610
rect 21968 19558 21980 19610
rect 22032 19558 22044 19610
rect 22096 19558 28734 19610
rect 28786 19558 28798 19610
rect 28850 19558 28862 19610
rect 28914 19558 28926 19610
rect 28978 19558 28990 19610
rect 29042 19558 29048 19610
rect 1104 19536 29048 19558
rect 3142 19456 3148 19508
rect 3200 19496 3206 19508
rect 5902 19496 5908 19508
rect 3200 19468 5212 19496
rect 5863 19468 5908 19496
rect 3200 19456 3206 19468
rect 4338 19428 4344 19440
rect 4299 19400 4344 19428
rect 4338 19388 4344 19400
rect 4396 19388 4402 19440
rect 2961 19363 3019 19369
rect 2961 19329 2973 19363
rect 3007 19360 3019 19363
rect 3007 19332 4844 19360
rect 3007 19329 3019 19332
rect 2961 19323 3019 19329
rect 2774 19252 2780 19304
rect 2832 19292 2838 19304
rect 3142 19292 3148 19304
rect 2832 19264 2877 19292
rect 3103 19264 3148 19292
rect 2832 19252 2838 19264
rect 3142 19252 3148 19264
rect 3200 19252 3206 19304
rect 3234 19252 3240 19304
rect 3292 19292 3298 19304
rect 4816 19292 4844 19332
rect 4890 19320 4896 19372
rect 4948 19360 4954 19372
rect 5184 19369 5212 19468
rect 5902 19456 5908 19468
rect 5960 19456 5966 19508
rect 6638 19496 6644 19508
rect 6599 19468 6644 19496
rect 6638 19456 6644 19468
rect 6696 19456 6702 19508
rect 7742 19456 7748 19508
rect 7800 19496 7806 19508
rect 8573 19499 8631 19505
rect 8573 19496 8585 19499
rect 7800 19468 8585 19496
rect 7800 19456 7806 19468
rect 8573 19465 8585 19468
rect 8619 19465 8631 19499
rect 9490 19496 9496 19508
rect 9451 19468 9496 19496
rect 8573 19459 8631 19465
rect 9490 19456 9496 19468
rect 9548 19456 9554 19508
rect 11606 19456 11612 19508
rect 11664 19496 11670 19508
rect 11701 19499 11759 19505
rect 11701 19496 11713 19499
rect 11664 19468 11713 19496
rect 11664 19456 11670 19468
rect 11701 19465 11713 19468
rect 11747 19465 11759 19499
rect 13262 19496 13268 19508
rect 11701 19459 11759 19465
rect 11808 19468 13268 19496
rect 7098 19428 7104 19440
rect 5276 19400 7104 19428
rect 5077 19363 5135 19369
rect 4948 19332 4993 19360
rect 4948 19320 4954 19332
rect 5077 19329 5089 19363
rect 5123 19329 5135 19363
rect 5077 19323 5135 19329
rect 5169 19363 5227 19369
rect 5169 19329 5181 19363
rect 5215 19329 5227 19363
rect 5169 19323 5227 19329
rect 5092 19292 5120 19323
rect 5276 19292 5304 19400
rect 7098 19388 7104 19400
rect 7156 19388 7162 19440
rect 7460 19431 7518 19437
rect 7460 19397 7472 19431
rect 7506 19428 7518 19431
rect 7558 19428 7564 19440
rect 7506 19400 7564 19428
rect 7506 19397 7518 19400
rect 7460 19391 7518 19397
rect 7558 19388 7564 19400
rect 7616 19388 7622 19440
rect 7650 19388 7656 19440
rect 7708 19428 7714 19440
rect 11808 19428 11836 19468
rect 13262 19456 13268 19468
rect 13320 19456 13326 19508
rect 16209 19499 16267 19505
rect 16209 19465 16221 19499
rect 16255 19496 16267 19499
rect 16298 19496 16304 19508
rect 16255 19468 16304 19496
rect 16255 19465 16267 19468
rect 16209 19459 16267 19465
rect 16298 19456 16304 19468
rect 16356 19456 16362 19508
rect 16850 19496 16856 19508
rect 16811 19468 16856 19496
rect 16850 19456 16856 19468
rect 16908 19456 16914 19508
rect 20898 19456 20904 19508
rect 20956 19496 20962 19508
rect 21085 19499 21143 19505
rect 21085 19496 21097 19499
rect 20956 19468 21097 19496
rect 20956 19456 20962 19468
rect 21085 19465 21097 19468
rect 21131 19465 21143 19499
rect 22186 19496 22192 19508
rect 22147 19468 22192 19496
rect 21085 19459 21143 19465
rect 12158 19428 12164 19440
rect 7708 19400 11836 19428
rect 12119 19400 12164 19428
rect 7708 19388 7714 19400
rect 5994 19360 6000 19372
rect 5955 19332 6000 19360
rect 5994 19320 6000 19332
rect 6052 19320 6058 19372
rect 6549 19363 6607 19369
rect 6549 19329 6561 19363
rect 6595 19360 6607 19363
rect 8294 19360 8300 19372
rect 6595 19332 8300 19360
rect 6595 19329 6607 19332
rect 6549 19323 6607 19329
rect 8294 19320 8300 19332
rect 8352 19360 8358 19372
rect 9306 19360 9312 19372
rect 8352 19332 9312 19360
rect 8352 19320 8358 19332
rect 9306 19320 9312 19332
rect 9364 19320 9370 19372
rect 9585 19363 9643 19369
rect 9585 19329 9597 19363
rect 9631 19360 9643 19363
rect 9766 19360 9772 19372
rect 9631 19332 9772 19360
rect 9631 19329 9643 19332
rect 9585 19323 9643 19329
rect 9766 19320 9772 19332
rect 9824 19320 9830 19372
rect 10336 19369 10364 19400
rect 12158 19388 12164 19400
rect 12216 19388 12222 19440
rect 16574 19388 16580 19440
rect 16632 19428 16638 19440
rect 17770 19428 17776 19440
rect 16632 19400 17776 19428
rect 16632 19388 16638 19400
rect 17770 19388 17776 19400
rect 17828 19428 17834 19440
rect 17954 19428 17960 19440
rect 17828 19400 17960 19428
rect 17828 19388 17834 19400
rect 17954 19388 17960 19400
rect 18012 19388 18018 19440
rect 20070 19428 20076 19440
rect 19720 19400 20076 19428
rect 10321 19363 10379 19369
rect 10321 19329 10333 19363
rect 10367 19329 10379 19363
rect 12066 19360 12072 19372
rect 12027 19332 12072 19360
rect 10321 19323 10379 19329
rect 12066 19320 12072 19332
rect 12124 19320 12130 19372
rect 12986 19320 12992 19372
rect 13044 19360 13050 19372
rect 13081 19363 13139 19369
rect 13081 19360 13093 19363
rect 13044 19332 13093 19360
rect 13044 19320 13050 19332
rect 13081 19329 13093 19332
rect 13127 19329 13139 19363
rect 13262 19360 13268 19372
rect 13223 19332 13268 19360
rect 13081 19323 13139 19329
rect 3292 19264 3337 19292
rect 4816 19264 4936 19292
rect 5092 19264 5304 19292
rect 3292 19252 3298 19264
rect 4908 19233 4936 19264
rect 7098 19252 7104 19304
rect 7156 19292 7162 19304
rect 7193 19295 7251 19301
rect 7193 19292 7205 19295
rect 7156 19264 7205 19292
rect 7156 19252 7162 19264
rect 7193 19261 7205 19264
rect 7239 19261 7251 19295
rect 7193 19255 7251 19261
rect 9490 19252 9496 19304
rect 9548 19292 9554 19304
rect 9677 19295 9735 19301
rect 9677 19292 9689 19295
rect 9548 19264 9689 19292
rect 9548 19252 9554 19264
rect 9677 19261 9689 19264
rect 9723 19292 9735 19295
rect 12253 19295 12311 19301
rect 12253 19292 12265 19295
rect 9723 19264 12265 19292
rect 9723 19261 9735 19264
rect 9677 19255 9735 19261
rect 12253 19261 12265 19264
rect 12299 19292 12311 19295
rect 12897 19295 12955 19301
rect 12897 19292 12909 19295
rect 12299 19264 12909 19292
rect 12299 19261 12311 19264
rect 12253 19255 12311 19261
rect 12897 19261 12909 19264
rect 12943 19261 12955 19295
rect 13096 19292 13124 19323
rect 13262 19320 13268 19332
rect 13320 19320 13326 19372
rect 13909 19363 13967 19369
rect 13909 19360 13921 19363
rect 13556 19332 13921 19360
rect 13556 19304 13584 19332
rect 13909 19329 13921 19332
rect 13955 19329 13967 19363
rect 14182 19360 14188 19372
rect 14143 19332 14188 19360
rect 13909 19323 13967 19329
rect 14182 19320 14188 19332
rect 14240 19320 14246 19372
rect 16022 19360 16028 19372
rect 15983 19332 16028 19360
rect 16022 19320 16028 19332
rect 16080 19320 16086 19372
rect 17034 19360 17040 19372
rect 16995 19332 17040 19360
rect 17034 19320 17040 19332
rect 17092 19320 17098 19372
rect 19720 19369 19748 19400
rect 20070 19388 20076 19400
rect 20128 19388 20134 19440
rect 21100 19428 21128 19459
rect 22186 19456 22192 19468
rect 22244 19456 22250 19508
rect 28074 19456 28080 19508
rect 28132 19496 28138 19508
rect 28261 19499 28319 19505
rect 28261 19496 28273 19499
rect 28132 19468 28273 19496
rect 28132 19456 28138 19468
rect 28261 19465 28273 19468
rect 28307 19465 28319 19499
rect 28261 19459 28319 19465
rect 21726 19428 21732 19440
rect 21100 19400 21732 19428
rect 21726 19388 21732 19400
rect 21784 19428 21790 19440
rect 21784 19400 22048 19428
rect 21784 19388 21790 19400
rect 19705 19363 19763 19369
rect 19705 19329 19717 19363
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 19972 19363 20030 19369
rect 19972 19329 19984 19363
rect 20018 19360 20030 19363
rect 21266 19360 21272 19372
rect 20018 19332 21272 19360
rect 20018 19329 20030 19332
rect 19972 19323 20030 19329
rect 21266 19320 21272 19332
rect 21324 19320 21330 19372
rect 22020 19369 22048 19400
rect 22005 19363 22063 19369
rect 22005 19329 22017 19363
rect 22051 19329 22063 19363
rect 22186 19360 22192 19372
rect 22147 19332 22192 19360
rect 22005 19323 22063 19329
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 22646 19360 22652 19372
rect 22607 19332 22652 19360
rect 22646 19320 22652 19332
rect 22704 19320 22710 19372
rect 22922 19369 22928 19372
rect 22916 19323 22928 19369
rect 22980 19360 22986 19372
rect 24949 19363 25007 19369
rect 22980 19332 23016 19360
rect 22922 19320 22928 19323
rect 22980 19320 22986 19332
rect 24949 19329 24961 19363
rect 24995 19360 25007 19363
rect 26145 19363 26203 19369
rect 26145 19360 26157 19363
rect 24995 19332 26157 19360
rect 24995 19329 25007 19332
rect 24949 19323 25007 19329
rect 26145 19329 26157 19332
rect 26191 19360 26203 19363
rect 26326 19360 26332 19372
rect 26191 19332 26332 19360
rect 26191 19329 26203 19332
rect 26145 19323 26203 19329
rect 26326 19320 26332 19332
rect 26384 19320 26390 19372
rect 27430 19360 27436 19372
rect 27391 19332 27436 19360
rect 27430 19320 27436 19332
rect 27488 19320 27494 19372
rect 13538 19292 13544 19304
rect 13096 19264 13544 19292
rect 12897 19255 12955 19261
rect 13538 19252 13544 19264
rect 13596 19252 13602 19304
rect 14277 19295 14335 19301
rect 14277 19261 14289 19295
rect 14323 19292 14335 19295
rect 14642 19292 14648 19304
rect 14323 19264 14648 19292
rect 14323 19261 14335 19264
rect 14277 19255 14335 19261
rect 14642 19252 14648 19264
rect 14700 19252 14706 19304
rect 15194 19252 15200 19304
rect 15252 19292 15258 19304
rect 15841 19295 15899 19301
rect 15841 19292 15853 19295
rect 15252 19264 15853 19292
rect 15252 19252 15258 19264
rect 15841 19261 15853 19264
rect 15887 19292 15899 19295
rect 17221 19295 17279 19301
rect 17221 19292 17233 19295
rect 15887 19264 17233 19292
rect 15887 19261 15899 19264
rect 15841 19255 15899 19261
rect 17221 19261 17233 19264
rect 17267 19261 17279 19295
rect 17221 19255 17279 19261
rect 17494 19252 17500 19304
rect 17552 19292 17558 19304
rect 19610 19292 19616 19304
rect 17552 19264 19616 19292
rect 17552 19252 17558 19264
rect 19610 19252 19616 19264
rect 19668 19252 19674 19304
rect 23842 19252 23848 19304
rect 23900 19292 23906 19304
rect 24581 19295 24639 19301
rect 24581 19292 24593 19295
rect 23900 19264 24593 19292
rect 23900 19252 23906 19264
rect 24581 19261 24593 19264
rect 24627 19261 24639 19295
rect 24581 19255 24639 19261
rect 24857 19295 24915 19301
rect 24857 19261 24869 19295
rect 24903 19261 24915 19295
rect 24857 19255 24915 19261
rect 4893 19227 4951 19233
rect 4893 19193 4905 19227
rect 4939 19193 4951 19227
rect 4893 19187 4951 19193
rect 10505 19227 10563 19233
rect 10505 19193 10517 19227
rect 10551 19224 10563 19227
rect 10594 19224 10600 19236
rect 10551 19196 10600 19224
rect 10551 19193 10563 19196
rect 10505 19187 10563 19193
rect 10594 19184 10600 19196
rect 10652 19184 10658 19236
rect 13630 19184 13636 19236
rect 13688 19224 13694 19236
rect 17512 19224 17540 19252
rect 22554 19224 22560 19236
rect 13688 19196 17540 19224
rect 22066 19196 22560 19224
rect 13688 19184 13694 19196
rect 4065 19159 4123 19165
rect 4065 19125 4077 19159
rect 4111 19156 4123 19159
rect 4246 19156 4252 19168
rect 4111 19128 4252 19156
rect 4111 19125 4123 19128
rect 4065 19119 4123 19125
rect 4246 19116 4252 19128
rect 4304 19156 4310 19168
rect 5074 19156 5080 19168
rect 4304 19128 5080 19156
rect 4304 19116 4310 19128
rect 5074 19116 5080 19128
rect 5132 19156 5138 19168
rect 7558 19156 7564 19168
rect 5132 19128 7564 19156
rect 5132 19116 5138 19128
rect 7558 19116 7564 19128
rect 7616 19116 7622 19168
rect 9125 19159 9183 19165
rect 9125 19125 9137 19159
rect 9171 19156 9183 19159
rect 9214 19156 9220 19168
rect 9171 19128 9220 19156
rect 9171 19125 9183 19128
rect 9125 19119 9183 19125
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 18230 19116 18236 19168
rect 18288 19156 18294 19168
rect 19886 19156 19892 19168
rect 18288 19128 19892 19156
rect 18288 19116 18294 19128
rect 19886 19116 19892 19128
rect 19944 19116 19950 19168
rect 21174 19116 21180 19168
rect 21232 19156 21238 19168
rect 22066 19156 22094 19196
rect 22554 19184 22560 19196
rect 22612 19184 22618 19236
rect 24026 19224 24032 19236
rect 23939 19196 24032 19224
rect 24026 19184 24032 19196
rect 24084 19224 24090 19236
rect 24872 19224 24900 19255
rect 26234 19252 26240 19304
rect 26292 19292 26298 19304
rect 27341 19295 27399 19301
rect 27341 19292 27353 19295
rect 26292 19264 27353 19292
rect 26292 19252 26298 19264
rect 27341 19261 27353 19264
rect 27387 19261 27399 19295
rect 27341 19255 27399 19261
rect 24084 19196 24900 19224
rect 24084 19184 24090 19196
rect 21232 19128 22094 19156
rect 21232 19116 21238 19128
rect 25958 19116 25964 19168
rect 26016 19156 26022 19168
rect 26053 19159 26111 19165
rect 26053 19156 26065 19159
rect 26016 19128 26065 19156
rect 26016 19116 26022 19128
rect 26053 19125 26065 19128
rect 26099 19125 26111 19159
rect 26053 19119 26111 19125
rect 1104 19066 28888 19088
rect 1104 19014 4423 19066
rect 4475 19014 4487 19066
rect 4539 19014 4551 19066
rect 4603 19014 4615 19066
rect 4667 19014 4679 19066
rect 4731 19014 11369 19066
rect 11421 19014 11433 19066
rect 11485 19014 11497 19066
rect 11549 19014 11561 19066
rect 11613 19014 11625 19066
rect 11677 19014 18315 19066
rect 18367 19014 18379 19066
rect 18431 19014 18443 19066
rect 18495 19014 18507 19066
rect 18559 19014 18571 19066
rect 18623 19014 25261 19066
rect 25313 19014 25325 19066
rect 25377 19014 25389 19066
rect 25441 19014 25453 19066
rect 25505 19014 25517 19066
rect 25569 19014 28888 19066
rect 1104 18992 28888 19014
rect 9766 18912 9772 18964
rect 9824 18952 9830 18964
rect 10505 18955 10563 18961
rect 10505 18952 10517 18955
rect 9824 18924 10517 18952
rect 9824 18912 9830 18924
rect 10505 18921 10517 18924
rect 10551 18921 10563 18955
rect 10505 18915 10563 18921
rect 12526 18912 12532 18964
rect 12584 18952 12590 18964
rect 12989 18955 13047 18961
rect 12989 18952 13001 18955
rect 12584 18924 13001 18952
rect 12584 18912 12590 18924
rect 12989 18921 13001 18924
rect 13035 18921 13047 18955
rect 21266 18952 21272 18964
rect 21227 18924 21272 18952
rect 12989 18915 13047 18921
rect 21266 18912 21272 18924
rect 21324 18912 21330 18964
rect 22922 18952 22928 18964
rect 22883 18924 22928 18952
rect 22922 18912 22928 18924
rect 22980 18912 22986 18964
rect 26326 18912 26332 18964
rect 26384 18952 26390 18964
rect 27433 18955 27491 18961
rect 27433 18952 27445 18955
rect 26384 18924 27445 18952
rect 26384 18912 26390 18924
rect 27433 18921 27445 18924
rect 27479 18921 27491 18955
rect 27433 18915 27491 18921
rect 5534 18844 5540 18896
rect 5592 18884 5598 18896
rect 16025 18887 16083 18893
rect 5592 18856 5948 18884
rect 5592 18844 5598 18856
rect 5920 18828 5948 18856
rect 16025 18853 16037 18887
rect 16071 18884 16083 18887
rect 17221 18887 17279 18893
rect 16071 18856 17172 18884
rect 16071 18853 16083 18856
rect 16025 18847 16083 18853
rect 2038 18776 2044 18828
rect 2096 18816 2102 18828
rect 2096 18788 4200 18816
rect 2096 18776 2102 18788
rect 2866 18708 2872 18760
rect 2924 18748 2930 18760
rect 4172 18757 4200 18788
rect 5902 18776 5908 18828
rect 5960 18816 5966 18828
rect 6733 18819 6791 18825
rect 5960 18788 6005 18816
rect 5960 18776 5966 18788
rect 6733 18785 6745 18819
rect 6779 18816 6791 18819
rect 7466 18816 7472 18828
rect 6779 18788 7472 18816
rect 6779 18785 6791 18788
rect 6733 18779 6791 18785
rect 7466 18776 7472 18788
rect 7524 18776 7530 18828
rect 13446 18825 13452 18828
rect 13432 18819 13452 18825
rect 13432 18816 13444 18819
rect 13359 18788 13444 18816
rect 13432 18785 13444 18788
rect 13504 18816 13510 18828
rect 17144 18816 17172 18856
rect 17221 18853 17233 18887
rect 17267 18884 17279 18887
rect 21174 18884 21180 18896
rect 17267 18856 21180 18884
rect 17267 18853 17279 18856
rect 17221 18847 17279 18853
rect 21174 18844 21180 18856
rect 21232 18844 21238 18896
rect 21560 18856 22094 18884
rect 21560 18816 21588 18856
rect 21726 18816 21732 18828
rect 13504 18788 16988 18816
rect 17144 18788 21588 18816
rect 21687 18788 21732 18816
rect 13432 18779 13452 18785
rect 13446 18776 13452 18779
rect 13504 18776 13510 18788
rect 5816 18760 5868 18766
rect 3973 18751 4031 18757
rect 3973 18748 3985 18751
rect 2924 18720 3985 18748
rect 2924 18708 2930 18720
rect 3973 18717 3985 18720
rect 4019 18717 4031 18751
rect 3973 18711 4031 18717
rect 4157 18751 4215 18757
rect 4157 18717 4169 18751
rect 4203 18717 4215 18751
rect 4157 18711 4215 18717
rect 9125 18751 9183 18757
rect 9125 18717 9137 18751
rect 9171 18717 9183 18751
rect 9125 18711 9183 18717
rect 5816 18702 5868 18708
rect 4338 18680 4344 18692
rect 4299 18652 4344 18680
rect 4338 18640 4344 18652
rect 4396 18640 4402 18692
rect 9140 18680 9168 18711
rect 9214 18708 9220 18760
rect 9272 18748 9278 18760
rect 9381 18751 9439 18757
rect 9381 18748 9393 18751
rect 9272 18720 9393 18748
rect 9272 18708 9278 18720
rect 9381 18717 9393 18720
rect 9427 18717 9439 18751
rect 9381 18711 9439 18717
rect 13538 18708 13544 18760
rect 13596 18748 13602 18760
rect 13633 18751 13691 18757
rect 13633 18748 13645 18751
rect 13596 18720 13645 18748
rect 13596 18708 13602 18720
rect 13633 18717 13645 18720
rect 13679 18717 13691 18751
rect 13633 18711 13691 18717
rect 13725 18751 13783 18757
rect 13725 18717 13737 18751
rect 13771 18748 13783 18751
rect 14734 18748 14740 18760
rect 13771 18720 14740 18748
rect 13771 18717 13783 18720
rect 13725 18711 13783 18717
rect 14734 18708 14740 18720
rect 14792 18708 14798 18760
rect 15286 18708 15292 18760
rect 15344 18748 15350 18760
rect 16960 18757 16988 18788
rect 21726 18776 21732 18788
rect 21784 18776 21790 18828
rect 21836 18825 21864 18856
rect 21821 18819 21879 18825
rect 21821 18785 21833 18819
rect 21867 18785 21879 18819
rect 22066 18816 22094 18856
rect 22186 18844 22192 18896
rect 22244 18884 22250 18896
rect 22244 18856 24992 18884
rect 22244 18844 22250 18856
rect 23477 18819 23535 18825
rect 23477 18816 23489 18819
rect 22066 18788 23489 18816
rect 21821 18779 21879 18785
rect 23477 18785 23489 18788
rect 23523 18816 23535 18819
rect 23523 18788 24900 18816
rect 23523 18785 23535 18788
rect 23477 18779 23535 18785
rect 15933 18751 15991 18757
rect 15933 18748 15945 18751
rect 15344 18720 15945 18748
rect 15344 18708 15350 18720
rect 15933 18717 15945 18720
rect 15979 18717 15991 18751
rect 15933 18711 15991 18717
rect 16117 18751 16175 18757
rect 16117 18717 16129 18751
rect 16163 18717 16175 18751
rect 16117 18711 16175 18717
rect 16761 18751 16819 18757
rect 16761 18717 16773 18751
rect 16807 18717 16819 18751
rect 16761 18711 16819 18717
rect 16945 18751 17003 18757
rect 16945 18717 16957 18751
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 17313 18751 17371 18757
rect 17313 18717 17325 18751
rect 17359 18748 17371 18751
rect 17402 18748 17408 18760
rect 17359 18720 17408 18748
rect 17359 18717 17371 18720
rect 17313 18711 17371 18717
rect 10594 18680 10600 18692
rect 9140 18652 10600 18680
rect 10594 18640 10600 18652
rect 10652 18640 10658 18692
rect 13170 18680 13176 18692
rect 13131 18652 13176 18680
rect 13170 18640 13176 18652
rect 13228 18640 13234 18692
rect 14274 18640 14280 18692
rect 14332 18680 14338 18692
rect 16132 18680 16160 18711
rect 14332 18652 16160 18680
rect 14332 18640 14338 18652
rect 13541 18615 13599 18621
rect 13541 18581 13553 18615
rect 13587 18612 13599 18615
rect 13630 18612 13636 18624
rect 13587 18584 13636 18612
rect 13587 18581 13599 18584
rect 13541 18575 13599 18581
rect 13630 18572 13636 18584
rect 13688 18572 13694 18624
rect 16776 18612 16804 18711
rect 17402 18708 17408 18720
rect 17460 18708 17466 18760
rect 18230 18748 18236 18760
rect 18191 18720 18236 18748
rect 18230 18708 18236 18720
rect 18288 18708 18294 18760
rect 18509 18751 18567 18757
rect 18509 18717 18521 18751
rect 18555 18748 18567 18751
rect 19794 18748 19800 18760
rect 18555 18720 19800 18748
rect 18555 18717 18567 18720
rect 18509 18711 18567 18717
rect 19794 18708 19800 18720
rect 19852 18708 19858 18760
rect 19886 18708 19892 18760
rect 19944 18748 19950 18760
rect 20806 18748 20812 18760
rect 19944 18720 19989 18748
rect 20767 18720 20812 18748
rect 19944 18708 19950 18720
rect 20806 18708 20812 18720
rect 20864 18708 20870 18760
rect 23385 18751 23443 18757
rect 23385 18717 23397 18751
rect 23431 18748 23443 18751
rect 24026 18748 24032 18760
rect 23431 18720 24032 18748
rect 23431 18717 23443 18720
rect 23385 18711 23443 18717
rect 24026 18708 24032 18720
rect 24084 18708 24090 18760
rect 24872 18680 24900 18788
rect 24964 18757 24992 18856
rect 25958 18816 25964 18828
rect 25919 18788 25964 18816
rect 25958 18776 25964 18788
rect 26016 18776 26022 18828
rect 24949 18751 25007 18757
rect 24949 18717 24961 18751
rect 24995 18717 25007 18751
rect 24949 18711 25007 18717
rect 25041 18751 25099 18757
rect 25041 18717 25053 18751
rect 25087 18748 25099 18751
rect 25685 18751 25743 18757
rect 25685 18748 25697 18751
rect 25087 18720 25697 18748
rect 25087 18717 25099 18720
rect 25041 18711 25099 18717
rect 25685 18717 25697 18720
rect 25731 18717 25743 18751
rect 25685 18711 25743 18717
rect 25130 18680 25136 18692
rect 18708 18652 19656 18680
rect 24872 18652 25136 18680
rect 18708 18612 18736 18652
rect 18874 18612 18880 18624
rect 16776 18584 18736 18612
rect 18835 18584 18880 18612
rect 18874 18572 18880 18584
rect 18932 18572 18938 18624
rect 19628 18612 19656 18652
rect 25130 18640 25136 18652
rect 25188 18640 25194 18692
rect 26602 18640 26608 18692
rect 26660 18640 26666 18692
rect 20254 18612 20260 18624
rect 19628 18584 20260 18612
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 21634 18612 21640 18624
rect 21595 18584 21640 18612
rect 21634 18572 21640 18584
rect 21692 18572 21698 18624
rect 23014 18572 23020 18624
rect 23072 18612 23078 18624
rect 23293 18615 23351 18621
rect 23293 18612 23305 18615
rect 23072 18584 23305 18612
rect 23072 18572 23078 18584
rect 23293 18581 23305 18584
rect 23339 18581 23351 18615
rect 23293 18575 23351 18581
rect 1104 18522 29048 18544
rect 1104 18470 7896 18522
rect 7948 18470 7960 18522
rect 8012 18470 8024 18522
rect 8076 18470 8088 18522
rect 8140 18470 8152 18522
rect 8204 18470 14842 18522
rect 14894 18470 14906 18522
rect 14958 18470 14970 18522
rect 15022 18470 15034 18522
rect 15086 18470 15098 18522
rect 15150 18470 21788 18522
rect 21840 18470 21852 18522
rect 21904 18470 21916 18522
rect 21968 18470 21980 18522
rect 22032 18470 22044 18522
rect 22096 18470 28734 18522
rect 28786 18470 28798 18522
rect 28850 18470 28862 18522
rect 28914 18470 28926 18522
rect 28978 18470 28990 18522
rect 29042 18470 29048 18522
rect 1104 18448 29048 18470
rect 4893 18411 4951 18417
rect 4893 18408 4905 18411
rect 2884 18380 4905 18408
rect 2884 18352 2912 18380
rect 4893 18377 4905 18380
rect 4939 18377 4951 18411
rect 4893 18371 4951 18377
rect 14734 18368 14740 18420
rect 14792 18408 14798 18420
rect 14829 18411 14887 18417
rect 14829 18408 14841 18411
rect 14792 18380 14841 18408
rect 14792 18368 14798 18380
rect 14829 18377 14841 18380
rect 14875 18377 14887 18411
rect 17402 18408 17408 18420
rect 17363 18380 17408 18408
rect 14829 18371 14887 18377
rect 17402 18368 17408 18380
rect 17460 18368 17466 18420
rect 19978 18368 19984 18420
rect 20036 18408 20042 18420
rect 20441 18411 20499 18417
rect 20441 18408 20453 18411
rect 20036 18380 20453 18408
rect 20036 18368 20042 18380
rect 20441 18377 20453 18380
rect 20487 18408 20499 18411
rect 22186 18408 22192 18420
rect 20487 18380 22192 18408
rect 20487 18377 20499 18380
rect 20441 18371 20499 18377
rect 22186 18368 22192 18380
rect 22244 18368 22250 18420
rect 26602 18408 26608 18420
rect 26563 18380 26608 18408
rect 26602 18368 26608 18380
rect 26660 18368 26666 18420
rect 2866 18340 2872 18352
rect 2827 18312 2872 18340
rect 2866 18300 2872 18312
rect 2924 18300 2930 18352
rect 5810 18300 5816 18352
rect 5868 18340 5874 18352
rect 7837 18343 7895 18349
rect 7837 18340 7849 18343
rect 5868 18312 7849 18340
rect 5868 18300 5874 18312
rect 7837 18309 7849 18312
rect 7883 18309 7895 18343
rect 9582 18340 9588 18352
rect 9543 18312 9588 18340
rect 7837 18303 7895 18309
rect 9582 18300 9588 18312
rect 9640 18300 9646 18352
rect 17221 18343 17279 18349
rect 17221 18309 17233 18343
rect 17267 18340 17279 18343
rect 17494 18340 17500 18352
rect 17267 18312 17500 18340
rect 17267 18309 17279 18312
rect 17221 18303 17279 18309
rect 17494 18300 17500 18312
rect 17552 18300 17558 18352
rect 18874 18300 18880 18352
rect 18932 18340 18938 18352
rect 18932 18312 19458 18340
rect 18932 18300 18938 18312
rect 20254 18300 20260 18352
rect 20312 18340 20318 18352
rect 24670 18340 24676 18352
rect 20312 18312 24676 18340
rect 20312 18300 20318 18312
rect 24670 18300 24676 18312
rect 24728 18300 24734 18352
rect 3970 18232 3976 18284
rect 4028 18232 4034 18284
rect 4801 18275 4859 18281
rect 4801 18272 4813 18275
rect 4356 18244 4813 18272
rect 4356 18213 4384 18244
rect 4801 18241 4813 18244
rect 4847 18241 4859 18275
rect 6730 18272 6736 18284
rect 6691 18244 6736 18272
rect 4801 18235 4859 18241
rect 6730 18232 6736 18244
rect 6788 18232 6794 18284
rect 12802 18232 12808 18284
rect 12860 18272 12866 18284
rect 13078 18272 13084 18284
rect 12860 18244 13084 18272
rect 12860 18232 12866 18244
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 13541 18275 13599 18281
rect 13541 18241 13553 18275
rect 13587 18272 13599 18275
rect 13722 18272 13728 18284
rect 13587 18244 13728 18272
rect 13587 18241 13599 18244
rect 13541 18235 13599 18241
rect 13722 18232 13728 18244
rect 13780 18232 13786 18284
rect 13909 18275 13967 18281
rect 13909 18241 13921 18275
rect 13955 18272 13967 18275
rect 14642 18272 14648 18284
rect 13955 18244 14648 18272
rect 13955 18241 13967 18244
rect 13909 18235 13967 18241
rect 14642 18232 14648 18244
rect 14700 18232 14706 18284
rect 14921 18275 14979 18281
rect 14921 18241 14933 18275
rect 14967 18241 14979 18275
rect 14921 18235 14979 18241
rect 24949 18275 25007 18281
rect 24949 18241 24961 18275
rect 24995 18272 25007 18275
rect 25130 18272 25136 18284
rect 24995 18244 25136 18272
rect 24995 18241 25007 18244
rect 24949 18235 25007 18241
rect 2593 18207 2651 18213
rect 2593 18173 2605 18207
rect 2639 18173 2651 18207
rect 2593 18167 2651 18173
rect 4341 18207 4399 18213
rect 4341 18173 4353 18207
rect 4387 18173 4399 18207
rect 4341 18167 4399 18173
rect 2608 18068 2636 18167
rect 13814 18164 13820 18216
rect 13872 18204 13878 18216
rect 14093 18207 14151 18213
rect 14093 18204 14105 18207
rect 13872 18176 14105 18204
rect 13872 18164 13878 18176
rect 14093 18173 14105 18176
rect 14139 18173 14151 18207
rect 14093 18167 14151 18173
rect 14274 18164 14280 18216
rect 14332 18204 14338 18216
rect 14936 18204 14964 18235
rect 25130 18232 25136 18244
rect 25188 18232 25194 18284
rect 25774 18272 25780 18284
rect 25735 18244 25780 18272
rect 25774 18232 25780 18244
rect 25832 18232 25838 18284
rect 26234 18272 26240 18284
rect 26195 18244 26240 18272
rect 26234 18232 26240 18244
rect 26292 18232 26298 18284
rect 18690 18204 18696 18216
rect 14332 18176 14964 18204
rect 18651 18176 18696 18204
rect 14332 18164 14338 18176
rect 18690 18164 18696 18176
rect 18748 18164 18754 18216
rect 18969 18207 19027 18213
rect 18969 18173 18981 18207
rect 19015 18204 19027 18207
rect 19702 18204 19708 18216
rect 19015 18176 19708 18204
rect 19015 18173 19027 18176
rect 18969 18167 19027 18173
rect 19702 18164 19708 18176
rect 19760 18164 19766 18216
rect 13538 18136 13544 18148
rect 13499 18108 13544 18136
rect 13538 18096 13544 18108
rect 13596 18096 13602 18148
rect 16574 18096 16580 18148
rect 16632 18136 16638 18148
rect 16853 18139 16911 18145
rect 16853 18136 16865 18139
rect 16632 18108 16865 18136
rect 16632 18096 16638 18108
rect 16853 18105 16865 18108
rect 16899 18105 16911 18139
rect 16853 18099 16911 18105
rect 2866 18068 2872 18080
rect 2608 18040 2872 18068
rect 2866 18028 2872 18040
rect 2924 18028 2930 18080
rect 6546 18028 6552 18080
rect 6604 18068 6610 18080
rect 6641 18071 6699 18077
rect 6641 18068 6653 18071
rect 6604 18040 6653 18068
rect 6604 18028 6610 18040
rect 6641 18037 6653 18040
rect 6687 18037 6699 18071
rect 6641 18031 6699 18037
rect 13078 18028 13084 18080
rect 13136 18068 13142 18080
rect 14366 18068 14372 18080
rect 13136 18040 14372 18068
rect 13136 18028 13142 18040
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 15286 18028 15292 18080
rect 15344 18068 15350 18080
rect 16942 18068 16948 18080
rect 15344 18040 16948 18068
rect 15344 18028 15350 18040
rect 16942 18028 16948 18040
rect 17000 18068 17006 18080
rect 17221 18071 17279 18077
rect 17221 18068 17233 18071
rect 17000 18040 17233 18068
rect 17000 18028 17006 18040
rect 17221 18037 17233 18040
rect 17267 18037 17279 18071
rect 24854 18068 24860 18080
rect 24815 18040 24860 18068
rect 17221 18031 17279 18037
rect 24854 18028 24860 18040
rect 24912 18028 24918 18080
rect 1104 17978 28888 18000
rect 1104 17926 4423 17978
rect 4475 17926 4487 17978
rect 4539 17926 4551 17978
rect 4603 17926 4615 17978
rect 4667 17926 4679 17978
rect 4731 17926 11369 17978
rect 11421 17926 11433 17978
rect 11485 17926 11497 17978
rect 11549 17926 11561 17978
rect 11613 17926 11625 17978
rect 11677 17926 18315 17978
rect 18367 17926 18379 17978
rect 18431 17926 18443 17978
rect 18495 17926 18507 17978
rect 18559 17926 18571 17978
rect 18623 17926 25261 17978
rect 25313 17926 25325 17978
rect 25377 17926 25389 17978
rect 25441 17926 25453 17978
rect 25505 17926 25517 17978
rect 25569 17926 28888 17978
rect 1104 17904 28888 17926
rect 2866 17864 2872 17876
rect 2827 17836 2872 17864
rect 2866 17824 2872 17836
rect 2924 17824 2930 17876
rect 3970 17824 3976 17876
rect 4028 17864 4034 17876
rect 4065 17867 4123 17873
rect 4065 17864 4077 17867
rect 4028 17836 4077 17864
rect 4028 17824 4034 17836
rect 4065 17833 4077 17836
rect 4111 17833 4123 17867
rect 4065 17827 4123 17833
rect 9677 17867 9735 17873
rect 9677 17833 9689 17867
rect 9723 17864 9735 17867
rect 11238 17864 11244 17876
rect 9723 17836 11244 17864
rect 9723 17833 9735 17836
rect 9677 17827 9735 17833
rect 11238 17824 11244 17836
rect 11296 17824 11302 17876
rect 19702 17824 19708 17876
rect 19760 17864 19766 17876
rect 19889 17867 19947 17873
rect 19889 17864 19901 17867
rect 19760 17836 19901 17864
rect 19760 17824 19766 17836
rect 19889 17833 19901 17836
rect 19935 17833 19947 17867
rect 19889 17827 19947 17833
rect 8294 17728 8300 17740
rect 5552 17700 8300 17728
rect 2958 17660 2964 17672
rect 2919 17632 2964 17660
rect 2958 17620 2964 17632
rect 3016 17620 3022 17672
rect 3234 17620 3240 17672
rect 3292 17660 3298 17672
rect 5552 17669 5580 17700
rect 8294 17688 8300 17700
rect 8352 17688 8358 17740
rect 9398 17728 9404 17740
rect 9359 17700 9404 17728
rect 9398 17688 9404 17700
rect 9456 17688 9462 17740
rect 10594 17688 10600 17740
rect 10652 17728 10658 17740
rect 11793 17731 11851 17737
rect 11793 17728 11805 17731
rect 10652 17700 11805 17728
rect 10652 17688 10658 17700
rect 11793 17697 11805 17700
rect 11839 17697 11851 17731
rect 11793 17691 11851 17697
rect 13170 17688 13176 17740
rect 13228 17728 13234 17740
rect 15565 17731 15623 17737
rect 15565 17728 15577 17731
rect 13228 17700 15577 17728
rect 13228 17688 13234 17700
rect 15565 17697 15577 17700
rect 15611 17697 15623 17731
rect 15565 17691 15623 17697
rect 22741 17731 22799 17737
rect 22741 17697 22753 17731
rect 22787 17728 22799 17731
rect 23106 17728 23112 17740
rect 22787 17700 23112 17728
rect 22787 17697 22799 17700
rect 22741 17691 22799 17697
rect 23106 17688 23112 17700
rect 23164 17688 23170 17740
rect 4157 17663 4215 17669
rect 4157 17660 4169 17663
rect 3292 17632 4169 17660
rect 3292 17620 3298 17632
rect 4157 17629 4169 17632
rect 4203 17629 4215 17663
rect 4157 17623 4215 17629
rect 5537 17663 5595 17669
rect 5537 17629 5549 17663
rect 5583 17629 5595 17663
rect 5537 17623 5595 17629
rect 6181 17663 6239 17669
rect 6181 17629 6193 17663
rect 6227 17629 6239 17663
rect 6181 17623 6239 17629
rect 6196 17592 6224 17623
rect 6730 17620 6736 17672
rect 6788 17660 6794 17672
rect 7282 17660 7288 17672
rect 6788 17632 7288 17660
rect 6788 17620 6794 17632
rect 7282 17620 7288 17632
rect 7340 17660 7346 17672
rect 9309 17663 9367 17669
rect 9309 17660 9321 17663
rect 7340 17632 9321 17660
rect 7340 17620 7346 17632
rect 9309 17629 9321 17632
rect 9355 17629 9367 17663
rect 9309 17623 9367 17629
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14553 17663 14611 17669
rect 14553 17660 14565 17663
rect 13872 17632 14565 17660
rect 13872 17620 13878 17632
rect 14553 17629 14565 17632
rect 14599 17629 14611 17663
rect 19978 17660 19984 17672
rect 19939 17632 19984 17660
rect 14553 17623 14611 17629
rect 19978 17620 19984 17632
rect 20036 17620 20042 17672
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17660 24639 17663
rect 24670 17660 24676 17672
rect 24627 17632 24676 17660
rect 24627 17629 24639 17632
rect 24581 17623 24639 17629
rect 24670 17620 24676 17632
rect 24728 17620 24734 17672
rect 24854 17669 24860 17672
rect 24848 17623 24860 17669
rect 24912 17660 24918 17672
rect 24912 17632 24948 17660
rect 24854 17620 24860 17623
rect 24912 17620 24918 17632
rect 27614 17620 27620 17672
rect 27672 17660 27678 17672
rect 27893 17663 27951 17669
rect 27893 17660 27905 17663
rect 27672 17632 27905 17660
rect 27672 17620 27678 17632
rect 27893 17629 27905 17632
rect 27939 17629 27951 17663
rect 27893 17623 27951 17629
rect 6362 17592 6368 17604
rect 6196 17564 6368 17592
rect 6362 17552 6368 17564
rect 6420 17592 6426 17604
rect 7193 17595 7251 17601
rect 6420 17564 6960 17592
rect 6420 17552 6426 17564
rect 5445 17527 5503 17533
rect 5445 17493 5457 17527
rect 5491 17524 5503 17527
rect 6822 17524 6828 17536
rect 5491 17496 6828 17524
rect 5491 17493 5503 17496
rect 5445 17487 5503 17493
rect 6822 17484 6828 17496
rect 6880 17484 6886 17536
rect 6932 17524 6960 17564
rect 7193 17561 7205 17595
rect 7239 17592 7251 17595
rect 7374 17592 7380 17604
rect 7239 17564 7380 17592
rect 7239 17561 7251 17564
rect 7193 17555 7251 17561
rect 7374 17552 7380 17564
rect 7432 17552 7438 17604
rect 12060 17595 12118 17601
rect 12060 17561 12072 17595
rect 12106 17592 12118 17595
rect 12342 17592 12348 17604
rect 12106 17564 12348 17592
rect 12106 17561 12118 17564
rect 12060 17555 12118 17561
rect 12342 17552 12348 17564
rect 12400 17552 12406 17604
rect 13722 17552 13728 17604
rect 13780 17592 13786 17604
rect 14277 17595 14335 17601
rect 14277 17592 14289 17595
rect 13780 17564 14289 17592
rect 13780 17552 13786 17564
rect 14277 17561 14289 17564
rect 14323 17561 14335 17595
rect 14642 17592 14648 17604
rect 14603 17564 14648 17592
rect 14277 17555 14335 17561
rect 14642 17552 14648 17564
rect 14700 17552 14706 17604
rect 15013 17595 15071 17601
rect 15013 17561 15025 17595
rect 15059 17592 15071 17595
rect 15194 17592 15200 17604
rect 15059 17564 15200 17592
rect 15059 17561 15071 17564
rect 15013 17555 15071 17561
rect 15194 17552 15200 17564
rect 15252 17552 15258 17604
rect 15832 17595 15890 17601
rect 15832 17561 15844 17595
rect 15878 17592 15890 17595
rect 16850 17592 16856 17604
rect 15878 17564 16856 17592
rect 15878 17561 15890 17564
rect 15832 17555 15890 17561
rect 16850 17552 16856 17564
rect 16908 17552 16914 17604
rect 21634 17552 21640 17604
rect 21692 17592 21698 17604
rect 22465 17595 22523 17601
rect 22465 17592 22477 17595
rect 21692 17564 22477 17592
rect 21692 17552 21698 17564
rect 22465 17561 22477 17564
rect 22511 17561 22523 17595
rect 28166 17592 28172 17604
rect 28127 17564 28172 17592
rect 22465 17555 22523 17561
rect 28166 17552 28172 17564
rect 28224 17552 28230 17604
rect 9950 17524 9956 17536
rect 6932 17496 9956 17524
rect 9950 17484 9956 17496
rect 10008 17484 10014 17536
rect 12986 17484 12992 17536
rect 13044 17524 13050 17536
rect 13173 17527 13231 17533
rect 13173 17524 13185 17527
rect 13044 17496 13185 17524
rect 13044 17484 13050 17496
rect 13173 17493 13185 17496
rect 13219 17493 13231 17527
rect 13173 17487 13231 17493
rect 14366 17484 14372 17536
rect 14424 17524 14430 17536
rect 14461 17527 14519 17533
rect 14461 17524 14473 17527
rect 14424 17496 14473 17524
rect 14424 17484 14430 17496
rect 14461 17493 14473 17496
rect 14507 17493 14519 17527
rect 14461 17487 14519 17493
rect 16945 17527 17003 17533
rect 16945 17493 16957 17527
rect 16991 17524 17003 17527
rect 17218 17524 17224 17536
rect 16991 17496 17224 17524
rect 16991 17493 17003 17496
rect 16945 17487 17003 17493
rect 17218 17484 17224 17496
rect 17276 17484 17282 17536
rect 22097 17527 22155 17533
rect 22097 17493 22109 17527
rect 22143 17524 22155 17527
rect 22278 17524 22284 17536
rect 22143 17496 22284 17524
rect 22143 17493 22155 17496
rect 22097 17487 22155 17493
rect 22278 17484 22284 17496
rect 22336 17484 22342 17536
rect 22557 17527 22615 17533
rect 22557 17493 22569 17527
rect 22603 17524 22615 17527
rect 24026 17524 24032 17536
rect 22603 17496 24032 17524
rect 22603 17493 22615 17496
rect 22557 17487 22615 17493
rect 24026 17484 24032 17496
rect 24084 17484 24090 17536
rect 25130 17484 25136 17536
rect 25188 17524 25194 17536
rect 25314 17524 25320 17536
rect 25188 17496 25320 17524
rect 25188 17484 25194 17496
rect 25314 17484 25320 17496
rect 25372 17524 25378 17536
rect 25961 17527 26019 17533
rect 25961 17524 25973 17527
rect 25372 17496 25973 17524
rect 25372 17484 25378 17496
rect 25961 17493 25973 17496
rect 26007 17493 26019 17527
rect 25961 17487 26019 17493
rect 1104 17434 29048 17456
rect 1104 17382 7896 17434
rect 7948 17382 7960 17434
rect 8012 17382 8024 17434
rect 8076 17382 8088 17434
rect 8140 17382 8152 17434
rect 8204 17382 14842 17434
rect 14894 17382 14906 17434
rect 14958 17382 14970 17434
rect 15022 17382 15034 17434
rect 15086 17382 15098 17434
rect 15150 17382 21788 17434
rect 21840 17382 21852 17434
rect 21904 17382 21916 17434
rect 21968 17382 21980 17434
rect 22032 17382 22044 17434
rect 22096 17382 28734 17434
rect 28786 17382 28798 17434
rect 28850 17382 28862 17434
rect 28914 17382 28926 17434
rect 28978 17382 28990 17434
rect 29042 17382 29048 17434
rect 1104 17360 29048 17382
rect 6730 17320 6736 17332
rect 4448 17292 6736 17320
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17184 2835 17187
rect 2958 17184 2964 17196
rect 2823 17156 2964 17184
rect 2823 17153 2835 17156
rect 2777 17147 2835 17153
rect 2958 17144 2964 17156
rect 3016 17184 3022 17196
rect 4062 17184 4068 17196
rect 3016 17156 4068 17184
rect 3016 17144 3022 17156
rect 4062 17144 4068 17156
rect 4120 17144 4126 17196
rect 4448 17193 4476 17292
rect 6730 17280 6736 17292
rect 6788 17280 6794 17332
rect 14366 17320 14372 17332
rect 13924 17292 14372 17320
rect 13924 17261 13952 17292
rect 14366 17280 14372 17292
rect 14424 17280 14430 17332
rect 16850 17280 16856 17332
rect 16908 17320 16914 17332
rect 16945 17323 17003 17329
rect 16945 17320 16957 17323
rect 16908 17292 16957 17320
rect 16908 17280 16914 17292
rect 16945 17289 16957 17292
rect 16991 17289 17003 17323
rect 27617 17323 27675 17329
rect 16945 17283 17003 17289
rect 22066 17292 24716 17320
rect 13909 17255 13967 17261
rect 13909 17221 13921 17255
rect 13955 17221 13967 17255
rect 14461 17255 14519 17261
rect 14461 17252 14473 17255
rect 13909 17215 13967 17221
rect 14108 17224 14473 17252
rect 5816 17196 5868 17202
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17153 4491 17187
rect 4433 17147 4491 17153
rect 5902 17144 5908 17196
rect 5960 17184 5966 17196
rect 7285 17187 7343 17193
rect 5960 17156 6053 17184
rect 5960 17144 5966 17156
rect 7285 17153 7297 17187
rect 7331 17184 7343 17187
rect 7650 17184 7656 17196
rect 7331 17156 7656 17184
rect 7331 17153 7343 17156
rect 7285 17147 7343 17153
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 10594 17144 10600 17196
rect 10652 17184 10658 17196
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 10652 17156 11713 17184
rect 10652 17144 10658 17156
rect 11701 17153 11713 17156
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 11790 17144 11796 17196
rect 11848 17184 11854 17196
rect 11957 17187 12015 17193
rect 11957 17184 11969 17187
rect 11848 17156 11969 17184
rect 11848 17144 11854 17156
rect 11957 17153 11969 17156
rect 12003 17153 12015 17187
rect 11957 17147 12015 17153
rect 13078 17144 13084 17196
rect 13136 17184 13142 17196
rect 13814 17184 13820 17196
rect 13136 17156 13820 17184
rect 13136 17144 13142 17156
rect 13814 17144 13820 17156
rect 13872 17144 13878 17196
rect 14001 17187 14059 17193
rect 14001 17153 14013 17187
rect 14047 17153 14059 17187
rect 14001 17147 14059 17153
rect 5816 17138 5868 17144
rect 4985 17119 5043 17125
rect 4985 17085 4997 17119
rect 5031 17085 5043 17119
rect 5920 17116 5948 17144
rect 7374 17116 7380 17128
rect 5920 17088 7380 17116
rect 4985 17079 5043 17085
rect 5000 17048 5028 17079
rect 7374 17076 7380 17088
rect 7432 17076 7438 17128
rect 13722 17076 13728 17128
rect 13780 17116 13786 17128
rect 14016 17116 14044 17147
rect 13780 17088 14044 17116
rect 13780 17076 13786 17088
rect 5534 17048 5540 17060
rect 5000 17020 5540 17048
rect 5534 17008 5540 17020
rect 5592 17008 5598 17060
rect 12986 17008 12992 17060
rect 13044 17048 13050 17060
rect 14108 17048 14136 17224
rect 14461 17221 14473 17224
rect 14507 17252 14519 17255
rect 14642 17252 14648 17264
rect 14507 17224 14648 17252
rect 14507 17221 14519 17224
rect 14461 17215 14519 17221
rect 14642 17212 14648 17224
rect 14700 17212 14706 17264
rect 17218 17252 17224 17264
rect 17144 17224 17224 17252
rect 15010 17144 15016 17196
rect 15068 17184 15074 17196
rect 15068 17156 15113 17184
rect 15068 17144 15074 17156
rect 15194 17144 15200 17196
rect 15252 17184 15258 17196
rect 17045 17185 17103 17191
rect 15252 17156 15297 17184
rect 15252 17144 15258 17156
rect 17045 17151 17057 17185
rect 17091 17182 17103 17185
rect 17144 17182 17172 17224
rect 17218 17212 17224 17224
rect 17276 17252 17282 17264
rect 22066 17252 22094 17292
rect 22278 17252 22284 17264
rect 17276 17224 22094 17252
rect 22239 17224 22284 17252
rect 17276 17212 17282 17224
rect 22278 17212 22284 17224
rect 22336 17212 22342 17264
rect 22738 17212 22744 17264
rect 22796 17212 22802 17264
rect 24026 17252 24032 17264
rect 23987 17224 24032 17252
rect 24026 17212 24032 17224
rect 24084 17252 24090 17264
rect 24688 17252 24716 17292
rect 27617 17289 27629 17323
rect 27663 17320 27675 17323
rect 27890 17320 27896 17332
rect 27663 17292 27896 17320
rect 27663 17289 27675 17292
rect 27617 17283 27675 17289
rect 27890 17280 27896 17292
rect 27948 17280 27954 17332
rect 25038 17252 25044 17264
rect 24084 17224 24532 17252
rect 24084 17212 24090 17224
rect 24504 17196 24532 17224
rect 24688 17224 25044 17252
rect 24486 17184 24492 17196
rect 17091 17154 17172 17182
rect 24399 17156 24492 17184
rect 17091 17151 17103 17154
rect 17045 17145 17103 17151
rect 24486 17144 24492 17156
rect 24544 17144 24550 17196
rect 24688 17193 24716 17224
rect 25038 17212 25044 17224
rect 25096 17212 25102 17264
rect 26237 17255 26295 17261
rect 26237 17221 26249 17255
rect 26283 17252 26295 17255
rect 27246 17252 27252 17264
rect 26283 17224 27252 17252
rect 26283 17221 26295 17224
rect 26237 17215 26295 17221
rect 27246 17212 27252 17224
rect 27304 17212 27310 17264
rect 24673 17187 24731 17193
rect 24673 17153 24685 17187
rect 24719 17153 24731 17187
rect 24673 17147 24731 17153
rect 24762 17144 24768 17196
rect 24820 17184 24826 17196
rect 24949 17187 25007 17193
rect 24949 17184 24961 17187
rect 24820 17156 24961 17184
rect 24820 17144 24826 17156
rect 24949 17153 24961 17156
rect 24995 17153 25007 17187
rect 25314 17184 25320 17196
rect 25275 17156 25320 17184
rect 24949 17147 25007 17153
rect 25314 17144 25320 17156
rect 25372 17144 25378 17196
rect 26145 17187 26203 17193
rect 26145 17153 26157 17187
rect 26191 17153 26203 17187
rect 26326 17184 26332 17196
rect 26287 17156 26332 17184
rect 26145 17147 26203 17153
rect 14369 17119 14427 17125
rect 14369 17085 14381 17119
rect 14415 17116 14427 17119
rect 14734 17116 14740 17128
rect 14415 17088 14740 17116
rect 14415 17085 14427 17088
rect 14369 17079 14427 17085
rect 14734 17076 14740 17088
rect 14792 17116 14798 17128
rect 15286 17116 15292 17128
rect 14792 17088 15292 17116
rect 14792 17076 14798 17088
rect 15286 17076 15292 17088
rect 15344 17076 15350 17128
rect 15381 17119 15439 17125
rect 15381 17085 15393 17119
rect 15427 17116 15439 17119
rect 22005 17119 22063 17125
rect 15427 17088 15792 17116
rect 15427 17085 15439 17088
rect 15381 17079 15439 17085
rect 13044 17020 14136 17048
rect 13044 17008 13050 17020
rect 14274 17008 14280 17060
rect 14332 17048 14338 17060
rect 15010 17048 15016 17060
rect 14332 17020 15016 17048
rect 14332 17008 14338 17020
rect 15010 17008 15016 17020
rect 15068 17008 15074 17060
rect 15764 16992 15792 17088
rect 22005 17085 22017 17119
rect 22051 17116 22063 17119
rect 22278 17116 22284 17128
rect 22051 17088 22284 17116
rect 22051 17085 22063 17088
rect 22005 17079 22063 17085
rect 22278 17076 22284 17088
rect 22336 17116 22342 17128
rect 22646 17116 22652 17128
rect 22336 17088 22652 17116
rect 22336 17076 22342 17088
rect 22646 17076 22652 17088
rect 22704 17076 22710 17128
rect 24857 17119 24915 17125
rect 24857 17085 24869 17119
rect 24903 17116 24915 17119
rect 26160 17116 26188 17147
rect 26326 17144 26332 17156
rect 26384 17144 26390 17196
rect 26878 17144 26884 17196
rect 26936 17184 26942 17196
rect 27157 17187 27215 17193
rect 27157 17184 27169 17187
rect 26936 17156 27169 17184
rect 26936 17144 26942 17156
rect 27157 17153 27169 17156
rect 27203 17153 27215 17187
rect 27157 17147 27215 17153
rect 27433 17187 27491 17193
rect 27433 17153 27445 17187
rect 27479 17153 27491 17187
rect 27433 17147 27491 17153
rect 24903 17088 26188 17116
rect 26344 17116 26372 17144
rect 27448 17116 27476 17147
rect 26344 17088 27476 17116
rect 24903 17085 24915 17088
rect 24857 17079 24915 17085
rect 2314 16940 2320 16992
rect 2372 16980 2378 16992
rect 2685 16983 2743 16989
rect 2685 16980 2697 16983
rect 2372 16952 2697 16980
rect 2372 16940 2378 16952
rect 2685 16949 2697 16952
rect 2731 16949 2743 16983
rect 2685 16943 2743 16949
rect 4341 16983 4399 16989
rect 4341 16949 4353 16983
rect 4387 16980 4399 16983
rect 5718 16980 5724 16992
rect 4387 16952 5724 16980
rect 4387 16949 4399 16952
rect 4341 16943 4399 16949
rect 5718 16940 5724 16952
rect 5776 16940 5782 16992
rect 9493 16983 9551 16989
rect 9493 16949 9505 16983
rect 9539 16980 9551 16983
rect 9674 16980 9680 16992
rect 9539 16952 9680 16980
rect 9539 16949 9551 16952
rect 9493 16943 9551 16949
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 13078 16980 13084 16992
rect 13039 16952 13084 16980
rect 13078 16940 13084 16952
rect 13136 16940 13142 16992
rect 14550 16940 14556 16992
rect 14608 16980 14614 16992
rect 15194 16980 15200 16992
rect 14608 16952 15200 16980
rect 14608 16940 14614 16952
rect 15194 16940 15200 16952
rect 15252 16940 15258 16992
rect 15746 16940 15752 16992
rect 15804 16980 15810 16992
rect 18230 16980 18236 16992
rect 15804 16952 18236 16980
rect 15804 16940 15810 16952
rect 18230 16940 18236 16952
rect 18288 16940 18294 16992
rect 1104 16890 28888 16912
rect 1104 16838 4423 16890
rect 4475 16838 4487 16890
rect 4539 16838 4551 16890
rect 4603 16838 4615 16890
rect 4667 16838 4679 16890
rect 4731 16838 11369 16890
rect 11421 16838 11433 16890
rect 11485 16838 11497 16890
rect 11549 16838 11561 16890
rect 11613 16838 11625 16890
rect 11677 16838 18315 16890
rect 18367 16838 18379 16890
rect 18431 16838 18443 16890
rect 18495 16838 18507 16890
rect 18559 16838 18571 16890
rect 18623 16838 25261 16890
rect 25313 16838 25325 16890
rect 25377 16838 25389 16890
rect 25441 16838 25453 16890
rect 25505 16838 25517 16890
rect 25569 16838 28888 16890
rect 1104 16816 28888 16838
rect 8294 16776 8300 16788
rect 8255 16748 8300 16776
rect 8294 16736 8300 16748
rect 8352 16736 8358 16788
rect 10594 16776 10600 16788
rect 9140 16748 10600 16776
rect 6546 16640 6552 16652
rect 6507 16612 6552 16640
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 6822 16640 6828 16652
rect 6783 16612 6828 16640
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 9140 16649 9168 16748
rect 10594 16736 10600 16748
rect 10652 16736 10658 16788
rect 12342 16776 12348 16788
rect 12303 16748 12348 16776
rect 12342 16736 12348 16748
rect 12400 16736 12406 16788
rect 16209 16779 16267 16785
rect 16209 16745 16221 16779
rect 16255 16776 16267 16779
rect 23106 16776 23112 16788
rect 16255 16748 23112 16776
rect 16255 16745 16267 16748
rect 16209 16739 16267 16745
rect 23106 16736 23112 16748
rect 23164 16736 23170 16788
rect 25225 16779 25283 16785
rect 25225 16745 25237 16779
rect 25271 16776 25283 16779
rect 26326 16776 26332 16788
rect 25271 16748 26332 16776
rect 25271 16745 25283 16748
rect 25225 16739 25283 16745
rect 26326 16736 26332 16748
rect 26384 16736 26390 16788
rect 27614 16776 27620 16788
rect 27575 16748 27620 16776
rect 27614 16736 27620 16748
rect 27672 16736 27678 16788
rect 16574 16708 16580 16720
rect 14292 16680 16580 16708
rect 9125 16643 9183 16649
rect 9125 16609 9137 16643
rect 9171 16609 9183 16643
rect 11698 16640 11704 16652
rect 11659 16612 11704 16640
rect 9125 16603 9183 16609
rect 11698 16600 11704 16612
rect 11756 16600 11762 16652
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16640 11943 16643
rect 11931 16612 12434 16640
rect 11931 16609 11943 16612
rect 11885 16603 11943 16609
rect 2501 16575 2559 16581
rect 2501 16541 2513 16575
rect 2547 16572 2559 16575
rect 2590 16572 2596 16584
rect 2547 16544 2596 16572
rect 2547 16541 2559 16544
rect 2501 16535 2559 16541
rect 2590 16532 2596 16544
rect 2648 16532 2654 16584
rect 3234 16532 3240 16584
rect 3292 16572 3298 16584
rect 3329 16575 3387 16581
rect 3329 16572 3341 16575
rect 3292 16544 3341 16572
rect 3292 16532 3298 16544
rect 3329 16541 3341 16544
rect 3375 16541 3387 16575
rect 12250 16572 12256 16584
rect 3329 16535 3387 16541
rect 8128 16544 12256 16572
rect 6932 16476 7314 16504
rect 2038 16396 2044 16448
rect 2096 16436 2102 16448
rect 2409 16439 2467 16445
rect 2409 16436 2421 16439
rect 2096 16408 2421 16436
rect 2096 16396 2102 16408
rect 2409 16405 2421 16408
rect 2455 16405 2467 16439
rect 2409 16399 2467 16405
rect 3237 16439 3295 16445
rect 3237 16405 3249 16439
rect 3283 16436 3295 16439
rect 3326 16436 3332 16448
rect 3283 16408 3332 16436
rect 3283 16405 3295 16408
rect 3237 16399 3295 16405
rect 3326 16396 3332 16408
rect 3384 16396 3390 16448
rect 5534 16396 5540 16448
rect 5592 16436 5598 16448
rect 6932 16436 6960 16476
rect 5592 16408 6960 16436
rect 5592 16396 5598 16408
rect 7006 16396 7012 16448
rect 7064 16436 7070 16448
rect 8128 16436 8156 16544
rect 12250 16532 12256 16544
rect 12308 16532 12314 16584
rect 12406 16572 12434 16612
rect 13078 16600 13084 16652
rect 13136 16640 13142 16652
rect 13633 16643 13691 16649
rect 13633 16640 13645 16643
rect 13136 16612 13645 16640
rect 13136 16600 13142 16612
rect 13633 16609 13645 16612
rect 13679 16609 13691 16643
rect 13633 16603 13691 16609
rect 14182 16600 14188 16652
rect 14240 16640 14246 16652
rect 14292 16640 14320 16680
rect 16574 16668 16580 16680
rect 16632 16668 16638 16720
rect 24026 16708 24032 16720
rect 23939 16680 24032 16708
rect 24026 16668 24032 16680
rect 24084 16708 24090 16720
rect 24673 16711 24731 16717
rect 24673 16708 24685 16711
rect 24084 16680 24685 16708
rect 24084 16668 24090 16680
rect 24673 16677 24685 16680
rect 24719 16708 24731 16711
rect 24762 16708 24768 16720
rect 24719 16680 24768 16708
rect 24719 16677 24731 16680
rect 24673 16671 24731 16677
rect 24762 16668 24768 16680
rect 24820 16668 24826 16720
rect 14642 16640 14648 16652
rect 14240 16612 14320 16640
rect 14603 16612 14648 16640
rect 14240 16600 14246 16612
rect 12986 16572 12992 16584
rect 12406 16544 12992 16572
rect 12986 16532 12992 16544
rect 13044 16532 13050 16584
rect 13170 16572 13176 16584
rect 13131 16544 13176 16572
rect 13170 16532 13176 16544
rect 13228 16532 13234 16584
rect 13722 16572 13728 16584
rect 13280 16544 13728 16572
rect 9214 16464 9220 16516
rect 9272 16504 9278 16516
rect 9370 16507 9428 16513
rect 9370 16504 9382 16507
rect 9272 16476 9382 16504
rect 9272 16464 9278 16476
rect 9370 16473 9382 16476
rect 9416 16473 9428 16507
rect 9370 16467 9428 16473
rect 12894 16464 12900 16516
rect 12952 16504 12958 16516
rect 13081 16507 13139 16513
rect 13081 16504 13093 16507
rect 12952 16476 13093 16504
rect 12952 16464 12958 16476
rect 13081 16473 13093 16476
rect 13127 16504 13139 16507
rect 13280 16504 13308 16544
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 14292 16581 14320 16612
rect 14642 16600 14648 16612
rect 14700 16600 14706 16652
rect 14277 16575 14335 16581
rect 14277 16541 14289 16575
rect 14323 16541 14335 16575
rect 14734 16572 14740 16584
rect 14695 16544 14740 16572
rect 14277 16535 14335 16541
rect 14734 16532 14740 16544
rect 14792 16532 14798 16584
rect 15194 16532 15200 16584
rect 15252 16572 15258 16584
rect 16117 16575 16175 16581
rect 16117 16572 16129 16575
rect 15252 16544 16129 16572
rect 15252 16532 15258 16544
rect 16117 16541 16129 16544
rect 16163 16541 16175 16575
rect 16592 16572 16620 16668
rect 18230 16640 18236 16652
rect 18191 16612 18236 16640
rect 18230 16600 18236 16612
rect 18288 16600 18294 16652
rect 18417 16643 18475 16649
rect 18417 16609 18429 16643
rect 18463 16640 18475 16643
rect 20622 16640 20628 16652
rect 18463 16612 20628 16640
rect 18463 16609 18475 16612
rect 18417 16603 18475 16609
rect 20622 16600 20628 16612
rect 20680 16600 20686 16652
rect 22278 16640 22284 16652
rect 22239 16612 22284 16640
rect 22278 16600 22284 16612
rect 22336 16600 22342 16652
rect 26878 16600 26884 16652
rect 26936 16640 26942 16652
rect 27157 16643 27215 16649
rect 27157 16640 27169 16643
rect 26936 16612 27169 16640
rect 26936 16600 26942 16612
rect 27157 16609 27169 16612
rect 27203 16609 27215 16643
rect 27157 16603 27215 16609
rect 16669 16575 16727 16581
rect 16669 16572 16681 16575
rect 16592 16544 16681 16572
rect 16117 16535 16175 16541
rect 16669 16541 16681 16544
rect 16715 16541 16727 16575
rect 16669 16535 16727 16541
rect 24486 16532 24492 16584
rect 24544 16572 24550 16584
rect 24857 16575 24915 16581
rect 24857 16572 24869 16575
rect 24544 16544 24869 16572
rect 24544 16532 24550 16544
rect 24857 16541 24869 16544
rect 24903 16541 24915 16575
rect 25038 16572 25044 16584
rect 24999 16544 25044 16572
rect 24857 16535 24915 16541
rect 25038 16532 25044 16544
rect 25096 16532 25102 16584
rect 27246 16572 27252 16584
rect 27207 16544 27252 16572
rect 27246 16532 27252 16544
rect 27304 16532 27310 16584
rect 13127 16476 13308 16504
rect 13541 16507 13599 16513
rect 13127 16473 13139 16476
rect 13081 16467 13139 16473
rect 13541 16473 13553 16507
rect 13587 16504 13599 16507
rect 13814 16504 13820 16516
rect 13587 16476 13820 16504
rect 13587 16473 13599 16476
rect 13541 16467 13599 16473
rect 13814 16464 13820 16476
rect 13872 16464 13878 16516
rect 14090 16464 14096 16516
rect 14148 16504 14154 16516
rect 18509 16507 18567 16513
rect 18509 16504 18521 16507
rect 14148 16476 18521 16504
rect 14148 16464 14154 16476
rect 18509 16473 18521 16476
rect 18555 16504 18567 16507
rect 22462 16504 22468 16516
rect 18555 16476 22468 16504
rect 18555 16473 18567 16476
rect 18509 16467 18567 16473
rect 22462 16464 22468 16476
rect 22520 16464 22526 16516
rect 22557 16507 22615 16513
rect 22557 16473 22569 16507
rect 22603 16473 22615 16507
rect 22557 16467 22615 16473
rect 7064 16408 8156 16436
rect 7064 16396 7070 16408
rect 9490 16396 9496 16448
rect 9548 16436 9554 16448
rect 10505 16439 10563 16445
rect 10505 16436 10517 16439
rect 9548 16408 10517 16436
rect 9548 16396 9554 16408
rect 10505 16405 10517 16408
rect 10551 16405 10563 16439
rect 10505 16399 10563 16405
rect 11977 16439 12035 16445
rect 11977 16405 11989 16439
rect 12023 16436 12035 16439
rect 12066 16436 12072 16448
rect 12023 16408 12072 16436
rect 12023 16405 12035 16408
rect 11977 16399 12035 16405
rect 12066 16396 12072 16408
rect 12124 16396 12130 16448
rect 18874 16436 18880 16448
rect 18835 16408 18880 16436
rect 18874 16396 18880 16408
rect 18932 16396 18938 16448
rect 22572 16436 22600 16467
rect 22830 16464 22836 16516
rect 22888 16504 22894 16516
rect 24949 16507 25007 16513
rect 22888 16476 23046 16504
rect 22888 16464 22894 16476
rect 24949 16473 24961 16507
rect 24995 16504 25007 16507
rect 25130 16504 25136 16516
rect 24995 16476 25136 16504
rect 24995 16473 25007 16476
rect 24949 16467 25007 16473
rect 25130 16464 25136 16476
rect 25188 16464 25194 16516
rect 22922 16436 22928 16448
rect 22572 16408 22928 16436
rect 22922 16396 22928 16408
rect 22980 16396 22986 16448
rect 1104 16346 29048 16368
rect 1104 16294 7896 16346
rect 7948 16294 7960 16346
rect 8012 16294 8024 16346
rect 8076 16294 8088 16346
rect 8140 16294 8152 16346
rect 8204 16294 14842 16346
rect 14894 16294 14906 16346
rect 14958 16294 14970 16346
rect 15022 16294 15034 16346
rect 15086 16294 15098 16346
rect 15150 16294 21788 16346
rect 21840 16294 21852 16346
rect 21904 16294 21916 16346
rect 21968 16294 21980 16346
rect 22032 16294 22044 16346
rect 22096 16294 28734 16346
rect 28786 16294 28798 16346
rect 28850 16294 28862 16346
rect 28914 16294 28926 16346
rect 28978 16294 28990 16346
rect 29042 16294 29048 16346
rect 1104 16272 29048 16294
rect 9125 16235 9183 16241
rect 9125 16201 9137 16235
rect 9171 16232 9183 16235
rect 9214 16232 9220 16244
rect 9171 16204 9220 16232
rect 9171 16201 9183 16204
rect 9125 16195 9183 16201
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 9398 16192 9404 16244
rect 9456 16232 9462 16244
rect 9585 16235 9643 16241
rect 9585 16232 9597 16235
rect 9456 16204 9597 16232
rect 9456 16192 9462 16204
rect 9585 16201 9597 16204
rect 9631 16201 9643 16235
rect 9585 16195 9643 16201
rect 11701 16235 11759 16241
rect 11701 16201 11713 16235
rect 11747 16232 11759 16235
rect 11790 16232 11796 16244
rect 11747 16204 11796 16232
rect 11747 16201 11759 16204
rect 11701 16195 11759 16201
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 12161 16235 12219 16241
rect 12161 16201 12173 16235
rect 12207 16232 12219 16235
rect 13078 16232 13084 16244
rect 12207 16204 13084 16232
rect 12207 16201 12219 16204
rect 12161 16195 12219 16201
rect 13078 16192 13084 16204
rect 13136 16192 13142 16244
rect 13446 16232 13452 16244
rect 13407 16204 13452 16232
rect 13446 16192 13452 16204
rect 13504 16192 13510 16244
rect 22557 16235 22615 16241
rect 15672 16204 20714 16232
rect 2314 16164 2320 16176
rect 2275 16136 2320 16164
rect 2314 16124 2320 16136
rect 2372 16124 2378 16176
rect 3326 16124 3332 16176
rect 3384 16124 3390 16176
rect 4062 16164 4068 16176
rect 4023 16136 4068 16164
rect 4062 16124 4068 16136
rect 4120 16124 4126 16176
rect 9306 16124 9312 16176
rect 9364 16164 9370 16176
rect 9493 16167 9551 16173
rect 9493 16164 9505 16167
rect 9364 16136 9505 16164
rect 9364 16124 9370 16136
rect 9493 16133 9505 16136
rect 9539 16133 9551 16167
rect 9493 16127 9551 16133
rect 10704 16136 12204 16164
rect 2038 16096 2044 16108
rect 1999 16068 2044 16096
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 5810 16056 5816 16108
rect 5868 16096 5874 16108
rect 10704 16105 10732 16136
rect 10689 16099 10747 16105
rect 5868 16068 6946 16096
rect 5868 16056 5874 16068
rect 10689 16065 10701 16099
rect 10735 16065 10747 16099
rect 10689 16059 10747 16065
rect 11974 16056 11980 16108
rect 12032 16096 12038 16108
rect 12069 16099 12127 16105
rect 12069 16096 12081 16099
rect 12032 16068 12081 16096
rect 12032 16056 12038 16068
rect 12069 16065 12081 16068
rect 12115 16065 12127 16099
rect 12176 16096 12204 16136
rect 12250 16124 12256 16176
rect 12308 16164 12314 16176
rect 15672 16164 15700 16204
rect 15930 16164 15936 16176
rect 12308 16136 15700 16164
rect 15891 16136 15936 16164
rect 12308 16124 12314 16136
rect 15930 16124 15936 16136
rect 15988 16164 15994 16176
rect 16482 16164 16488 16176
rect 15988 16136 16488 16164
rect 15988 16124 15994 16136
rect 16482 16124 16488 16136
rect 16540 16164 16546 16176
rect 16540 16136 18828 16164
rect 16540 16124 16546 16136
rect 12618 16096 12624 16108
rect 12176 16068 12624 16096
rect 12069 16059 12127 16065
rect 12618 16056 12624 16068
rect 12676 16096 12682 16108
rect 13170 16096 13176 16108
rect 12676 16068 13176 16096
rect 12676 16056 12682 16068
rect 13170 16056 13176 16068
rect 13228 16096 13234 16108
rect 13722 16096 13728 16108
rect 13228 16068 13728 16096
rect 13228 16056 13234 16068
rect 13722 16056 13728 16068
rect 13780 16056 13786 16108
rect 14734 16096 14740 16108
rect 14695 16068 14740 16096
rect 14734 16056 14740 16068
rect 14792 16056 14798 16108
rect 17770 16105 17776 16108
rect 17764 16059 17776 16105
rect 17828 16096 17834 16108
rect 17828 16068 17864 16096
rect 17770 16056 17776 16059
rect 17828 16056 17834 16068
rect 6546 16028 6552 16040
rect 6507 16000 6552 16028
rect 6546 15988 6552 16000
rect 6604 15988 6610 16040
rect 7374 16028 7380 16040
rect 7335 16000 7380 16028
rect 7374 15988 7380 16000
rect 7432 15988 7438 16040
rect 9582 15988 9588 16040
rect 9640 16028 9646 16040
rect 9677 16031 9735 16037
rect 9677 16028 9689 16031
rect 9640 16000 9689 16028
rect 9640 15988 9646 16000
rect 9677 15997 9689 16000
rect 9723 15997 9735 16031
rect 9677 15991 9735 15997
rect 10965 16031 11023 16037
rect 10965 15997 10977 16031
rect 11011 15997 11023 16031
rect 10965 15991 11023 15997
rect 10980 15960 11008 15991
rect 11054 15988 11060 16040
rect 11112 16028 11118 16040
rect 11698 16028 11704 16040
rect 11112 16000 11704 16028
rect 11112 15988 11118 16000
rect 11698 15988 11704 16000
rect 11756 16028 11762 16040
rect 12253 16031 12311 16037
rect 12253 16028 12265 16031
rect 11756 16000 12265 16028
rect 11756 15988 11762 16000
rect 12253 15997 12265 16000
rect 12299 15997 12311 16031
rect 15746 16028 15752 16040
rect 15707 16000 15752 16028
rect 12253 15991 12311 15997
rect 15746 15988 15752 16000
rect 15804 15988 15810 16040
rect 15841 16031 15899 16037
rect 15841 15997 15853 16031
rect 15887 16028 15899 16031
rect 17402 16028 17408 16040
rect 15887 16000 17408 16028
rect 15887 15997 15899 16000
rect 15841 15991 15899 15997
rect 17402 15988 17408 16000
rect 17460 15988 17466 16040
rect 17494 15988 17500 16040
rect 17552 16028 17558 16040
rect 17552 16000 17597 16028
rect 17552 15988 17558 16000
rect 12434 15960 12440 15972
rect 10980 15932 12440 15960
rect 12434 15920 12440 15932
rect 12492 15960 12498 15972
rect 12894 15960 12900 15972
rect 12492 15932 12900 15960
rect 12492 15920 12498 15932
rect 12894 15920 12900 15932
rect 12952 15920 12958 15972
rect 16666 15960 16672 15972
rect 14752 15932 16672 15960
rect 10962 15852 10968 15904
rect 11020 15892 11026 15904
rect 11057 15895 11115 15901
rect 11057 15892 11069 15895
rect 11020 15864 11069 15892
rect 11020 15852 11026 15864
rect 11057 15861 11069 15864
rect 11103 15861 11115 15895
rect 11057 15855 11115 15861
rect 11974 15852 11980 15904
rect 12032 15892 12038 15904
rect 14458 15892 14464 15904
rect 12032 15864 14464 15892
rect 12032 15852 12038 15864
rect 14458 15852 14464 15864
rect 14516 15892 14522 15904
rect 14752 15892 14780 15932
rect 16666 15920 16672 15932
rect 16724 15920 16730 15972
rect 18800 15960 18828 16136
rect 18874 16124 18880 16176
rect 18932 16164 18938 16176
rect 19582 16167 19640 16173
rect 19582 16164 19594 16167
rect 18932 16136 19594 16164
rect 18932 16124 18938 16136
rect 19582 16133 19594 16136
rect 19628 16133 19640 16167
rect 20686 16164 20714 16204
rect 22557 16201 22569 16235
rect 22603 16232 22615 16235
rect 22738 16232 22744 16244
rect 22603 16204 22744 16232
rect 22603 16201 22615 16204
rect 22557 16195 22615 16201
rect 22738 16192 22744 16204
rect 22796 16192 22802 16244
rect 22922 16192 22928 16244
rect 22980 16232 22986 16244
rect 23017 16235 23075 16241
rect 23017 16232 23029 16235
rect 22980 16204 23029 16232
rect 22980 16192 22986 16204
rect 23017 16201 23029 16204
rect 23063 16201 23075 16235
rect 23017 16195 23075 16201
rect 23477 16235 23535 16241
rect 23477 16201 23489 16235
rect 23523 16232 23535 16235
rect 24026 16232 24032 16244
rect 23523 16204 24032 16232
rect 23523 16201 23535 16204
rect 23477 16195 23535 16201
rect 24026 16192 24032 16204
rect 24084 16192 24090 16244
rect 20686 16136 22416 16164
rect 19582 16127 19640 16133
rect 22388 16108 22416 16136
rect 22462 16124 22468 16176
rect 22520 16164 22526 16176
rect 22520 16136 23060 16164
rect 22520 16124 22526 16136
rect 23032 16108 23060 16136
rect 19337 16099 19395 16105
rect 19337 16065 19349 16099
rect 19383 16096 19395 16099
rect 22370 16096 22376 16108
rect 19383 16068 20714 16096
rect 22283 16068 22376 16096
rect 19383 16065 19395 16068
rect 19337 16059 19395 16065
rect 20686 16028 20714 16068
rect 22370 16056 22376 16068
rect 22428 16056 22434 16108
rect 22557 16099 22615 16105
rect 22557 16065 22569 16099
rect 22603 16096 22615 16099
rect 22922 16096 22928 16108
rect 22603 16068 22928 16096
rect 22603 16065 22615 16068
rect 22557 16059 22615 16065
rect 22278 16028 22284 16040
rect 20686 16000 22284 16028
rect 22278 15988 22284 16000
rect 22336 16028 22342 16040
rect 22572 16028 22600 16059
rect 22922 16056 22928 16068
rect 22980 16056 22986 16108
rect 23014 16056 23020 16108
rect 23072 16096 23078 16108
rect 23385 16099 23443 16105
rect 23385 16096 23397 16099
rect 23072 16068 23397 16096
rect 23072 16056 23078 16068
rect 23385 16065 23397 16068
rect 23431 16065 23443 16099
rect 23385 16059 23443 16065
rect 22336 16000 22600 16028
rect 22336 15988 22342 16000
rect 23106 15988 23112 16040
rect 23164 16028 23170 16040
rect 23661 16031 23719 16037
rect 23661 16028 23673 16031
rect 23164 16000 23673 16028
rect 23164 15988 23170 16000
rect 23661 15997 23673 16000
rect 23707 16028 23719 16031
rect 23842 16028 23848 16040
rect 23707 16000 23848 16028
rect 23707 15997 23719 16000
rect 23661 15991 23719 15997
rect 23842 15988 23848 16000
rect 23900 15988 23906 16040
rect 18800 15932 19380 15960
rect 14516 15864 14780 15892
rect 16301 15895 16359 15901
rect 14516 15852 14522 15864
rect 16301 15861 16313 15895
rect 16347 15892 16359 15895
rect 16574 15892 16580 15904
rect 16347 15864 16580 15892
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 16574 15852 16580 15864
rect 16632 15852 16638 15904
rect 18874 15892 18880 15904
rect 18835 15864 18880 15892
rect 18874 15852 18880 15864
rect 18932 15852 18938 15904
rect 19352 15892 19380 15932
rect 20622 15920 20628 15972
rect 20680 15960 20686 15972
rect 20717 15963 20775 15969
rect 20717 15960 20729 15963
rect 20680 15932 20729 15960
rect 20680 15920 20686 15932
rect 20717 15929 20729 15932
rect 20763 15929 20775 15963
rect 20717 15923 20775 15929
rect 21634 15892 21640 15904
rect 19352 15864 21640 15892
rect 21634 15852 21640 15864
rect 21692 15852 21698 15904
rect 1104 15802 28888 15824
rect 1104 15750 4423 15802
rect 4475 15750 4487 15802
rect 4539 15750 4551 15802
rect 4603 15750 4615 15802
rect 4667 15750 4679 15802
rect 4731 15750 11369 15802
rect 11421 15750 11433 15802
rect 11485 15750 11497 15802
rect 11549 15750 11561 15802
rect 11613 15750 11625 15802
rect 11677 15750 18315 15802
rect 18367 15750 18379 15802
rect 18431 15750 18443 15802
rect 18495 15750 18507 15802
rect 18559 15750 18571 15802
rect 18623 15750 25261 15802
rect 25313 15750 25325 15802
rect 25377 15750 25389 15802
rect 25441 15750 25453 15802
rect 25505 15750 25517 15802
rect 25569 15750 28888 15802
rect 1104 15728 28888 15750
rect 7282 15688 7288 15700
rect 7243 15660 7288 15688
rect 7282 15648 7288 15660
rect 7340 15648 7346 15700
rect 17402 15648 17408 15700
rect 17460 15688 17466 15700
rect 17865 15691 17923 15697
rect 17865 15688 17877 15691
rect 17460 15660 17877 15688
rect 17460 15648 17466 15660
rect 17865 15657 17877 15660
rect 17911 15657 17923 15691
rect 22830 15688 22836 15700
rect 22791 15660 22836 15688
rect 17865 15651 17923 15657
rect 22830 15648 22836 15660
rect 22888 15648 22894 15700
rect 11054 15580 11060 15632
rect 11112 15620 11118 15632
rect 14090 15620 14096 15632
rect 11112 15592 14096 15620
rect 11112 15580 11118 15592
rect 14090 15580 14096 15592
rect 14148 15580 14154 15632
rect 4338 15512 4344 15564
rect 4396 15552 4402 15564
rect 4396 15524 9812 15552
rect 4396 15512 4402 15524
rect 1949 15487 2007 15493
rect 1949 15453 1961 15487
rect 1995 15453 2007 15487
rect 2590 15484 2596 15496
rect 2551 15456 2596 15484
rect 1949 15447 2007 15453
rect 1964 15416 1992 15447
rect 2590 15444 2596 15456
rect 2648 15444 2654 15496
rect 3234 15444 3240 15496
rect 3292 15484 3298 15496
rect 3329 15487 3387 15493
rect 3329 15484 3341 15487
rect 3292 15456 3341 15484
rect 3292 15444 3298 15456
rect 3329 15453 3341 15456
rect 3375 15453 3387 15487
rect 5534 15484 5540 15496
rect 5495 15456 5540 15484
rect 3329 15447 3387 15453
rect 5534 15444 5540 15456
rect 5592 15444 5598 15496
rect 9674 15484 9680 15496
rect 9635 15456 9680 15484
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 9784 15484 9812 15524
rect 10962 15512 10968 15564
rect 11020 15552 11026 15564
rect 11333 15555 11391 15561
rect 11333 15552 11345 15555
rect 11020 15524 11345 15552
rect 11020 15512 11026 15524
rect 11333 15521 11345 15524
rect 11379 15521 11391 15555
rect 11333 15515 11391 15521
rect 12434 15512 12440 15564
rect 12492 15552 12498 15564
rect 20349 15555 20407 15561
rect 12492 15524 12537 15552
rect 12492 15512 12498 15524
rect 20349 15521 20361 15555
rect 20395 15552 20407 15555
rect 20530 15552 20536 15564
rect 20395 15524 20536 15552
rect 20395 15521 20407 15524
rect 20349 15515 20407 15521
rect 20530 15512 20536 15524
rect 20588 15512 20594 15564
rect 20625 15555 20683 15561
rect 20625 15521 20637 15555
rect 20671 15552 20683 15555
rect 20898 15552 20904 15564
rect 20671 15524 20904 15552
rect 20671 15521 20683 15524
rect 20625 15515 20683 15521
rect 20898 15512 20904 15524
rect 20956 15512 20962 15564
rect 14277 15487 14335 15493
rect 14277 15484 14289 15487
rect 9784 15456 14289 15484
rect 14277 15453 14289 15456
rect 14323 15453 14335 15487
rect 14277 15447 14335 15453
rect 16485 15487 16543 15493
rect 16485 15453 16497 15487
rect 16531 15453 16543 15487
rect 16485 15447 16543 15453
rect 2774 15416 2780 15428
rect 1964 15388 2780 15416
rect 2774 15376 2780 15388
rect 2832 15376 2838 15428
rect 5718 15376 5724 15428
rect 5776 15416 5782 15428
rect 5813 15419 5871 15425
rect 5813 15416 5825 15419
rect 5776 15388 5825 15416
rect 5776 15376 5782 15388
rect 5813 15385 5825 15388
rect 5859 15385 5871 15419
rect 5813 15379 5871 15385
rect 6546 15376 6552 15428
rect 6604 15376 6610 15428
rect 9950 15416 9956 15428
rect 9911 15388 9956 15416
rect 9950 15376 9956 15388
rect 10008 15376 10014 15428
rect 12618 15416 12624 15428
rect 12579 15388 12624 15416
rect 12618 15376 12624 15388
rect 12676 15376 12682 15428
rect 12802 15416 12808 15428
rect 12763 15388 12808 15416
rect 12802 15376 12808 15388
rect 12860 15376 12866 15428
rect 12986 15376 12992 15428
rect 13044 15416 13050 15428
rect 13173 15419 13231 15425
rect 13173 15416 13185 15419
rect 13044 15388 13185 15416
rect 13044 15376 13050 15388
rect 13173 15385 13185 15388
rect 13219 15416 13231 15419
rect 13262 15416 13268 15428
rect 13219 15388 13268 15416
rect 13219 15385 13231 15388
rect 13173 15379 13231 15385
rect 13262 15376 13268 15388
rect 13320 15376 13326 15428
rect 16500 15416 16528 15447
rect 16574 15444 16580 15496
rect 16632 15484 16638 15496
rect 16741 15487 16799 15493
rect 16741 15484 16753 15487
rect 16632 15456 16753 15484
rect 16632 15444 16638 15456
rect 16741 15453 16753 15456
rect 16787 15453 16799 15487
rect 16741 15447 16799 15453
rect 20257 15487 20315 15493
rect 20257 15453 20269 15487
rect 20303 15484 20315 15487
rect 20714 15484 20720 15496
rect 20303 15456 20720 15484
rect 20303 15453 20315 15456
rect 20257 15447 20315 15453
rect 20714 15444 20720 15456
rect 20772 15444 20778 15496
rect 22370 15444 22376 15496
rect 22428 15484 22434 15496
rect 22741 15487 22799 15493
rect 22741 15484 22753 15487
rect 22428 15456 22753 15484
rect 22428 15444 22434 15456
rect 22741 15453 22753 15456
rect 22787 15453 22799 15487
rect 22922 15484 22928 15496
rect 22883 15456 22928 15484
rect 22741 15447 22799 15453
rect 22922 15444 22928 15456
rect 22980 15444 22986 15496
rect 26142 15484 26148 15496
rect 26103 15456 26148 15484
rect 26142 15444 26148 15456
rect 26200 15444 26206 15496
rect 17494 15416 17500 15428
rect 16500 15388 17500 15416
rect 17494 15376 17500 15388
rect 17552 15376 17558 15428
rect 1854 15348 1860 15360
rect 1815 15320 1860 15348
rect 1854 15308 1860 15320
rect 1912 15308 1918 15360
rect 2498 15348 2504 15360
rect 2459 15320 2504 15348
rect 2498 15308 2504 15320
rect 2556 15308 2562 15360
rect 3234 15348 3240 15360
rect 3195 15320 3240 15348
rect 3234 15308 3240 15320
rect 3292 15308 3298 15360
rect 10502 15308 10508 15360
rect 10560 15348 10566 15360
rect 10781 15351 10839 15357
rect 10781 15348 10793 15351
rect 10560 15320 10793 15348
rect 10560 15308 10566 15320
rect 10781 15317 10793 15320
rect 10827 15317 10839 15351
rect 10781 15311 10839 15317
rect 11054 15308 11060 15360
rect 11112 15348 11118 15360
rect 11149 15351 11207 15357
rect 11149 15348 11161 15351
rect 11112 15320 11161 15348
rect 11112 15308 11118 15320
rect 11149 15317 11161 15320
rect 11195 15317 11207 15351
rect 11149 15311 11207 15317
rect 11238 15308 11244 15360
rect 11296 15348 11302 15360
rect 12713 15351 12771 15357
rect 11296 15320 11341 15348
rect 11296 15308 11302 15320
rect 12713 15317 12725 15351
rect 12759 15348 12771 15351
rect 13446 15348 13452 15360
rect 12759 15320 13452 15348
rect 12759 15317 12771 15320
rect 12713 15311 12771 15317
rect 13446 15308 13452 15320
rect 13504 15308 13510 15360
rect 14734 15308 14740 15360
rect 14792 15348 14798 15360
rect 15565 15351 15623 15357
rect 15565 15348 15577 15351
rect 14792 15320 15577 15348
rect 14792 15308 14798 15320
rect 15565 15317 15577 15320
rect 15611 15317 15623 15351
rect 15565 15311 15623 15317
rect 25958 15308 25964 15360
rect 26016 15348 26022 15360
rect 26053 15351 26111 15357
rect 26053 15348 26065 15351
rect 26016 15320 26065 15348
rect 26016 15308 26022 15320
rect 26053 15317 26065 15320
rect 26099 15317 26111 15351
rect 26053 15311 26111 15317
rect 1104 15258 29048 15280
rect 1104 15206 7896 15258
rect 7948 15206 7960 15258
rect 8012 15206 8024 15258
rect 8076 15206 8088 15258
rect 8140 15206 8152 15258
rect 8204 15206 14842 15258
rect 14894 15206 14906 15258
rect 14958 15206 14970 15258
rect 15022 15206 15034 15258
rect 15086 15206 15098 15258
rect 15150 15206 21788 15258
rect 21840 15206 21852 15258
rect 21904 15206 21916 15258
rect 21968 15206 21980 15258
rect 22032 15206 22044 15258
rect 22096 15206 28734 15258
rect 28786 15206 28798 15258
rect 28850 15206 28862 15258
rect 28914 15206 28926 15258
rect 28978 15206 28990 15258
rect 29042 15206 29048 15258
rect 1104 15184 29048 15206
rect 17770 15104 17776 15156
rect 17828 15144 17834 15156
rect 17865 15147 17923 15153
rect 17865 15144 17877 15147
rect 17828 15116 17877 15144
rect 17828 15104 17834 15116
rect 17865 15113 17877 15116
rect 17911 15113 17923 15147
rect 17865 15107 17923 15113
rect 17954 15104 17960 15156
rect 18012 15144 18018 15156
rect 18233 15147 18291 15153
rect 18233 15144 18245 15147
rect 18012 15116 18245 15144
rect 18012 15104 18018 15116
rect 18233 15113 18245 15116
rect 18279 15113 18291 15147
rect 24946 15144 24952 15156
rect 24907 15116 24952 15144
rect 18233 15107 18291 15113
rect 24946 15104 24952 15116
rect 25004 15104 25010 15156
rect 2225 15079 2283 15085
rect 2225 15045 2237 15079
rect 2271 15076 2283 15079
rect 2498 15076 2504 15088
rect 2271 15048 2504 15076
rect 2271 15045 2283 15048
rect 2225 15039 2283 15045
rect 2498 15036 2504 15048
rect 2556 15036 2562 15088
rect 3234 15036 3240 15088
rect 3292 15036 3298 15088
rect 14921 15079 14979 15085
rect 14921 15076 14933 15079
rect 13372 15048 14933 15076
rect 1854 14968 1860 15020
rect 1912 15008 1918 15020
rect 1949 15011 2007 15017
rect 1949 15008 1961 15011
rect 1912 14980 1961 15008
rect 1912 14968 1918 14980
rect 1949 14977 1961 14980
rect 1995 14977 2007 15011
rect 5074 15008 5080 15020
rect 5035 14980 5080 15008
rect 1949 14971 2007 14977
rect 5074 14968 5080 14980
rect 5132 14968 5138 15020
rect 6546 15008 6552 15020
rect 6507 14980 6552 15008
rect 6546 14968 6552 14980
rect 6604 14968 6610 15020
rect 7466 15008 7472 15020
rect 7427 14980 7472 15008
rect 7466 14968 7472 14980
rect 7524 14968 7530 15020
rect 9944 15011 10002 15017
rect 9944 14977 9956 15011
rect 9990 15008 10002 15011
rect 10410 15008 10416 15020
rect 9990 14980 10416 15008
rect 9990 14977 10002 14980
rect 9944 14971 10002 14977
rect 10410 14968 10416 14980
rect 10468 14968 10474 15020
rect 11238 14968 11244 15020
rect 11296 15008 11302 15020
rect 12342 15008 12348 15020
rect 11296 14980 12348 15008
rect 11296 14968 11302 14980
rect 12342 14968 12348 14980
rect 12400 15008 12406 15020
rect 13372 15017 13400 15048
rect 14921 15045 14933 15048
rect 14967 15045 14979 15079
rect 14921 15039 14979 15045
rect 19260 15048 21404 15076
rect 13357 15011 13415 15017
rect 13357 15008 13369 15011
rect 12400 14980 13369 15008
rect 12400 14968 12406 14980
rect 13357 14977 13369 14980
rect 13403 14977 13415 15011
rect 13357 14971 13415 14977
rect 13446 14968 13452 15020
rect 13504 15008 13510 15020
rect 13504 14980 13549 15008
rect 13504 14968 13510 14980
rect 13722 14968 13728 15020
rect 13780 15008 13786 15020
rect 13909 15011 13967 15017
rect 13909 15008 13921 15011
rect 13780 14980 13921 15008
rect 13780 14968 13786 14980
rect 13909 14977 13921 14980
rect 13955 14977 13967 15011
rect 15013 15011 15071 15017
rect 13909 14971 13967 14977
rect 14016 14980 14780 15008
rect 15013 15006 15025 15011
rect 2590 14900 2596 14952
rect 2648 14940 2654 14952
rect 3973 14943 4031 14949
rect 3973 14940 3985 14943
rect 2648 14912 3985 14940
rect 2648 14900 2654 14912
rect 3973 14909 3985 14912
rect 4019 14909 4031 14943
rect 3973 14903 4031 14909
rect 4801 14943 4859 14949
rect 4801 14909 4813 14943
rect 4847 14940 4859 14943
rect 6564 14940 6592 14968
rect 4847 14912 6592 14940
rect 9677 14943 9735 14949
rect 4847 14909 4859 14912
rect 4801 14903 4859 14909
rect 9677 14909 9689 14943
rect 9723 14909 9735 14943
rect 9677 14903 9735 14909
rect 6638 14804 6644 14816
rect 6599 14776 6644 14804
rect 6638 14764 6644 14776
rect 6696 14764 6702 14816
rect 7558 14804 7564 14816
rect 7519 14776 7564 14804
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 9692 14804 9720 14903
rect 12894 14900 12900 14952
rect 12952 14940 12958 14952
rect 13633 14943 13691 14949
rect 13633 14940 13645 14943
rect 12952 14912 13645 14940
rect 12952 14900 12958 14912
rect 13633 14909 13645 14912
rect 13679 14940 13691 14943
rect 14016 14940 14044 14980
rect 13679 14912 14044 14940
rect 14752 14940 14780 14980
rect 14936 14978 15025 15006
rect 14936 14940 14964 14978
rect 15013 14977 15025 14978
rect 15059 14977 15071 15011
rect 15013 14971 15071 14977
rect 15105 15011 15163 15017
rect 15105 14977 15117 15011
rect 15151 14977 15163 15011
rect 15562 15008 15568 15020
rect 15523 14980 15568 15008
rect 15105 14971 15163 14977
rect 15120 14940 15148 14971
rect 15562 14968 15568 14980
rect 15620 14968 15626 15020
rect 19260 15017 19288 15048
rect 21376 15020 21404 15048
rect 24762 15036 24768 15088
rect 24820 15076 24826 15088
rect 24820 15036 24854 15076
rect 25038 15036 25044 15088
rect 25096 15076 25102 15088
rect 25096 15048 27384 15076
rect 25096 15036 25102 15048
rect 18325 15011 18383 15017
rect 18325 14977 18337 15011
rect 18371 15008 18383 15011
rect 19245 15011 19303 15017
rect 18371 14980 18920 15008
rect 18371 14977 18383 14980
rect 18325 14971 18383 14977
rect 18892 14952 18920 14980
rect 19245 14977 19257 15011
rect 19291 14977 19303 15011
rect 19245 14971 19303 14977
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 21358 15008 21364 15020
rect 20772 14980 20865 15008
rect 21319 14980 21364 15008
rect 20772 14968 20778 14980
rect 21358 14968 21364 14980
rect 21416 14968 21422 15020
rect 24826 15017 24854 15036
rect 24826 15011 24907 15017
rect 24826 14980 24861 15011
rect 24849 14977 24861 14980
rect 24895 15008 24907 15011
rect 26786 15008 26792 15020
rect 24895 14980 24957 15008
rect 26266 14980 26792 15008
rect 24895 14977 24907 14980
rect 24849 14971 24907 14977
rect 26786 14968 26792 14980
rect 26844 14968 26850 15020
rect 27356 15017 27384 15048
rect 27341 15011 27399 15017
rect 27341 14977 27353 15011
rect 27387 15008 27399 15011
rect 27982 15008 27988 15020
rect 27387 14980 27988 15008
rect 27387 14977 27399 14980
rect 27341 14971 27399 14977
rect 27982 14968 27988 14980
rect 28040 14968 28046 15020
rect 14752 14912 14964 14940
rect 15028 14912 15148 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 14274 14872 14280 14884
rect 14235 14844 14280 14872
rect 14274 14832 14280 14844
rect 14332 14872 14338 14884
rect 14826 14872 14832 14884
rect 14332 14844 14832 14872
rect 14332 14832 14338 14844
rect 14826 14832 14832 14844
rect 14884 14832 14890 14884
rect 9950 14804 9956 14816
rect 9692 14776 9956 14804
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 10870 14764 10876 14816
rect 10928 14804 10934 14816
rect 11057 14807 11115 14813
rect 11057 14804 11069 14807
rect 10928 14776 11069 14804
rect 10928 14764 10934 14776
rect 11057 14773 11069 14776
rect 11103 14804 11115 14807
rect 13446 14804 13452 14816
rect 11103 14776 13452 14804
rect 11103 14773 11115 14776
rect 11057 14767 11115 14773
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 13722 14764 13728 14816
rect 13780 14804 13786 14816
rect 15028 14804 15056 14912
rect 15286 14900 15292 14952
rect 15344 14940 15350 14952
rect 15473 14943 15531 14949
rect 15473 14940 15485 14943
rect 15344 14912 15485 14940
rect 15344 14900 15350 14912
rect 15473 14909 15485 14912
rect 15519 14940 15531 14943
rect 16022 14940 16028 14952
rect 15519 14912 16028 14940
rect 15519 14909 15531 14912
rect 15473 14903 15531 14909
rect 16022 14900 16028 14912
rect 16080 14900 16086 14952
rect 18230 14900 18236 14952
rect 18288 14940 18294 14952
rect 18417 14943 18475 14949
rect 18417 14940 18429 14943
rect 18288 14912 18429 14940
rect 18288 14900 18294 14912
rect 18417 14909 18429 14912
rect 18463 14909 18475 14943
rect 18417 14903 18475 14909
rect 18874 14900 18880 14952
rect 18932 14940 18938 14952
rect 19153 14943 19211 14949
rect 19153 14940 19165 14943
rect 18932 14912 19165 14940
rect 18932 14900 18938 14912
rect 19153 14909 19165 14912
rect 19199 14909 19211 14943
rect 20732 14940 20760 14968
rect 25777 14943 25835 14949
rect 20732 14912 24854 14940
rect 19153 14903 19211 14909
rect 19610 14804 19616 14816
rect 13780 14776 15056 14804
rect 19571 14776 19616 14804
rect 13780 14764 13786 14776
rect 19610 14764 19616 14776
rect 19668 14764 19674 14816
rect 20346 14764 20352 14816
rect 20404 14804 20410 14816
rect 20625 14807 20683 14813
rect 20625 14804 20637 14807
rect 20404 14776 20637 14804
rect 20404 14764 20410 14776
rect 20625 14773 20637 14776
rect 20671 14773 20683 14807
rect 21266 14804 21272 14816
rect 21227 14776 21272 14804
rect 20625 14767 20683 14773
rect 21266 14764 21272 14776
rect 21324 14764 21330 14816
rect 24826 14804 24854 14912
rect 25777 14909 25789 14943
rect 25823 14940 25835 14943
rect 26510 14940 26516 14952
rect 25823 14912 26372 14940
rect 26471 14912 26516 14940
rect 25823 14909 25835 14912
rect 25777 14903 25835 14909
rect 26142 14872 26148 14884
rect 25056 14844 26148 14872
rect 25056 14804 25084 14844
rect 26142 14832 26148 14844
rect 26200 14832 26206 14884
rect 26344 14872 26372 14912
rect 26510 14900 26516 14912
rect 26568 14900 26574 14952
rect 27430 14872 27436 14884
rect 26344 14844 27436 14872
rect 27430 14832 27436 14844
rect 27488 14832 27494 14884
rect 27246 14804 27252 14816
rect 24826 14776 25084 14804
rect 27207 14776 27252 14804
rect 27246 14764 27252 14776
rect 27304 14764 27310 14816
rect 1104 14714 28888 14736
rect 1104 14662 4423 14714
rect 4475 14662 4487 14714
rect 4539 14662 4551 14714
rect 4603 14662 4615 14714
rect 4667 14662 4679 14714
rect 4731 14662 11369 14714
rect 11421 14662 11433 14714
rect 11485 14662 11497 14714
rect 11549 14662 11561 14714
rect 11613 14662 11625 14714
rect 11677 14662 18315 14714
rect 18367 14662 18379 14714
rect 18431 14662 18443 14714
rect 18495 14662 18507 14714
rect 18559 14662 18571 14714
rect 18623 14662 25261 14714
rect 25313 14662 25325 14714
rect 25377 14662 25389 14714
rect 25441 14662 25453 14714
rect 25505 14662 25517 14714
rect 25569 14662 28888 14714
rect 1104 14640 28888 14662
rect 5552 14572 8340 14600
rect 5552 14544 5580 14572
rect 5534 14532 5540 14544
rect 2148 14504 5540 14532
rect 2148 14405 2176 14504
rect 5534 14492 5540 14504
rect 5592 14492 5598 14544
rect 6546 14464 6552 14476
rect 5184 14436 6552 14464
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14365 2191 14399
rect 2133 14359 2191 14365
rect 2774 14356 2780 14408
rect 2832 14396 2838 14408
rect 2832 14368 2877 14396
rect 2832 14356 2838 14368
rect 3050 14356 3056 14408
rect 3108 14396 3114 14408
rect 5184 14405 5212 14436
rect 6546 14424 6552 14436
rect 6604 14424 6610 14476
rect 3421 14399 3479 14405
rect 3421 14396 3433 14399
rect 3108 14368 3433 14396
rect 3108 14356 3114 14368
rect 3421 14365 3433 14368
rect 3467 14396 3479 14399
rect 5169 14399 5227 14405
rect 5169 14396 5181 14399
rect 3467 14368 5181 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 5169 14365 5181 14368
rect 5215 14365 5227 14399
rect 5169 14359 5227 14365
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 8312 14405 8340 14572
rect 9582 14560 9588 14612
rect 9640 14600 9646 14612
rect 9640 14572 11192 14600
rect 9640 14560 9646 14572
rect 11164 14532 11192 14572
rect 11238 14560 11244 14612
rect 11296 14600 11302 14612
rect 11609 14603 11667 14609
rect 11609 14600 11621 14603
rect 11296 14572 11621 14600
rect 11296 14560 11302 14572
rect 11609 14569 11621 14572
rect 11655 14569 11667 14603
rect 11609 14563 11667 14569
rect 12437 14603 12495 14609
rect 12437 14569 12449 14603
rect 12483 14600 12495 14603
rect 12802 14600 12808 14612
rect 12483 14572 12808 14600
rect 12483 14569 12495 14572
rect 12437 14563 12495 14569
rect 12802 14560 12808 14572
rect 12860 14560 12866 14612
rect 13446 14560 13452 14612
rect 13504 14600 13510 14612
rect 15562 14600 15568 14612
rect 13504 14572 15568 14600
rect 13504 14560 13510 14572
rect 15562 14560 15568 14572
rect 15620 14560 15626 14612
rect 26142 14560 26148 14612
rect 26200 14600 26206 14612
rect 27433 14603 27491 14609
rect 27433 14600 27445 14603
rect 26200 14572 27445 14600
rect 26200 14560 26206 14572
rect 27433 14569 27445 14572
rect 27479 14569 27491 14603
rect 27433 14563 27491 14569
rect 18690 14532 18696 14544
rect 11164 14504 18696 14532
rect 18690 14492 18696 14504
rect 18748 14492 18754 14544
rect 10502 14464 10508 14476
rect 10463 14436 10508 14464
rect 10502 14424 10508 14436
rect 10560 14424 10566 14476
rect 12894 14424 12900 14476
rect 12952 14464 12958 14476
rect 12989 14467 13047 14473
rect 12989 14464 13001 14467
rect 12952 14436 13001 14464
rect 12952 14424 12958 14436
rect 12989 14433 13001 14436
rect 13035 14433 13047 14467
rect 12989 14427 13047 14433
rect 13725 14467 13783 14473
rect 13725 14433 13737 14467
rect 13771 14464 13783 14467
rect 14182 14464 14188 14476
rect 13771 14436 14188 14464
rect 13771 14433 13783 14436
rect 13725 14427 13783 14433
rect 14182 14424 14188 14436
rect 14240 14464 14246 14476
rect 20346 14464 20352 14476
rect 14240 14436 15700 14464
rect 20307 14436 20352 14464
rect 14240 14424 14246 14436
rect 5629 14399 5687 14405
rect 5629 14396 5641 14399
rect 5592 14368 5641 14396
rect 5592 14356 5598 14368
rect 5629 14365 5641 14368
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14396 8355 14399
rect 9582 14396 9588 14408
rect 8343 14368 9588 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 9582 14356 9588 14368
rect 9640 14356 9646 14408
rect 9950 14356 9956 14408
rect 10008 14396 10014 14408
rect 10229 14399 10287 14405
rect 10229 14396 10241 14399
rect 10008 14368 10241 14396
rect 10008 14356 10014 14368
rect 10229 14365 10241 14368
rect 10275 14365 10287 14399
rect 12342 14396 12348 14408
rect 12303 14368 12348 14396
rect 10229 14359 10287 14365
rect 12342 14356 12348 14368
rect 12400 14396 12406 14408
rect 14461 14399 14519 14405
rect 14461 14396 14473 14399
rect 12400 14368 14473 14396
rect 12400 14356 12406 14368
rect 5902 14328 5908 14340
rect 5863 14300 5908 14328
rect 5902 14288 5908 14300
rect 5960 14288 5966 14340
rect 6638 14288 6644 14340
rect 6696 14288 6702 14340
rect 7466 14288 7472 14340
rect 7524 14328 7530 14340
rect 7653 14331 7711 14337
rect 7653 14328 7665 14331
rect 7524 14300 7665 14328
rect 7524 14288 7530 14300
rect 7653 14297 7665 14300
rect 7699 14297 7711 14331
rect 7653 14291 7711 14297
rect 12618 14288 12624 14340
rect 12676 14328 12682 14340
rect 13372 14337 13400 14368
rect 14461 14365 14473 14368
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 14550 14356 14556 14408
rect 14608 14396 14614 14408
rect 14737 14399 14795 14405
rect 14737 14396 14749 14399
rect 14608 14368 14749 14396
rect 14608 14356 14614 14368
rect 14737 14365 14749 14368
rect 14783 14365 14795 14399
rect 14737 14359 14795 14365
rect 14826 14356 14832 14408
rect 14884 14396 14890 14408
rect 15672 14405 15700 14436
rect 20346 14424 20352 14436
rect 20404 14424 20410 14476
rect 20625 14467 20683 14473
rect 20625 14433 20637 14467
rect 20671 14464 20683 14467
rect 21266 14464 21272 14476
rect 20671 14436 21272 14464
rect 20671 14433 20683 14436
rect 20625 14427 20683 14433
rect 21266 14424 21272 14436
rect 21324 14424 21330 14476
rect 21358 14424 21364 14476
rect 21416 14464 21422 14476
rect 22373 14467 22431 14473
rect 22373 14464 22385 14467
rect 21416 14436 22385 14464
rect 21416 14424 21422 14436
rect 22373 14433 22385 14436
rect 22419 14433 22431 14467
rect 22373 14427 22431 14433
rect 24946 14424 24952 14476
rect 25004 14464 25010 14476
rect 25685 14467 25743 14473
rect 25685 14464 25697 14467
rect 25004 14436 25697 14464
rect 25004 14424 25010 14436
rect 25685 14433 25697 14436
rect 25731 14433 25743 14467
rect 25958 14464 25964 14476
rect 25919 14436 25964 14464
rect 25685 14427 25743 14433
rect 25958 14424 25964 14436
rect 26016 14424 26022 14476
rect 15473 14399 15531 14405
rect 14884 14368 14929 14396
rect 14884 14356 14890 14368
rect 15473 14365 15485 14399
rect 15519 14365 15531 14399
rect 15473 14359 15531 14365
rect 15657 14399 15715 14405
rect 15657 14365 15669 14399
rect 15703 14365 15715 14399
rect 15657 14359 15715 14365
rect 13173 14331 13231 14337
rect 13173 14328 13185 14331
rect 12676 14300 13185 14328
rect 12676 14288 12682 14300
rect 13173 14297 13185 14300
rect 13219 14297 13231 14331
rect 13173 14291 13231 14297
rect 13357 14331 13415 14337
rect 13357 14297 13369 14331
rect 13403 14297 13415 14331
rect 13357 14291 13415 14297
rect 13814 14288 13820 14340
rect 13872 14328 13878 14340
rect 14366 14328 14372 14340
rect 13872 14300 14372 14328
rect 13872 14288 13878 14300
rect 14366 14288 14372 14300
rect 14424 14328 14430 14340
rect 14645 14331 14703 14337
rect 14645 14328 14657 14331
rect 14424 14300 14657 14328
rect 14424 14288 14430 14300
rect 14645 14297 14657 14300
rect 14691 14328 14703 14331
rect 15488 14328 15516 14359
rect 14691 14300 15516 14328
rect 15841 14331 15899 14337
rect 14691 14297 14703 14300
rect 14645 14291 14703 14297
rect 15841 14297 15853 14331
rect 15887 14328 15899 14331
rect 17494 14328 17500 14340
rect 15887 14300 17500 14328
rect 15887 14297 15899 14300
rect 15841 14291 15899 14297
rect 17494 14288 17500 14300
rect 17552 14288 17558 14340
rect 21174 14288 21180 14340
rect 21232 14288 21238 14340
rect 26510 14288 26516 14340
rect 26568 14288 26574 14340
rect 1578 14220 1584 14272
rect 1636 14260 1642 14272
rect 2041 14263 2099 14269
rect 2041 14260 2053 14263
rect 1636 14232 2053 14260
rect 1636 14220 1642 14232
rect 2041 14229 2053 14232
rect 2087 14229 2099 14263
rect 2041 14223 2099 14229
rect 2314 14220 2320 14272
rect 2372 14260 2378 14272
rect 2685 14263 2743 14269
rect 2685 14260 2697 14263
rect 2372 14232 2697 14260
rect 2372 14220 2378 14232
rect 2685 14229 2697 14232
rect 2731 14229 2743 14263
rect 3326 14260 3332 14272
rect 3287 14232 3332 14260
rect 2685 14223 2743 14229
rect 3326 14220 3332 14232
rect 3384 14220 3390 14272
rect 5074 14260 5080 14272
rect 5035 14232 5080 14260
rect 5074 14220 5080 14232
rect 5132 14220 5138 14272
rect 8202 14260 8208 14272
rect 8163 14232 8208 14260
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 13265 14263 13323 14269
rect 13265 14229 13277 14263
rect 13311 14260 13323 14263
rect 13446 14260 13452 14272
rect 13311 14232 13452 14260
rect 13311 14229 13323 14232
rect 13265 14223 13323 14229
rect 13446 14220 13452 14232
rect 13504 14220 13510 14272
rect 15013 14263 15071 14269
rect 15013 14229 15025 14263
rect 15059 14260 15071 14263
rect 15654 14260 15660 14272
rect 15059 14232 15660 14260
rect 15059 14229 15071 14232
rect 15013 14223 15071 14229
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 17218 14220 17224 14272
rect 17276 14260 17282 14272
rect 20714 14260 20720 14272
rect 17276 14232 20720 14260
rect 17276 14220 17282 14232
rect 20714 14220 20720 14232
rect 20772 14220 20778 14272
rect 1104 14170 29048 14192
rect 1104 14118 7896 14170
rect 7948 14118 7960 14170
rect 8012 14118 8024 14170
rect 8076 14118 8088 14170
rect 8140 14118 8152 14170
rect 8204 14118 14842 14170
rect 14894 14118 14906 14170
rect 14958 14118 14970 14170
rect 15022 14118 15034 14170
rect 15086 14118 15098 14170
rect 15150 14118 21788 14170
rect 21840 14118 21852 14170
rect 21904 14118 21916 14170
rect 21968 14118 21980 14170
rect 22032 14118 22044 14170
rect 22096 14118 28734 14170
rect 28786 14118 28798 14170
rect 28850 14118 28862 14170
rect 28914 14118 28926 14170
rect 28978 14118 28990 14170
rect 29042 14118 29048 14170
rect 1104 14096 29048 14118
rect 5534 14056 5540 14068
rect 5495 14028 5540 14056
rect 5534 14016 5540 14028
rect 5592 14016 5598 14068
rect 5902 14016 5908 14068
rect 5960 14056 5966 14068
rect 6641 14059 6699 14065
rect 6641 14056 6653 14059
rect 5960 14028 6653 14056
rect 5960 14016 5966 14028
rect 6641 14025 6653 14028
rect 6687 14025 6699 14059
rect 6641 14019 6699 14025
rect 9582 14016 9588 14068
rect 9640 14056 9646 14068
rect 9677 14059 9735 14065
rect 9677 14056 9689 14059
rect 9640 14028 9689 14056
rect 9640 14016 9646 14028
rect 9677 14025 9689 14028
rect 9723 14025 9735 14059
rect 10410 14056 10416 14068
rect 10371 14028 10416 14056
rect 9677 14019 9735 14025
rect 10410 14016 10416 14028
rect 10468 14016 10474 14068
rect 10870 14056 10876 14068
rect 10831 14028 10876 14056
rect 10870 14016 10876 14028
rect 10928 14016 10934 14068
rect 14274 14056 14280 14068
rect 12912 14028 14280 14056
rect 2314 13988 2320 14000
rect 2275 13960 2320 13988
rect 2314 13948 2320 13960
rect 2372 13948 2378 14000
rect 3326 13948 3332 14000
rect 3384 13948 3390 14000
rect 8202 13988 8208 14000
rect 8163 13960 8208 13988
rect 8202 13948 8208 13960
rect 8260 13948 8266 14000
rect 9858 13988 9864 14000
rect 9430 13960 9864 13988
rect 9858 13948 9864 13960
rect 9916 13948 9922 14000
rect 4798 13920 4804 13932
rect 4759 13892 4804 13920
rect 4798 13880 4804 13892
rect 4856 13920 4862 13932
rect 5445 13923 5503 13929
rect 5445 13920 5457 13923
rect 4856 13892 5457 13920
rect 4856 13880 4862 13892
rect 5445 13889 5457 13892
rect 5491 13889 5503 13923
rect 5445 13883 5503 13889
rect 6733 13923 6791 13929
rect 6733 13889 6745 13923
rect 6779 13920 6791 13923
rect 7466 13920 7472 13932
rect 6779 13892 7472 13920
rect 6779 13889 6791 13892
rect 6733 13883 6791 13889
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 7558 13880 7564 13932
rect 7616 13920 7622 13932
rect 7929 13923 7987 13929
rect 7929 13920 7941 13923
rect 7616 13892 7941 13920
rect 7616 13880 7622 13892
rect 7929 13889 7941 13892
rect 7975 13889 7987 13923
rect 10778 13920 10784 13932
rect 10739 13892 10784 13920
rect 7929 13883 7987 13889
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 12158 13920 12164 13932
rect 12119 13892 12164 13920
rect 12158 13880 12164 13892
rect 12216 13880 12222 13932
rect 12912 13929 12940 14028
rect 14274 14016 14280 14028
rect 14332 14016 14338 14068
rect 14737 14059 14795 14065
rect 14737 14025 14749 14059
rect 14783 14056 14795 14059
rect 15378 14056 15384 14068
rect 14783 14028 15384 14056
rect 14783 14025 14795 14028
rect 14737 14019 14795 14025
rect 15378 14016 15384 14028
rect 15436 14016 15442 14068
rect 24762 14056 24768 14068
rect 20686 14028 24768 14056
rect 13446 13948 13452 14000
rect 13504 13988 13510 14000
rect 15749 13991 15807 13997
rect 15749 13988 15761 13991
rect 13504 13960 15761 13988
rect 13504 13948 13510 13960
rect 15749 13957 15761 13960
rect 15795 13957 15807 13991
rect 15749 13951 15807 13957
rect 16042 13991 16100 13997
rect 16042 13957 16054 13991
rect 16088 13988 16100 13991
rect 17218 13988 17224 14000
rect 16088 13960 17224 13988
rect 16088 13957 16100 13960
rect 16042 13951 16100 13957
rect 17218 13948 17224 13960
rect 17276 13948 17282 14000
rect 20686 13988 20714 14028
rect 24762 14016 24768 14028
rect 24820 14016 24826 14068
rect 17696 13960 18276 13988
rect 12897 13923 12955 13929
rect 12897 13889 12909 13923
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 13624 13923 13682 13929
rect 13624 13889 13636 13923
rect 13670 13920 13682 13923
rect 14182 13920 14188 13932
rect 13670 13892 14188 13920
rect 13670 13889 13682 13892
rect 13624 13883 13682 13889
rect 14182 13880 14188 13892
rect 14240 13880 14246 13932
rect 15470 13920 15476 13932
rect 14384 13892 15476 13920
rect 2038 13852 2044 13864
rect 1999 13824 2044 13852
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 2774 13812 2780 13864
rect 2832 13852 2838 13864
rect 4065 13855 4123 13861
rect 4065 13852 4077 13855
rect 2832 13824 4077 13852
rect 2832 13812 2838 13824
rect 4065 13821 4077 13824
rect 4111 13821 4123 13855
rect 4065 13815 4123 13821
rect 4893 13855 4951 13861
rect 4893 13821 4905 13855
rect 4939 13852 4951 13855
rect 5810 13852 5816 13864
rect 4939 13824 5816 13852
rect 4939 13821 4951 13824
rect 4893 13815 4951 13821
rect 5810 13812 5816 13824
rect 5868 13812 5874 13864
rect 10962 13852 10968 13864
rect 10923 13824 10968 13852
rect 10962 13812 10968 13824
rect 11020 13812 11026 13864
rect 12529 13855 12587 13861
rect 12529 13821 12541 13855
rect 12575 13852 12587 13855
rect 12618 13852 12624 13864
rect 12575 13824 12624 13852
rect 12575 13821 12587 13824
rect 12529 13815 12587 13821
rect 12618 13812 12624 13824
rect 12676 13812 12682 13864
rect 13357 13855 13415 13861
rect 13357 13821 13369 13855
rect 13403 13821 13415 13855
rect 13357 13815 13415 13821
rect 13372 13728 13400 13815
rect 13354 13716 13360 13728
rect 13267 13688 13360 13716
rect 13354 13676 13360 13688
rect 13412 13716 13418 13728
rect 14384 13716 14412 13892
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 15654 13920 15660 13932
rect 15615 13892 15660 13920
rect 15654 13880 15660 13892
rect 15712 13880 15718 13932
rect 15893 13923 15951 13929
rect 15893 13889 15905 13923
rect 15939 13920 15951 13923
rect 17313 13923 17371 13929
rect 15939 13892 17264 13920
rect 15939 13889 15951 13892
rect 15893 13883 15951 13889
rect 17236 13852 17264 13892
rect 17313 13889 17325 13923
rect 17359 13920 17371 13923
rect 17402 13920 17408 13932
rect 17359 13892 17408 13920
rect 17359 13889 17371 13892
rect 17313 13883 17371 13889
rect 17402 13880 17408 13892
rect 17460 13880 17466 13932
rect 17497 13923 17555 13929
rect 17696 13926 17724 13960
rect 17497 13889 17509 13923
rect 17543 13920 17555 13923
rect 17604 13920 17724 13926
rect 17543 13898 17724 13920
rect 17543 13892 17632 13898
rect 17543 13889 17555 13892
rect 17497 13883 17555 13889
rect 17770 13880 17776 13932
rect 17828 13920 17834 13932
rect 18141 13923 18199 13929
rect 18141 13920 18153 13923
rect 17828 13892 18153 13920
rect 17828 13880 17834 13892
rect 18141 13889 18153 13892
rect 18187 13889 18199 13923
rect 18248 13920 18276 13960
rect 19260 13960 20714 13988
rect 18325 13923 18383 13929
rect 18325 13920 18337 13923
rect 18248 13892 18337 13920
rect 18141 13883 18199 13889
rect 18325 13889 18337 13892
rect 18371 13920 18383 13923
rect 19260 13920 19288 13960
rect 21174 13948 21180 14000
rect 21232 13988 21238 14000
rect 21232 13960 21277 13988
rect 21232 13948 21238 13960
rect 27798 13948 27804 14000
rect 27856 13988 27862 14000
rect 27985 13991 28043 13997
rect 27985 13988 27997 13991
rect 27856 13960 27997 13988
rect 27856 13948 27862 13960
rect 27985 13957 27997 13960
rect 28031 13957 28043 13991
rect 27985 13951 28043 13957
rect 27344 13932 27396 13938
rect 21450 13920 21456 13932
rect 18371 13892 19288 13920
rect 21114 13892 21456 13920
rect 18371 13889 18383 13892
rect 18325 13883 18383 13889
rect 21450 13880 21456 13892
rect 21508 13880 21514 13932
rect 21542 13880 21548 13932
rect 21600 13920 21606 13932
rect 23106 13929 23112 13932
rect 22833 13923 22891 13929
rect 22833 13920 22845 13923
rect 21600 13892 22845 13920
rect 21600 13880 21606 13892
rect 22833 13889 22845 13892
rect 22879 13889 22891 13923
rect 22833 13883 22891 13889
rect 23100 13883 23112 13929
rect 23164 13920 23170 13932
rect 26418 13920 26424 13932
rect 23164 13892 23200 13920
rect 26379 13892 26424 13920
rect 23106 13880 23112 13883
rect 23164 13880 23170 13892
rect 26418 13880 26424 13892
rect 26476 13880 26482 13932
rect 26786 13880 26792 13932
rect 26844 13920 26850 13932
rect 26844 13892 27344 13920
rect 26844 13880 26850 13892
rect 17420 13852 17448 13880
rect 17586 13852 17592 13864
rect 17236 13824 17356 13852
rect 17420 13824 17592 13852
rect 17328 13784 17356 13824
rect 17586 13812 17592 13824
rect 17644 13812 17650 13864
rect 17681 13855 17739 13861
rect 17681 13821 17693 13855
rect 17727 13852 17739 13855
rect 17954 13852 17960 13864
rect 17727 13824 17960 13852
rect 17727 13821 17739 13824
rect 17681 13815 17739 13821
rect 17954 13812 17960 13824
rect 18012 13812 18018 13864
rect 19426 13852 19432 13864
rect 18064 13824 19432 13852
rect 18064 13784 18092 13824
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 20622 13852 20628 13864
rect 20535 13824 20628 13852
rect 20622 13812 20628 13824
rect 20680 13852 20686 13864
rect 20806 13852 20812 13864
rect 20680 13824 20812 13852
rect 20680 13812 20686 13824
rect 20806 13812 20812 13824
rect 20864 13812 20870 13864
rect 17328 13756 18092 13784
rect 21082 13744 21088 13796
rect 21140 13784 21146 13796
rect 21560 13784 21588 13880
rect 27344 13874 27396 13880
rect 27430 13812 27436 13864
rect 27488 13852 27494 13864
rect 27488 13824 27533 13852
rect 27488 13812 27494 13824
rect 21140 13756 21588 13784
rect 21140 13744 21146 13756
rect 18230 13716 18236 13728
rect 13412 13688 14412 13716
rect 18191 13688 18236 13716
rect 13412 13676 13418 13688
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 23566 13676 23572 13728
rect 23624 13716 23630 13728
rect 24213 13719 24271 13725
rect 24213 13716 24225 13719
rect 23624 13688 24225 13716
rect 23624 13676 23630 13688
rect 24213 13685 24225 13688
rect 24259 13685 24271 13719
rect 24213 13679 24271 13685
rect 26234 13676 26240 13728
rect 26292 13716 26298 13728
rect 26329 13719 26387 13725
rect 26329 13716 26341 13719
rect 26292 13688 26341 13716
rect 26292 13676 26298 13688
rect 26329 13685 26341 13688
rect 26375 13685 26387 13719
rect 26329 13679 26387 13685
rect 1104 13626 28888 13648
rect 1104 13574 4423 13626
rect 4475 13574 4487 13626
rect 4539 13574 4551 13626
rect 4603 13574 4615 13626
rect 4667 13574 4679 13626
rect 4731 13574 11369 13626
rect 11421 13574 11433 13626
rect 11485 13574 11497 13626
rect 11549 13574 11561 13626
rect 11613 13574 11625 13626
rect 11677 13574 18315 13626
rect 18367 13574 18379 13626
rect 18431 13574 18443 13626
rect 18495 13574 18507 13626
rect 18559 13574 18571 13626
rect 18623 13574 25261 13626
rect 25313 13574 25325 13626
rect 25377 13574 25389 13626
rect 25441 13574 25453 13626
rect 25505 13574 25517 13626
rect 25569 13574 28888 13626
rect 1104 13552 28888 13574
rect 2038 13472 2044 13524
rect 2096 13512 2102 13524
rect 2317 13515 2375 13521
rect 2317 13512 2329 13515
rect 2096 13484 2329 13512
rect 2096 13472 2102 13484
rect 2317 13481 2329 13484
rect 2363 13481 2375 13515
rect 10873 13515 10931 13521
rect 10873 13512 10885 13515
rect 2317 13475 2375 13481
rect 6564 13484 10885 13512
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13376 4123 13379
rect 4798 13376 4804 13388
rect 4111 13348 4804 13376
rect 4111 13345 4123 13348
rect 4065 13339 4123 13345
rect 4798 13336 4804 13348
rect 4856 13336 4862 13388
rect 5810 13376 5816 13388
rect 5771 13348 5816 13376
rect 5810 13336 5816 13348
rect 5868 13336 5874 13388
rect 6089 13379 6147 13385
rect 6089 13345 6101 13379
rect 6135 13376 6147 13379
rect 6564 13376 6592 13484
rect 10873 13481 10885 13484
rect 10919 13481 10931 13515
rect 23106 13512 23112 13524
rect 23067 13484 23112 13512
rect 10873 13475 10931 13481
rect 23106 13472 23112 13484
rect 23164 13472 23170 13524
rect 27982 13512 27988 13524
rect 27943 13484 27988 13512
rect 27982 13472 27988 13484
rect 28040 13472 28046 13524
rect 9858 13444 9864 13456
rect 9819 13416 9864 13444
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 14642 13444 14648 13456
rect 11716 13416 14648 13444
rect 6135 13348 6592 13376
rect 6135 13345 6147 13348
rect 6089 13339 6147 13345
rect 11716 13320 11744 13416
rect 14642 13404 14648 13416
rect 14700 13404 14706 13456
rect 23584 13416 24900 13444
rect 23584 13388 23612 13416
rect 12621 13379 12679 13385
rect 12621 13376 12633 13379
rect 11808 13348 12633 13376
rect 1765 13311 1823 13317
rect 1765 13277 1777 13311
rect 1811 13308 1823 13311
rect 2409 13311 2467 13317
rect 2409 13308 2421 13311
rect 1811 13280 2421 13308
rect 1811 13277 1823 13280
rect 1765 13271 1823 13277
rect 2409 13277 2421 13280
rect 2455 13277 2467 13311
rect 3050 13308 3056 13320
rect 3011 13280 3056 13308
rect 2409 13271 2467 13277
rect 2424 13240 2452 13271
rect 3050 13268 3056 13280
rect 3108 13268 3114 13320
rect 6546 13308 6552 13320
rect 6507 13280 6552 13308
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 9769 13311 9827 13317
rect 9769 13277 9781 13311
rect 9815 13308 9827 13311
rect 9950 13308 9956 13320
rect 9815 13280 9956 13308
rect 9815 13277 9827 13280
rect 9769 13271 9827 13277
rect 9950 13268 9956 13280
rect 10008 13268 10014 13320
rect 10962 13308 10968 13320
rect 10923 13280 10968 13308
rect 10962 13268 10968 13280
rect 11020 13268 11026 13320
rect 11698 13308 11704 13320
rect 11659 13280 11704 13308
rect 11698 13268 11704 13280
rect 11756 13268 11762 13320
rect 3602 13240 3608 13252
rect 2424 13212 3608 13240
rect 3602 13200 3608 13212
rect 3660 13200 3666 13252
rect 5074 13200 5080 13252
rect 5132 13200 5138 13252
rect 6638 13200 6644 13252
rect 6696 13240 6702 13252
rect 6794 13243 6852 13249
rect 6794 13240 6806 13243
rect 6696 13212 6806 13240
rect 6696 13200 6702 13212
rect 6794 13209 6806 13212
rect 6840 13209 6852 13243
rect 6794 13203 6852 13209
rect 7190 13200 7196 13252
rect 7248 13240 7254 13252
rect 9306 13240 9312 13252
rect 7248 13212 9312 13240
rect 7248 13200 7254 13212
rect 9306 13200 9312 13212
rect 9364 13240 9370 13252
rect 11808 13240 11836 13348
rect 12621 13345 12633 13348
rect 12667 13345 12679 13379
rect 23566 13376 23572 13388
rect 12621 13339 12679 13345
rect 12728 13348 14412 13376
rect 12158 13308 12164 13320
rect 12119 13280 12164 13308
rect 12158 13268 12164 13280
rect 12216 13308 12222 13320
rect 12728 13317 12756 13348
rect 14384 13320 14412 13348
rect 16776 13348 19840 13376
rect 23527 13348 23572 13376
rect 12713 13311 12771 13317
rect 12713 13308 12725 13311
rect 12216 13280 12725 13308
rect 12216 13268 12222 13280
rect 12713 13277 12725 13280
rect 12759 13277 12771 13311
rect 12986 13308 12992 13320
rect 12947 13280 12992 13308
rect 12713 13271 12771 13277
rect 12986 13268 12992 13280
rect 13044 13268 13050 13320
rect 14366 13268 14372 13320
rect 14424 13308 14430 13320
rect 14645 13311 14703 13317
rect 14645 13308 14657 13311
rect 14424 13280 14657 13308
rect 14424 13268 14430 13280
rect 14645 13277 14657 13280
rect 14691 13277 14703 13311
rect 14645 13271 14703 13277
rect 14921 13311 14979 13317
rect 14921 13277 14933 13311
rect 14967 13308 14979 13311
rect 15286 13308 15292 13320
rect 14967 13280 15292 13308
rect 14967 13277 14979 13280
rect 14921 13271 14979 13277
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 15749 13311 15807 13317
rect 15749 13308 15761 13311
rect 15528 13280 15761 13308
rect 15528 13268 15534 13280
rect 15749 13277 15761 13280
rect 15795 13308 15807 13311
rect 16482 13308 16488 13320
rect 15795 13280 16488 13308
rect 15795 13277 15807 13280
rect 15749 13271 15807 13277
rect 16482 13268 16488 13280
rect 16540 13308 16546 13320
rect 16776 13308 16804 13348
rect 17586 13308 17592 13320
rect 16540 13280 16804 13308
rect 17547 13280 17592 13308
rect 16540 13268 16546 13280
rect 17586 13268 17592 13280
rect 17644 13268 17650 13320
rect 17678 13268 17684 13320
rect 17736 13308 17742 13320
rect 17954 13308 17960 13320
rect 17736 13280 17781 13308
rect 17915 13280 17960 13308
rect 17736 13268 17742 13280
rect 17954 13268 17960 13280
rect 18012 13268 18018 13320
rect 18095 13311 18153 13317
rect 18095 13277 18107 13311
rect 18141 13308 18153 13311
rect 18230 13308 18236 13320
rect 18141 13280 18236 13308
rect 18141 13277 18153 13280
rect 18095 13271 18153 13277
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 19518 13308 19524 13320
rect 19479 13280 19524 13308
rect 19518 13268 19524 13280
rect 19576 13268 19582 13320
rect 19705 13311 19763 13317
rect 19705 13277 19717 13311
rect 19751 13277 19763 13311
rect 19705 13271 19763 13277
rect 9364 13212 11836 13240
rect 12069 13243 12127 13249
rect 9364 13200 9370 13212
rect 12069 13209 12081 13243
rect 12115 13240 12127 13243
rect 12802 13240 12808 13252
rect 12115 13212 12808 13240
rect 12115 13209 12127 13212
rect 12069 13203 12127 13209
rect 12802 13200 12808 13212
rect 12860 13200 12866 13252
rect 14553 13243 14611 13249
rect 14553 13209 14565 13243
rect 14599 13240 14611 13243
rect 16016 13243 16074 13249
rect 14599 13212 14688 13240
rect 14599 13209 14611 13212
rect 14553 13203 14611 13209
rect 14660 13184 14688 13212
rect 16016 13209 16028 13243
rect 16062 13240 16074 13243
rect 16850 13240 16856 13252
rect 16062 13212 16856 13240
rect 16062 13209 16074 13212
rect 16016 13203 16074 13209
rect 16850 13200 16856 13212
rect 16908 13200 16914 13252
rect 17034 13200 17040 13252
rect 17092 13240 17098 13252
rect 17865 13243 17923 13249
rect 17865 13240 17877 13243
rect 17092 13212 17877 13240
rect 17092 13200 17098 13212
rect 17865 13209 17877 13212
rect 17911 13209 17923 13243
rect 19720 13240 19748 13271
rect 17865 13203 17923 13209
rect 18248 13212 19748 13240
rect 19812 13240 19840 13348
rect 23566 13336 23572 13348
rect 23624 13336 23630 13388
rect 23750 13376 23756 13388
rect 23711 13348 23756 13376
rect 23750 13336 23756 13348
rect 23808 13336 23814 13388
rect 24578 13376 24584 13388
rect 24539 13348 24584 13376
rect 24578 13336 24584 13348
rect 24636 13336 24642 13388
rect 24872 13385 24900 13416
rect 24857 13379 24915 13385
rect 24857 13345 24869 13379
rect 24903 13345 24915 13379
rect 26234 13376 26240 13388
rect 26195 13348 26240 13376
rect 24857 13339 24915 13345
rect 26234 13336 26240 13348
rect 26292 13336 26298 13388
rect 26513 13379 26571 13385
rect 26513 13345 26525 13379
rect 26559 13376 26571 13379
rect 27246 13376 27252 13388
rect 26559 13348 27252 13376
rect 26559 13345 26571 13348
rect 26513 13339 26571 13345
rect 27246 13336 27252 13348
rect 27304 13336 27310 13388
rect 19889 13311 19947 13317
rect 19889 13277 19901 13311
rect 19935 13308 19947 13311
rect 20990 13308 20996 13320
rect 19935 13280 20996 13308
rect 19935 13277 19947 13280
rect 19889 13271 19947 13277
rect 20990 13268 20996 13280
rect 21048 13268 21054 13320
rect 23474 13308 23480 13320
rect 23435 13280 23480 13308
rect 23474 13268 23480 13280
rect 23532 13268 23538 13320
rect 24949 13311 25007 13317
rect 24949 13277 24961 13311
rect 24995 13277 25007 13311
rect 24949 13271 25007 13277
rect 22281 13243 22339 13249
rect 22281 13240 22293 13243
rect 19812 13212 22293 13240
rect 1673 13175 1731 13181
rect 1673 13141 1685 13175
rect 1719 13172 1731 13175
rect 1854 13172 1860 13184
rect 1719 13144 1860 13172
rect 1719 13141 1731 13144
rect 1673 13135 1731 13141
rect 1854 13132 1860 13144
rect 1912 13132 1918 13184
rect 2958 13172 2964 13184
rect 2919 13144 2964 13172
rect 2958 13132 2964 13144
rect 3016 13132 3022 13184
rect 7006 13132 7012 13184
rect 7064 13172 7070 13184
rect 7929 13175 7987 13181
rect 7929 13172 7941 13175
rect 7064 13144 7941 13172
rect 7064 13132 7070 13144
rect 7929 13141 7941 13144
rect 7975 13141 7987 13175
rect 7929 13135 7987 13141
rect 11146 13132 11152 13184
rect 11204 13172 11210 13184
rect 11977 13175 12035 13181
rect 11977 13172 11989 13175
rect 11204 13144 11989 13172
rect 11204 13132 11210 13144
rect 11977 13141 11989 13144
rect 12023 13141 12035 13175
rect 11977 13135 12035 13141
rect 14642 13132 14648 13184
rect 14700 13132 14706 13184
rect 16942 13132 16948 13184
rect 17000 13172 17006 13184
rect 18248 13181 18276 13212
rect 22281 13209 22293 13212
rect 22327 13209 22339 13243
rect 24964 13240 24992 13271
rect 26418 13240 26424 13252
rect 24964 13212 26424 13240
rect 22281 13203 22339 13209
rect 26418 13200 26424 13212
rect 26476 13200 26482 13252
rect 27798 13240 27804 13252
rect 27738 13212 27804 13240
rect 27798 13200 27804 13212
rect 27856 13200 27862 13252
rect 17129 13175 17187 13181
rect 17129 13172 17141 13175
rect 17000 13144 17141 13172
rect 17000 13132 17006 13144
rect 17129 13141 17141 13144
rect 17175 13141 17187 13175
rect 17129 13135 17187 13141
rect 18233 13175 18291 13181
rect 18233 13141 18245 13175
rect 18279 13141 18291 13175
rect 18233 13135 18291 13141
rect 19426 13132 19432 13184
rect 19484 13172 19490 13184
rect 19521 13175 19579 13181
rect 19521 13172 19533 13175
rect 19484 13144 19533 13172
rect 19484 13132 19490 13144
rect 19521 13141 19533 13144
rect 19567 13172 19579 13175
rect 19978 13172 19984 13184
rect 19567 13144 19984 13172
rect 19567 13141 19579 13144
rect 19521 13135 19579 13141
rect 19978 13132 19984 13144
rect 20036 13132 20042 13184
rect 22370 13172 22376 13184
rect 22331 13144 22376 13172
rect 22370 13132 22376 13144
rect 22428 13132 22434 13184
rect 1104 13082 29048 13104
rect 1104 13030 7896 13082
rect 7948 13030 7960 13082
rect 8012 13030 8024 13082
rect 8076 13030 8088 13082
rect 8140 13030 8152 13082
rect 8204 13030 14842 13082
rect 14894 13030 14906 13082
rect 14958 13030 14970 13082
rect 15022 13030 15034 13082
rect 15086 13030 15098 13082
rect 15150 13030 21788 13082
rect 21840 13030 21852 13082
rect 21904 13030 21916 13082
rect 21968 13030 21980 13082
rect 22032 13030 22044 13082
rect 22096 13030 28734 13082
rect 28786 13030 28798 13082
rect 28850 13030 28862 13082
rect 28914 13030 28926 13082
rect 28978 13030 28990 13082
rect 29042 13030 29048 13082
rect 1104 13008 29048 13030
rect 6549 12971 6607 12977
rect 6549 12937 6561 12971
rect 6595 12968 6607 12971
rect 6638 12968 6644 12980
rect 6595 12940 6644 12968
rect 6595 12937 6607 12940
rect 6549 12931 6607 12937
rect 6638 12928 6644 12940
rect 6696 12928 6702 12980
rect 7006 12968 7012 12980
rect 6967 12940 7012 12968
rect 7006 12928 7012 12940
rect 7064 12928 7070 12980
rect 13446 12968 13452 12980
rect 12406 12940 13452 12968
rect 1854 12900 1860 12912
rect 1815 12872 1860 12900
rect 1854 12860 1860 12872
rect 1912 12860 1918 12912
rect 3602 12900 3608 12912
rect 3563 12872 3608 12900
rect 3602 12860 3608 12872
rect 3660 12860 3666 12912
rect 6086 12860 6092 12912
rect 6144 12900 6150 12912
rect 7024 12900 7052 12928
rect 10778 12900 10784 12912
rect 6144 12872 7052 12900
rect 9508 12872 10784 12900
rect 6144 12860 6150 12872
rect 1578 12832 1584 12844
rect 1539 12804 1584 12832
rect 1578 12792 1584 12804
rect 1636 12792 1642 12844
rect 2958 12792 2964 12844
rect 3016 12792 3022 12844
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 4798 12832 4804 12844
rect 4663 12804 4804 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 4798 12792 4804 12804
rect 4856 12792 4862 12844
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12832 5319 12835
rect 5718 12832 5724 12844
rect 5307 12804 5724 12832
rect 5307 12801 5319 12804
rect 5261 12795 5319 12801
rect 5718 12792 5724 12804
rect 5776 12832 5782 12844
rect 6546 12832 6552 12844
rect 5776 12804 6552 12832
rect 5776 12792 5782 12804
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 6917 12835 6975 12841
rect 6917 12801 6929 12835
rect 6963 12832 6975 12835
rect 9508 12832 9536 12872
rect 10778 12860 10784 12872
rect 10836 12860 10842 12912
rect 6963 12804 9536 12832
rect 9605 12835 9663 12841
rect 6963 12801 6975 12804
rect 6917 12795 6975 12801
rect 9605 12801 9617 12835
rect 9651 12832 9663 12835
rect 9766 12832 9772 12844
rect 9651 12804 9772 12832
rect 9651 12801 9663 12804
rect 9605 12795 9663 12801
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12832 10931 12835
rect 12406 12832 12434 12940
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 16850 12968 16856 12980
rect 16811 12940 16856 12968
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 16942 12928 16948 12980
rect 17000 12968 17006 12980
rect 17313 12971 17371 12977
rect 17313 12968 17325 12971
rect 17000 12940 17325 12968
rect 17000 12928 17006 12940
rect 17313 12937 17325 12940
rect 17359 12937 17371 12971
rect 20990 12968 20996 12980
rect 20951 12940 20996 12968
rect 17313 12931 17371 12937
rect 20990 12928 20996 12940
rect 21048 12928 21054 12980
rect 24578 12968 24584 12980
rect 21192 12940 24584 12968
rect 14734 12900 14740 12912
rect 14695 12872 14740 12900
rect 14734 12860 14740 12872
rect 14792 12860 14798 12912
rect 15378 12900 15384 12912
rect 15339 12872 15384 12900
rect 15378 12860 15384 12872
rect 15436 12860 15442 12912
rect 15749 12903 15807 12909
rect 15749 12869 15761 12903
rect 15795 12900 15807 12903
rect 17678 12900 17684 12912
rect 15795 12872 17684 12900
rect 15795 12869 15807 12872
rect 15749 12863 15807 12869
rect 17678 12860 17684 12872
rect 17736 12860 17742 12912
rect 21082 12900 21088 12912
rect 18892 12872 21088 12900
rect 10919 12804 12434 12832
rect 12529 12835 12587 12841
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 12529 12801 12541 12835
rect 12575 12832 12587 12835
rect 15565 12835 15623 12841
rect 12575 12804 15516 12832
rect 12575 12801 12587 12804
rect 12529 12795 12587 12801
rect 7190 12764 7196 12776
rect 7151 12736 7196 12764
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 9861 12767 9919 12773
rect 9861 12733 9873 12767
rect 9907 12733 9919 12767
rect 9861 12727 9919 12733
rect 12345 12767 12403 12773
rect 12345 12733 12357 12767
rect 12391 12764 12403 12767
rect 13354 12764 13360 12776
rect 12391 12736 13360 12764
rect 12391 12733 12403 12736
rect 12345 12727 12403 12733
rect 9876 12696 9904 12727
rect 13354 12724 13360 12736
rect 13412 12724 13418 12776
rect 9950 12696 9956 12708
rect 9876 12668 9956 12696
rect 9950 12656 9956 12668
rect 10008 12696 10014 12708
rect 10870 12696 10876 12708
rect 10008 12668 10876 12696
rect 10008 12656 10014 12668
rect 10870 12656 10876 12668
rect 10928 12656 10934 12708
rect 15488 12696 15516 12804
rect 15565 12801 15577 12835
rect 15611 12832 15623 12835
rect 15654 12832 15660 12844
rect 15611 12804 15660 12832
rect 15611 12801 15623 12804
rect 15565 12795 15623 12801
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 16666 12792 16672 12844
rect 16724 12832 16730 12844
rect 17218 12832 17224 12844
rect 16724 12804 17224 12832
rect 16724 12792 16730 12804
rect 17218 12792 17224 12804
rect 17276 12792 17282 12844
rect 18892 12841 18920 12872
rect 21082 12860 21088 12872
rect 21140 12860 21146 12912
rect 18877 12835 18935 12841
rect 18877 12832 18889 12835
rect 17328 12804 18889 12832
rect 17328 12696 17356 12804
rect 18877 12801 18889 12804
rect 18923 12801 18935 12835
rect 18877 12795 18935 12801
rect 19144 12835 19202 12841
rect 19144 12801 19156 12835
rect 19190 12832 19202 12835
rect 19426 12832 19432 12844
rect 19190 12804 19432 12832
rect 19190 12801 19202 12804
rect 19144 12795 19202 12801
rect 19426 12792 19432 12804
rect 19484 12792 19490 12844
rect 21192 12841 21220 12940
rect 24578 12928 24584 12940
rect 24636 12928 24642 12980
rect 21453 12903 21511 12909
rect 21453 12869 21465 12903
rect 21499 12900 21511 12903
rect 22462 12900 22468 12912
rect 21499 12872 22468 12900
rect 21499 12869 21511 12872
rect 21453 12863 21511 12869
rect 22462 12860 22468 12872
rect 22520 12860 22526 12912
rect 28166 12900 28172 12912
rect 28127 12872 28172 12900
rect 28166 12860 28172 12872
rect 28224 12860 28230 12912
rect 21177 12835 21235 12841
rect 21177 12801 21189 12835
rect 21223 12801 21235 12835
rect 21177 12795 21235 12801
rect 22281 12835 22339 12841
rect 22281 12801 22293 12835
rect 22327 12832 22339 12835
rect 22370 12832 22376 12844
rect 22327 12804 22376 12832
rect 22327 12801 22339 12804
rect 22281 12795 22339 12801
rect 22370 12792 22376 12804
rect 22428 12792 22434 12844
rect 22554 12841 22560 12844
rect 22548 12795 22560 12841
rect 22612 12832 22618 12844
rect 26326 12832 26332 12844
rect 22612 12804 22648 12832
rect 26287 12804 26332 12832
rect 22554 12792 22560 12795
rect 22612 12792 22618 12804
rect 26326 12792 26332 12804
rect 26384 12792 26390 12844
rect 26418 12792 26424 12844
rect 26476 12832 26482 12844
rect 27341 12835 27399 12841
rect 27341 12832 27353 12835
rect 26476 12804 27353 12832
rect 26476 12792 26482 12804
rect 27341 12801 27353 12804
rect 27387 12832 27399 12835
rect 27430 12832 27436 12844
rect 27387 12804 27436 12832
rect 27387 12801 27399 12804
rect 27341 12795 27399 12801
rect 27430 12792 27436 12804
rect 27488 12792 27494 12844
rect 27614 12792 27620 12844
rect 27672 12832 27678 12844
rect 27893 12835 27951 12841
rect 27893 12832 27905 12835
rect 27672 12804 27905 12832
rect 27672 12792 27678 12804
rect 27893 12801 27905 12804
rect 27939 12801 27951 12835
rect 27893 12795 27951 12801
rect 17494 12764 17500 12776
rect 17455 12736 17500 12764
rect 17494 12724 17500 12736
rect 17552 12724 17558 12776
rect 21266 12764 21272 12776
rect 21227 12736 21272 12764
rect 21266 12724 21272 12736
rect 21324 12724 21330 12776
rect 15488 12668 17356 12696
rect 5169 12631 5227 12637
rect 5169 12597 5181 12631
rect 5215 12628 5227 12631
rect 5442 12628 5448 12640
rect 5215 12600 5448 12628
rect 5215 12597 5227 12600
rect 5169 12591 5227 12597
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 8478 12628 8484 12640
rect 8439 12600 8484 12628
rect 8478 12588 8484 12600
rect 8536 12588 8542 12640
rect 10686 12588 10692 12640
rect 10744 12628 10750 12640
rect 10781 12631 10839 12637
rect 10781 12628 10793 12631
rect 10744 12600 10793 12628
rect 10744 12588 10750 12600
rect 10781 12597 10793 12600
rect 10827 12597 10839 12631
rect 17512 12628 17540 12724
rect 19794 12628 19800 12640
rect 17512 12600 19800 12628
rect 10781 12591 10839 12597
rect 19794 12588 19800 12600
rect 19852 12588 19858 12640
rect 19886 12588 19892 12640
rect 19944 12628 19950 12640
rect 20257 12631 20315 12637
rect 20257 12628 20269 12631
rect 19944 12600 20269 12628
rect 19944 12588 19950 12600
rect 20257 12597 20269 12600
rect 20303 12597 20315 12631
rect 20257 12591 20315 12597
rect 20898 12588 20904 12640
rect 20956 12628 20962 12640
rect 21177 12631 21235 12637
rect 21177 12628 21189 12631
rect 20956 12600 21189 12628
rect 20956 12588 20962 12600
rect 21177 12597 21189 12600
rect 21223 12597 21235 12631
rect 23658 12628 23664 12640
rect 23619 12600 23664 12628
rect 21177 12591 21235 12597
rect 23658 12588 23664 12600
rect 23716 12588 23722 12640
rect 26418 12628 26424 12640
rect 26379 12600 26424 12628
rect 26418 12588 26424 12600
rect 26476 12588 26482 12640
rect 26694 12588 26700 12640
rect 26752 12628 26758 12640
rect 27249 12631 27307 12637
rect 27249 12628 27261 12631
rect 26752 12600 27261 12628
rect 26752 12588 26758 12600
rect 27249 12597 27261 12600
rect 27295 12597 27307 12631
rect 27249 12591 27307 12597
rect 1104 12538 28888 12560
rect 1104 12486 4423 12538
rect 4475 12486 4487 12538
rect 4539 12486 4551 12538
rect 4603 12486 4615 12538
rect 4667 12486 4679 12538
rect 4731 12486 11369 12538
rect 11421 12486 11433 12538
rect 11485 12486 11497 12538
rect 11549 12486 11561 12538
rect 11613 12486 11625 12538
rect 11677 12486 18315 12538
rect 18367 12486 18379 12538
rect 18431 12486 18443 12538
rect 18495 12486 18507 12538
rect 18559 12486 18571 12538
rect 18623 12486 25261 12538
rect 25313 12486 25325 12538
rect 25377 12486 25389 12538
rect 25441 12486 25453 12538
rect 25505 12486 25517 12538
rect 25569 12486 28888 12538
rect 1104 12464 28888 12486
rect 9766 12384 9772 12436
rect 9824 12424 9830 12436
rect 9861 12427 9919 12433
rect 9861 12424 9873 12427
rect 9824 12396 9873 12424
rect 9824 12384 9830 12396
rect 9861 12393 9873 12396
rect 9907 12393 9919 12427
rect 9861 12387 9919 12393
rect 14182 12384 14188 12436
rect 14240 12424 14246 12436
rect 14277 12427 14335 12433
rect 14277 12424 14289 12427
rect 14240 12396 14289 12424
rect 14240 12384 14246 12396
rect 14277 12393 14289 12396
rect 14323 12393 14335 12427
rect 14277 12387 14335 12393
rect 15565 12427 15623 12433
rect 15565 12393 15577 12427
rect 15611 12424 15623 12427
rect 17034 12424 17040 12436
rect 15611 12396 17040 12424
rect 15611 12393 15623 12396
rect 15565 12387 15623 12393
rect 17034 12384 17040 12396
rect 17092 12384 17098 12436
rect 17221 12427 17279 12433
rect 17221 12393 17233 12427
rect 17267 12424 17279 12427
rect 17586 12424 17592 12436
rect 17267 12396 17592 12424
rect 17267 12393 17279 12396
rect 17221 12387 17279 12393
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 19426 12424 19432 12436
rect 19387 12396 19432 12424
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 21177 12427 21235 12433
rect 21177 12393 21189 12427
rect 21223 12424 21235 12427
rect 21266 12424 21272 12436
rect 21223 12396 21272 12424
rect 21223 12393 21235 12396
rect 21177 12387 21235 12393
rect 21266 12384 21272 12396
rect 21324 12384 21330 12436
rect 22554 12384 22560 12436
rect 22612 12424 22618 12436
rect 22649 12427 22707 12433
rect 22649 12424 22661 12427
rect 22612 12396 22661 12424
rect 22612 12384 22618 12396
rect 22649 12393 22661 12396
rect 22695 12393 22707 12427
rect 22649 12387 22707 12393
rect 27430 12384 27436 12436
rect 27488 12424 27494 12436
rect 28169 12427 28227 12433
rect 28169 12424 28181 12427
rect 27488 12396 28181 12424
rect 27488 12384 27494 12396
rect 28169 12393 28181 12396
rect 28215 12393 28227 12427
rect 28169 12387 28227 12393
rect 10778 12316 10784 12368
rect 10836 12356 10842 12368
rect 10836 12328 14044 12356
rect 10836 12316 10842 12328
rect 5718 12288 5724 12300
rect 5679 12260 5724 12288
rect 5718 12248 5724 12260
rect 5776 12248 5782 12300
rect 9306 12288 9312 12300
rect 9267 12260 9312 12288
rect 9306 12248 9312 12260
rect 9364 12248 9370 12300
rect 10962 12288 10968 12300
rect 10875 12260 10968 12288
rect 10962 12248 10968 12260
rect 11020 12288 11026 12300
rect 13906 12288 13912 12300
rect 11020 12260 13912 12288
rect 11020 12248 11026 12260
rect 13906 12248 13912 12260
rect 13964 12248 13970 12300
rect 14016 12232 14044 12328
rect 19794 12316 19800 12368
rect 19852 12356 19858 12368
rect 19852 12328 22094 12356
rect 19852 12316 19858 12328
rect 14826 12288 14832 12300
rect 14787 12260 14832 12288
rect 14826 12248 14832 12260
rect 14884 12248 14890 12300
rect 16942 12288 16948 12300
rect 16903 12260 16948 12288
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 19886 12288 19892 12300
rect 19847 12260 19892 12288
rect 19886 12248 19892 12260
rect 19944 12248 19950 12300
rect 19996 12297 20024 12328
rect 19981 12291 20039 12297
rect 19981 12257 19993 12291
rect 20027 12257 20039 12291
rect 19981 12251 20039 12257
rect 20070 12248 20076 12300
rect 20128 12288 20134 12300
rect 20717 12291 20775 12297
rect 20717 12288 20729 12291
rect 20128 12260 20729 12288
rect 20128 12248 20134 12260
rect 20717 12257 20729 12260
rect 20763 12257 20775 12291
rect 22066 12288 22094 12328
rect 23293 12291 23351 12297
rect 23293 12288 23305 12291
rect 22066 12260 23305 12288
rect 20717 12251 20775 12257
rect 23293 12257 23305 12260
rect 23339 12288 23351 12291
rect 23750 12288 23756 12300
rect 23339 12260 23756 12288
rect 23339 12257 23351 12260
rect 23293 12251 23351 12257
rect 23750 12248 23756 12260
rect 23808 12248 23814 12300
rect 26418 12288 26424 12300
rect 26379 12260 26424 12288
rect 26418 12248 26424 12260
rect 26476 12248 26482 12300
rect 26694 12288 26700 12300
rect 26655 12260 26700 12288
rect 26694 12248 26700 12260
rect 26752 12248 26758 12300
rect 4065 12223 4123 12229
rect 4065 12189 4077 12223
rect 4111 12220 4123 12223
rect 4890 12220 4896 12232
rect 4111 12192 4896 12220
rect 4111 12189 4123 12192
rect 4065 12183 4123 12189
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 8478 12180 8484 12232
rect 8536 12220 8542 12232
rect 9214 12220 9220 12232
rect 8536 12192 9220 12220
rect 8536 12180 8542 12192
rect 9214 12180 9220 12192
rect 9272 12220 9278 12232
rect 9401 12223 9459 12229
rect 9401 12220 9413 12223
rect 9272 12192 9413 12220
rect 9272 12180 9278 12192
rect 9401 12189 9413 12192
rect 9447 12189 9459 12223
rect 11238 12220 11244 12232
rect 11199 12192 11244 12220
rect 9401 12183 9459 12189
rect 11238 12180 11244 12192
rect 11296 12180 11302 12232
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 12805 12223 12863 12229
rect 12805 12189 12817 12223
rect 12851 12220 12863 12223
rect 13446 12220 13452 12232
rect 12851 12192 13452 12220
rect 12851 12189 12863 12192
rect 12805 12183 12863 12189
rect 4617 12155 4675 12161
rect 4617 12121 4629 12155
rect 4663 12152 4675 12155
rect 4798 12152 4804 12164
rect 4663 12124 4804 12152
rect 4663 12121 4675 12124
rect 4617 12115 4675 12121
rect 4798 12112 4804 12124
rect 4856 12112 4862 12164
rect 5988 12155 6046 12161
rect 5988 12121 6000 12155
rect 6034 12152 6046 12155
rect 6546 12152 6552 12164
rect 6034 12124 6552 12152
rect 6034 12121 6046 12124
rect 5988 12115 6046 12121
rect 6546 12112 6552 12124
rect 6604 12112 6610 12164
rect 10870 12112 10876 12164
rect 10928 12152 10934 12164
rect 11992 12152 12020 12183
rect 13446 12180 13452 12192
rect 13504 12180 13510 12232
rect 13998 12220 14004 12232
rect 13911 12192 14004 12220
rect 13998 12180 14004 12192
rect 14056 12220 14062 12232
rect 14645 12223 14703 12229
rect 14645 12220 14657 12223
rect 14056 12192 14657 12220
rect 14056 12180 14062 12192
rect 14645 12189 14657 12192
rect 14691 12189 14703 12223
rect 14645 12183 14703 12189
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12220 14795 12223
rect 15194 12220 15200 12232
rect 14783 12192 15200 12220
rect 14783 12189 14795 12192
rect 14737 12183 14795 12189
rect 10928 12124 12020 12152
rect 14660 12152 14688 12183
rect 15194 12180 15200 12192
rect 15252 12220 15258 12232
rect 15473 12223 15531 12229
rect 15473 12220 15485 12223
rect 15252 12192 15485 12220
rect 15252 12180 15258 12192
rect 15473 12189 15485 12192
rect 15519 12189 15531 12223
rect 15654 12220 15660 12232
rect 15615 12192 15660 12220
rect 15473 12183 15531 12189
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 16853 12223 16911 12229
rect 16853 12189 16865 12223
rect 16899 12189 16911 12223
rect 20806 12220 20812 12232
rect 20767 12192 20812 12220
rect 16853 12183 16911 12189
rect 16666 12152 16672 12164
rect 14660 12124 16672 12152
rect 10928 12112 10934 12124
rect 16666 12112 16672 12124
rect 16724 12112 16730 12164
rect 16868 12152 16896 12183
rect 20806 12180 20812 12192
rect 20864 12180 20870 12232
rect 23014 12220 23020 12232
rect 22975 12192 23020 12220
rect 23014 12180 23020 12192
rect 23072 12180 23078 12232
rect 23109 12223 23167 12229
rect 23109 12189 23121 12223
rect 23155 12220 23167 12223
rect 23658 12220 23664 12232
rect 23155 12192 23664 12220
rect 23155 12189 23167 12192
rect 23109 12183 23167 12189
rect 23658 12180 23664 12192
rect 23716 12180 23722 12232
rect 25685 12223 25743 12229
rect 25685 12220 25697 12223
rect 24826 12192 25697 12220
rect 24826 12152 24854 12192
rect 25685 12189 25697 12192
rect 25731 12220 25743 12223
rect 26326 12220 26332 12232
rect 25731 12192 26332 12220
rect 25731 12189 25743 12192
rect 25685 12183 25743 12189
rect 26326 12180 26332 12192
rect 26384 12180 26390 12232
rect 27982 12152 27988 12164
rect 16868 12124 24854 12152
rect 27922 12124 27988 12152
rect 27982 12112 27988 12124
rect 28040 12112 28046 12164
rect 7006 12044 7012 12096
rect 7064 12084 7070 12096
rect 7101 12087 7159 12093
rect 7101 12084 7113 12087
rect 7064 12056 7113 12084
rect 7064 12044 7070 12056
rect 7101 12053 7113 12056
rect 7147 12053 7159 12087
rect 9490 12084 9496 12096
rect 9403 12056 9496 12084
rect 7101 12047 7159 12053
rect 9490 12044 9496 12056
rect 9548 12084 9554 12096
rect 11882 12084 11888 12096
rect 9548 12056 11888 12084
rect 9548 12044 9554 12056
rect 11882 12044 11888 12056
rect 11940 12044 11946 12096
rect 12066 12084 12072 12096
rect 12027 12056 12072 12084
rect 12066 12044 12072 12056
rect 12124 12044 12130 12096
rect 12250 12044 12256 12096
rect 12308 12084 12314 12096
rect 12713 12087 12771 12093
rect 12713 12084 12725 12087
rect 12308 12056 12725 12084
rect 12308 12044 12314 12056
rect 12713 12053 12725 12056
rect 12759 12053 12771 12087
rect 16684 12084 16712 12112
rect 19797 12087 19855 12093
rect 19797 12084 19809 12087
rect 16684 12056 19809 12084
rect 12713 12047 12771 12053
rect 19797 12053 19809 12056
rect 19843 12053 19855 12087
rect 19797 12047 19855 12053
rect 25038 12044 25044 12096
rect 25096 12084 25102 12096
rect 25593 12087 25651 12093
rect 25593 12084 25605 12087
rect 25096 12056 25605 12084
rect 25096 12044 25102 12056
rect 25593 12053 25605 12056
rect 25639 12053 25651 12087
rect 25593 12047 25651 12053
rect 1104 11994 29048 12016
rect 1104 11942 7896 11994
rect 7948 11942 7960 11994
rect 8012 11942 8024 11994
rect 8076 11942 8088 11994
rect 8140 11942 8152 11994
rect 8204 11942 14842 11994
rect 14894 11942 14906 11994
rect 14958 11942 14970 11994
rect 15022 11942 15034 11994
rect 15086 11942 15098 11994
rect 15150 11942 21788 11994
rect 21840 11942 21852 11994
rect 21904 11942 21916 11994
rect 21968 11942 21980 11994
rect 22032 11942 22044 11994
rect 22096 11942 28734 11994
rect 28786 11942 28798 11994
rect 28850 11942 28862 11994
rect 28914 11942 28926 11994
rect 28978 11942 28990 11994
rect 29042 11942 29048 11994
rect 1104 11920 29048 11942
rect 6546 11880 6552 11892
rect 6507 11852 6552 11880
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 7006 11880 7012 11892
rect 6967 11852 7012 11880
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 11054 11880 11060 11892
rect 9692 11852 11060 11880
rect 9692 11756 9720 11852
rect 11054 11840 11060 11852
rect 11112 11840 11118 11892
rect 12066 11840 12072 11892
rect 12124 11880 12130 11892
rect 12124 11852 12434 11880
rect 12124 11840 12130 11852
rect 9858 11772 9864 11824
rect 9916 11812 9922 11824
rect 12250 11812 12256 11824
rect 9916 11784 11008 11812
rect 9916 11772 9922 11784
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11713 3111 11747
rect 3053 11707 3111 11713
rect 3237 11747 3295 11753
rect 3237 11713 3249 11747
rect 3283 11744 3295 11747
rect 4154 11744 4160 11756
rect 3283 11716 4160 11744
rect 3283 11713 3295 11716
rect 3237 11707 3295 11713
rect 2314 11676 2320 11688
rect 2275 11648 2320 11676
rect 2314 11636 2320 11648
rect 2372 11636 2378 11688
rect 3068 11676 3096 11707
rect 4154 11704 4160 11716
rect 4212 11704 4218 11756
rect 5353 11747 5411 11753
rect 5353 11713 5365 11747
rect 5399 11744 5411 11747
rect 6362 11744 6368 11756
rect 5399 11716 6368 11744
rect 5399 11713 5411 11716
rect 5353 11707 5411 11713
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11744 6975 11747
rect 9674 11744 9680 11756
rect 6963 11716 9680 11744
rect 6963 11713 6975 11716
rect 6917 11707 6975 11713
rect 9674 11704 9680 11716
rect 9732 11704 9738 11756
rect 10686 11744 10692 11756
rect 10647 11716 10692 11744
rect 10686 11704 10692 11716
rect 10744 11704 10750 11756
rect 10980 11753 11008 11784
rect 11716 11784 12256 11812
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11713 11023 11747
rect 11146 11744 11152 11756
rect 11107 11716 11152 11744
rect 10965 11707 11023 11713
rect 11146 11704 11152 11716
rect 11204 11704 11210 11756
rect 11716 11753 11744 11784
rect 12250 11772 12256 11784
rect 12308 11772 12314 11824
rect 12406 11812 12434 11852
rect 16758 11840 16764 11892
rect 16816 11880 16822 11892
rect 18233 11883 18291 11889
rect 18233 11880 18245 11883
rect 16816 11852 18245 11880
rect 16816 11840 16822 11852
rect 18233 11849 18245 11852
rect 18279 11880 18291 11883
rect 20070 11880 20076 11892
rect 18279 11852 20076 11880
rect 18279 11849 18291 11852
rect 18233 11843 18291 11849
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 26326 11840 26332 11892
rect 26384 11880 26390 11892
rect 26513 11883 26571 11889
rect 26513 11880 26525 11883
rect 26384 11852 26525 11880
rect 26384 11840 26390 11852
rect 26513 11849 26525 11852
rect 26559 11849 26571 11883
rect 26513 11843 26571 11849
rect 13722 11812 13728 11824
rect 12406 11784 12466 11812
rect 13635 11784 13728 11812
rect 13722 11772 13728 11784
rect 13780 11812 13786 11824
rect 16574 11812 16580 11824
rect 13780 11784 16580 11812
rect 13780 11772 13786 11784
rect 16574 11772 16580 11784
rect 16632 11772 16638 11824
rect 25038 11812 25044 11824
rect 24999 11784 25044 11812
rect 25038 11772 25044 11784
rect 25096 11772 25102 11824
rect 25682 11772 25688 11824
rect 25740 11772 25746 11824
rect 27982 11812 27988 11824
rect 27943 11784 27988 11812
rect 27982 11772 27988 11784
rect 28040 11772 28046 11824
rect 27344 11756 27396 11762
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 14642 11704 14648 11756
rect 14700 11744 14706 11756
rect 15013 11747 15071 11753
rect 15013 11744 15025 11747
rect 14700 11716 15025 11744
rect 14700 11704 14706 11716
rect 15013 11713 15025 11716
rect 15059 11713 15071 11747
rect 15013 11707 15071 11713
rect 16666 11704 16672 11756
rect 16724 11744 16730 11756
rect 17126 11753 17132 11756
rect 16853 11747 16911 11753
rect 16853 11744 16865 11747
rect 16724 11716 16865 11744
rect 16724 11704 16730 11716
rect 16853 11713 16865 11716
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 17120 11707 17132 11753
rect 17184 11744 17190 11756
rect 19705 11747 19763 11753
rect 17184 11716 17220 11744
rect 17126 11704 17132 11707
rect 17184 11704 17190 11716
rect 19705 11713 19717 11747
rect 19751 11713 19763 11747
rect 19705 11707 19763 11713
rect 4246 11676 4252 11688
rect 3068 11648 4252 11676
rect 4246 11636 4252 11648
rect 4304 11636 4310 11688
rect 7190 11676 7196 11688
rect 7151 11648 7196 11676
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 10778 11676 10784 11688
rect 10739 11648 10784 11676
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 10873 11679 10931 11685
rect 10873 11645 10885 11679
rect 10919 11676 10931 11679
rect 11974 11676 11980 11688
rect 10919 11648 11836 11676
rect 11935 11648 11980 11676
rect 10919 11645 10931 11648
rect 10873 11639 10931 11645
rect 11808 11552 11836 11648
rect 11974 11636 11980 11648
rect 12032 11636 12038 11688
rect 14734 11636 14740 11688
rect 14792 11676 14798 11688
rect 14921 11679 14979 11685
rect 14921 11676 14933 11679
rect 14792 11648 14933 11676
rect 14792 11636 14798 11648
rect 14921 11645 14933 11648
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 19720 11608 19748 11707
rect 20162 11704 20168 11756
rect 20220 11744 20226 11756
rect 23201 11747 23259 11753
rect 20220 11716 20562 11744
rect 20220 11704 20226 11716
rect 23201 11713 23213 11747
rect 23247 11744 23259 11747
rect 24029 11747 24087 11753
rect 24029 11744 24041 11747
rect 23247 11716 24041 11744
rect 23247 11713 23259 11716
rect 23201 11707 23259 11713
rect 24029 11713 24041 11716
rect 24075 11744 24087 11747
rect 24670 11744 24676 11756
rect 24075 11716 24676 11744
rect 24075 11713 24087 11716
rect 24029 11707 24087 11713
rect 24670 11704 24676 11716
rect 24728 11704 24734 11756
rect 27344 11698 27396 11704
rect 19797 11679 19855 11685
rect 19797 11645 19809 11679
rect 19843 11676 19855 11679
rect 19886 11676 19892 11688
rect 19843 11648 19892 11676
rect 19843 11645 19855 11648
rect 19797 11639 19855 11645
rect 19886 11636 19892 11648
rect 19944 11636 19950 11688
rect 20622 11676 20628 11688
rect 20583 11648 20628 11676
rect 20622 11636 20628 11648
rect 20680 11636 20686 11688
rect 21266 11636 21272 11688
rect 21324 11676 21330 11688
rect 21361 11679 21419 11685
rect 21361 11676 21373 11679
rect 21324 11648 21373 11676
rect 21324 11636 21330 11648
rect 21361 11645 21373 11648
rect 21407 11645 21419 11679
rect 21361 11639 21419 11645
rect 22462 11636 22468 11688
rect 22520 11676 22526 11688
rect 22833 11679 22891 11685
rect 22833 11676 22845 11679
rect 22520 11648 22845 11676
rect 22520 11636 22526 11648
rect 22833 11645 22845 11648
rect 22879 11645 22891 11679
rect 22833 11639 22891 11645
rect 23293 11679 23351 11685
rect 23293 11645 23305 11679
rect 23339 11676 23351 11679
rect 23658 11676 23664 11688
rect 23339 11648 23664 11676
rect 23339 11645 23351 11648
rect 23293 11639 23351 11645
rect 23658 11636 23664 11648
rect 23716 11636 23722 11688
rect 24762 11676 24768 11688
rect 24723 11648 24768 11676
rect 24762 11636 24768 11648
rect 24820 11636 24826 11688
rect 27433 11679 27491 11685
rect 27433 11645 27445 11679
rect 27479 11676 27491 11679
rect 27522 11676 27528 11688
rect 27479 11648 27528 11676
rect 27479 11645 27491 11648
rect 27433 11639 27491 11645
rect 27522 11636 27528 11648
rect 27580 11636 27586 11688
rect 20898 11608 20904 11620
rect 19720 11580 20904 11608
rect 20898 11568 20904 11580
rect 20956 11568 20962 11620
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 10505 11543 10563 11549
rect 10505 11540 10517 11543
rect 8536 11512 10517 11540
rect 8536 11500 8542 11512
rect 10505 11509 10517 11512
rect 10551 11509 10563 11543
rect 10505 11503 10563 11509
rect 11790 11500 11796 11552
rect 11848 11500 11854 11552
rect 15381 11543 15439 11549
rect 15381 11509 15393 11543
rect 15427 11540 15439 11543
rect 18138 11540 18144 11552
rect 15427 11512 18144 11540
rect 15427 11509 15439 11512
rect 15381 11503 15439 11509
rect 18138 11500 18144 11512
rect 18196 11500 18202 11552
rect 19334 11540 19340 11552
rect 19295 11512 19340 11540
rect 19334 11500 19340 11512
rect 19392 11500 19398 11552
rect 19518 11500 19524 11552
rect 19576 11540 19582 11552
rect 19886 11540 19892 11552
rect 19576 11512 19892 11540
rect 19576 11500 19582 11512
rect 19886 11500 19892 11512
rect 19944 11500 19950 11552
rect 23934 11540 23940 11552
rect 23895 11512 23940 11540
rect 23934 11500 23940 11512
rect 23992 11500 23998 11552
rect 1104 11450 28888 11472
rect 1104 11398 4423 11450
rect 4475 11398 4487 11450
rect 4539 11398 4551 11450
rect 4603 11398 4615 11450
rect 4667 11398 4679 11450
rect 4731 11398 11369 11450
rect 11421 11398 11433 11450
rect 11485 11398 11497 11450
rect 11549 11398 11561 11450
rect 11613 11398 11625 11450
rect 11677 11398 18315 11450
rect 18367 11398 18379 11450
rect 18431 11398 18443 11450
rect 18495 11398 18507 11450
rect 18559 11398 18571 11450
rect 18623 11398 25261 11450
rect 25313 11398 25325 11450
rect 25377 11398 25389 11450
rect 25441 11398 25453 11450
rect 25505 11398 25517 11450
rect 25569 11398 28888 11450
rect 1104 11376 28888 11398
rect 6362 11296 6368 11348
rect 6420 11336 6426 11348
rect 10781 11339 10839 11345
rect 6420 11308 7144 11336
rect 6420 11296 6426 11308
rect 2958 11228 2964 11280
rect 3016 11268 3022 11280
rect 3329 11271 3387 11277
rect 3329 11268 3341 11271
rect 3016 11240 3341 11268
rect 3016 11228 3022 11240
rect 3329 11237 3341 11240
rect 3375 11237 3387 11271
rect 3329 11231 3387 11237
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 6380 11200 6408 11296
rect 7006 11268 7012 11280
rect 6656 11240 7012 11268
rect 6656 11209 6684 11240
rect 7006 11228 7012 11240
rect 7064 11228 7070 11280
rect 7116 11268 7144 11308
rect 10781 11305 10793 11339
rect 10827 11336 10839 11339
rect 11974 11336 11980 11348
rect 10827 11308 11980 11336
rect 10827 11305 10839 11308
rect 10781 11299 10839 11305
rect 11974 11296 11980 11308
rect 12032 11296 12038 11348
rect 17126 11336 17132 11348
rect 17087 11308 17132 11336
rect 17126 11296 17132 11308
rect 17184 11296 17190 11348
rect 19610 11336 19616 11348
rect 19571 11308 19616 11336
rect 19610 11296 19616 11308
rect 19668 11296 19674 11348
rect 19886 11336 19892 11348
rect 19847 11308 19892 11336
rect 19886 11296 19892 11308
rect 19944 11296 19950 11348
rect 24762 11336 24768 11348
rect 24723 11308 24768 11336
rect 24762 11296 24768 11308
rect 24820 11296 24826 11348
rect 14182 11268 14188 11280
rect 7116 11240 14188 11268
rect 14182 11228 14188 11240
rect 14240 11228 14246 11280
rect 19702 11228 19708 11280
rect 19760 11268 19766 11280
rect 22373 11271 22431 11277
rect 22373 11268 22385 11271
rect 19760 11240 22385 11268
rect 19760 11228 19766 11240
rect 22373 11237 22385 11240
rect 22419 11237 22431 11271
rect 22373 11231 22431 11237
rect 5123 11172 6408 11200
rect 6641 11203 6699 11209
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 6641 11169 6653 11203
rect 6687 11169 6699 11203
rect 6641 11163 6699 11169
rect 6917 11203 6975 11209
rect 6917 11169 6929 11203
rect 6963 11200 6975 11203
rect 9030 11200 9036 11212
rect 6963 11172 9036 11200
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 9030 11160 9036 11172
rect 9088 11160 9094 11212
rect 9214 11200 9220 11212
rect 9175 11172 9220 11200
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11200 9735 11203
rect 10226 11200 10232 11212
rect 9723 11172 10232 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 10226 11160 10232 11172
rect 10284 11160 10290 11212
rect 11054 11160 11060 11212
rect 11112 11200 11118 11212
rect 14734 11200 14740 11212
rect 11112 11172 13860 11200
rect 14695 11172 14740 11200
rect 11112 11160 11118 11172
rect 1578 11132 1584 11144
rect 1539 11104 1584 11132
rect 1578 11092 1584 11104
rect 1636 11092 1642 11144
rect 5442 11132 5448 11144
rect 5403 11104 5448 11132
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 5626 11092 5632 11144
rect 5684 11132 5690 11144
rect 6549 11135 6607 11141
rect 6549 11132 6561 11135
rect 5684 11104 6561 11132
rect 5684 11092 5690 11104
rect 6549 11101 6561 11104
rect 6595 11132 6607 11135
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 6595 11104 7389 11132
rect 6595 11101 6607 11104
rect 6549 11095 6607 11101
rect 7377 11101 7389 11104
rect 7423 11101 7435 11135
rect 7377 11095 7435 11101
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11132 8355 11135
rect 9122 11132 9128 11144
rect 8343 11104 9128 11132
rect 8343 11101 8355 11104
rect 8297 11095 8355 11101
rect 9122 11092 9128 11104
rect 9180 11132 9186 11144
rect 9309 11135 9367 11141
rect 9309 11132 9321 11135
rect 9180 11104 9321 11132
rect 9180 11092 9186 11104
rect 9309 11101 9321 11104
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 10873 11135 10931 11141
rect 10873 11101 10885 11135
rect 10919 11132 10931 11135
rect 11238 11132 11244 11144
rect 10919 11104 11244 11132
rect 10919 11101 10931 11104
rect 10873 11095 10931 11101
rect 11238 11092 11244 11104
rect 11296 11132 11302 11144
rect 11793 11135 11851 11141
rect 11296 11104 11560 11132
rect 11296 11092 11302 11104
rect 1854 11064 1860 11076
rect 1815 11036 1860 11064
rect 1854 11024 1860 11036
rect 1912 11024 1918 11076
rect 2314 11024 2320 11076
rect 2372 11024 2378 11076
rect 11532 11073 11560 11104
rect 11793 11101 11805 11135
rect 11839 11132 11851 11135
rect 13722 11132 13728 11144
rect 11839 11104 13728 11132
rect 11839 11101 11851 11104
rect 11793 11095 11851 11101
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 13832 11132 13860 11172
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 14826 11160 14832 11212
rect 14884 11200 14890 11212
rect 14921 11203 14979 11209
rect 14921 11200 14933 11203
rect 14884 11172 14933 11200
rect 14884 11160 14890 11172
rect 14921 11169 14933 11172
rect 14967 11200 14979 11203
rect 16577 11203 16635 11209
rect 16577 11200 16589 11203
rect 14967 11172 16589 11200
rect 14967 11169 14979 11172
rect 14921 11163 14979 11169
rect 16577 11169 16589 11172
rect 16623 11200 16635 11203
rect 17402 11200 17408 11212
rect 16623 11172 17408 11200
rect 16623 11169 16635 11172
rect 16577 11163 16635 11169
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 19334 11160 19340 11212
rect 19392 11200 19398 11212
rect 19521 11203 19579 11209
rect 19521 11200 19533 11203
rect 19392 11172 19533 11200
rect 19392 11160 19398 11172
rect 19521 11169 19533 11172
rect 19567 11169 19579 11203
rect 20898 11200 20904 11212
rect 19521 11163 19579 11169
rect 20640 11172 20904 11200
rect 14645 11135 14703 11141
rect 14645 11132 14657 11135
rect 13832 11104 14657 11132
rect 14645 11101 14657 11104
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11132 16727 11135
rect 16758 11132 16764 11144
rect 16715 11104 16764 11132
rect 16715 11101 16727 11104
rect 16669 11095 16727 11101
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 18138 11092 18144 11144
rect 18196 11132 18202 11144
rect 20640 11141 20668 11172
rect 20898 11160 20904 11172
rect 20956 11200 20962 11212
rect 25682 11200 25688 11212
rect 20956 11172 22094 11200
rect 25643 11172 25688 11200
rect 20956 11160 20962 11172
rect 19705 11135 19763 11141
rect 19705 11132 19717 11135
rect 18196 11104 19717 11132
rect 18196 11092 18202 11104
rect 19705 11101 19717 11104
rect 19751 11101 19763 11135
rect 19705 11095 19763 11101
rect 20625 11135 20683 11141
rect 20625 11101 20637 11135
rect 20671 11101 20683 11135
rect 20625 11095 20683 11101
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 21085 11135 21143 11141
rect 21085 11132 21097 11135
rect 20772 11104 21097 11132
rect 20772 11092 20778 11104
rect 21085 11101 21097 11104
rect 21131 11101 21143 11135
rect 22066 11132 22094 11172
rect 25682 11160 25688 11172
rect 25740 11160 25746 11212
rect 26050 11160 26056 11212
rect 26108 11200 26114 11212
rect 27338 11200 27344 11212
rect 26108 11172 27344 11200
rect 26108 11160 26114 11172
rect 23293 11135 23351 11141
rect 23293 11132 23305 11135
rect 22066 11104 23305 11132
rect 21085 11095 21143 11101
rect 23293 11101 23305 11104
rect 23339 11101 23351 11135
rect 24670 11132 24676 11144
rect 24631 11104 24676 11132
rect 23293 11095 23351 11101
rect 24670 11092 24676 11104
rect 24728 11092 24734 11144
rect 26528 11118 26556 11172
rect 27338 11160 27344 11172
rect 27396 11160 27402 11212
rect 26602 11092 26608 11144
rect 26660 11132 26666 11144
rect 27522 11132 27528 11144
rect 26660 11104 27528 11132
rect 26660 11092 26666 11104
rect 27522 11092 27528 11104
rect 27580 11092 27586 11144
rect 11517 11067 11575 11073
rect 11517 11033 11529 11067
rect 11563 11064 11575 11067
rect 13078 11064 13084 11076
rect 11563 11036 13084 11064
rect 11563 11033 11575 11036
rect 11517 11027 11575 11033
rect 13078 11024 13084 11036
rect 13136 11024 13142 11076
rect 19426 11064 19432 11076
rect 13832 11036 19288 11064
rect 19387 11036 19432 11064
rect 7098 10956 7104 11008
rect 7156 10996 7162 11008
rect 7469 10999 7527 11005
rect 7469 10996 7481 10999
rect 7156 10968 7481 10996
rect 7156 10956 7162 10968
rect 7469 10965 7481 10968
rect 7515 10965 7527 10999
rect 7469 10959 7527 10965
rect 7650 10956 7656 11008
rect 7708 10996 7714 11008
rect 8205 10999 8263 11005
rect 8205 10996 8217 10999
rect 7708 10968 8217 10996
rect 7708 10956 7714 10968
rect 8205 10965 8217 10968
rect 8251 10965 8263 10999
rect 8205 10959 8263 10965
rect 12158 10956 12164 11008
rect 12216 10996 12222 11008
rect 13832 10996 13860 11036
rect 14274 10996 14280 11008
rect 12216 10968 13860 10996
rect 14235 10968 14280 10996
rect 12216 10956 12222 10968
rect 14274 10956 14280 10968
rect 14332 10956 14338 11008
rect 16776 11005 16804 11036
rect 16761 10999 16819 11005
rect 16761 10965 16773 10999
rect 16807 10996 16819 10999
rect 19260 10996 19288 11036
rect 19426 11024 19432 11036
rect 19484 11024 19490 11076
rect 23474 11064 23480 11076
rect 19536 11036 23480 11064
rect 19536 10996 19564 11036
rect 23474 11024 23480 11036
rect 23532 11064 23538 11076
rect 23658 11064 23664 11076
rect 23532 11036 23664 11064
rect 23532 11024 23538 11036
rect 23658 11024 23664 11036
rect 23716 11024 23722 11076
rect 20530 10996 20536 11008
rect 16807 10968 16841 10996
rect 19260 10968 19564 10996
rect 20491 10968 20536 10996
rect 16807 10965 16819 10968
rect 16761 10959 16819 10965
rect 20530 10956 20536 10968
rect 20588 10956 20594 11008
rect 22830 10956 22836 11008
rect 22888 10996 22894 11008
rect 23385 10999 23443 11005
rect 23385 10996 23397 10999
rect 22888 10968 23397 10996
rect 22888 10956 22894 10968
rect 23385 10965 23397 10968
rect 23431 10965 23443 10999
rect 23385 10959 23443 10965
rect 1104 10906 29048 10928
rect 1104 10854 7896 10906
rect 7948 10854 7960 10906
rect 8012 10854 8024 10906
rect 8076 10854 8088 10906
rect 8140 10854 8152 10906
rect 8204 10854 14842 10906
rect 14894 10854 14906 10906
rect 14958 10854 14970 10906
rect 15022 10854 15034 10906
rect 15086 10854 15098 10906
rect 15150 10854 21788 10906
rect 21840 10854 21852 10906
rect 21904 10854 21916 10906
rect 21968 10854 21980 10906
rect 22032 10854 22044 10906
rect 22096 10854 28734 10906
rect 28786 10854 28798 10906
rect 28850 10854 28862 10906
rect 28914 10854 28926 10906
rect 28978 10854 28990 10906
rect 29042 10854 29048 10906
rect 1104 10832 29048 10854
rect 1854 10752 1860 10804
rect 1912 10792 1918 10804
rect 2409 10795 2467 10801
rect 2409 10792 2421 10795
rect 1912 10764 2421 10792
rect 1912 10752 1918 10764
rect 2409 10761 2421 10764
rect 2455 10761 2467 10795
rect 2409 10755 2467 10761
rect 14645 10795 14703 10801
rect 14645 10761 14657 10795
rect 14691 10792 14703 10795
rect 14734 10792 14740 10804
rect 14691 10764 14740 10792
rect 14691 10761 14703 10764
rect 14645 10755 14703 10761
rect 14734 10752 14740 10764
rect 14792 10752 14798 10804
rect 23934 10792 23940 10804
rect 23124 10764 23940 10792
rect 7377 10727 7435 10733
rect 7377 10693 7389 10727
rect 7423 10724 7435 10727
rect 7650 10724 7656 10736
rect 7423 10696 7656 10724
rect 7423 10693 7435 10696
rect 7377 10687 7435 10693
rect 7650 10684 7656 10696
rect 7708 10684 7714 10736
rect 8110 10684 8116 10736
rect 8168 10684 8174 10736
rect 9122 10724 9128 10736
rect 9083 10696 9128 10724
rect 9122 10684 9128 10696
rect 9180 10684 9186 10736
rect 13532 10727 13590 10733
rect 13532 10693 13544 10727
rect 13578 10724 13590 10727
rect 14274 10724 14280 10736
rect 13578 10696 14280 10724
rect 13578 10693 13590 10696
rect 13532 10687 13590 10693
rect 14274 10684 14280 10696
rect 14332 10684 14338 10736
rect 19702 10724 19708 10736
rect 19663 10696 19708 10724
rect 19702 10684 19708 10696
rect 19760 10684 19766 10736
rect 23124 10733 23152 10764
rect 23934 10752 23940 10764
rect 23992 10752 23998 10804
rect 24581 10795 24639 10801
rect 24581 10761 24593 10795
rect 24627 10792 24639 10795
rect 24670 10792 24676 10804
rect 24627 10764 24676 10792
rect 24627 10761 24639 10764
rect 24581 10755 24639 10761
rect 24670 10752 24676 10764
rect 24728 10752 24734 10804
rect 23109 10727 23167 10733
rect 23109 10693 23121 10727
rect 23155 10693 23167 10727
rect 23109 10687 23167 10693
rect 24118 10684 24124 10736
rect 24176 10684 24182 10736
rect 2501 10659 2559 10665
rect 2501 10625 2513 10659
rect 2547 10656 2559 10659
rect 2958 10656 2964 10668
rect 2547 10628 2964 10656
rect 2547 10625 2559 10628
rect 2501 10619 2559 10625
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 4982 10616 4988 10668
rect 5040 10616 5046 10668
rect 7098 10656 7104 10668
rect 7059 10628 7104 10656
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 13265 10659 13323 10665
rect 13265 10625 13277 10659
rect 13311 10656 13323 10659
rect 14550 10656 14556 10668
rect 13311 10628 14556 10656
rect 13311 10625 13323 10628
rect 13265 10619 13323 10625
rect 14550 10616 14556 10628
rect 14608 10616 14614 10668
rect 17218 10656 17224 10668
rect 17131 10628 17224 10656
rect 17218 10616 17224 10628
rect 17276 10656 17282 10668
rect 19245 10659 19303 10665
rect 17276 10628 18644 10656
rect 17276 10616 17282 10628
rect 3053 10591 3111 10597
rect 3053 10557 3065 10591
rect 3099 10588 3111 10591
rect 3605 10591 3663 10597
rect 3605 10588 3617 10591
rect 3099 10560 3617 10588
rect 3099 10557 3111 10560
rect 3053 10551 3111 10557
rect 3605 10557 3617 10560
rect 3651 10557 3663 10591
rect 3605 10551 3663 10557
rect 3881 10591 3939 10597
rect 3881 10557 3893 10591
rect 3927 10588 3939 10591
rect 4338 10588 4344 10600
rect 3927 10560 4344 10588
rect 3927 10557 3939 10560
rect 3881 10551 3939 10557
rect 4338 10548 4344 10560
rect 4396 10548 4402 10600
rect 17313 10591 17371 10597
rect 17313 10557 17325 10591
rect 17359 10557 17371 10591
rect 17313 10551 17371 10557
rect 17328 10520 17356 10551
rect 17402 10548 17408 10600
rect 17460 10588 17466 10600
rect 18616 10588 18644 10628
rect 19245 10625 19257 10659
rect 19291 10656 19303 10659
rect 20806 10656 20812 10668
rect 19291 10628 20812 10656
rect 19291 10625 19303 10628
rect 19245 10619 19303 10625
rect 20806 10616 20812 10628
rect 20864 10616 20870 10668
rect 22830 10656 22836 10668
rect 22791 10628 22836 10656
rect 22830 10616 22836 10628
rect 22888 10616 22894 10668
rect 27890 10656 27896 10668
rect 27851 10628 27896 10656
rect 27890 10616 27896 10628
rect 27948 10616 27954 10668
rect 21450 10588 21456 10600
rect 17460 10560 17505 10588
rect 18616 10560 20392 10588
rect 21363 10560 21456 10588
rect 17460 10548 17466 10560
rect 17862 10520 17868 10532
rect 17328 10492 17868 10520
rect 17862 10480 17868 10492
rect 17920 10480 17926 10532
rect 5353 10455 5411 10461
rect 5353 10421 5365 10455
rect 5399 10452 5411 10455
rect 5626 10452 5632 10464
rect 5399 10424 5632 10452
rect 5399 10421 5411 10424
rect 5353 10415 5411 10421
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 16758 10412 16764 10464
rect 16816 10452 16822 10464
rect 16853 10455 16911 10461
rect 16853 10452 16865 10455
rect 16816 10424 16865 10452
rect 16816 10412 16822 10424
rect 16853 10421 16865 10424
rect 16899 10421 16911 10455
rect 16853 10415 16911 10421
rect 19153 10455 19211 10461
rect 19153 10421 19165 10455
rect 19199 10452 19211 10455
rect 20254 10452 20260 10464
rect 19199 10424 20260 10452
rect 19199 10421 19211 10424
rect 19153 10415 19211 10421
rect 20254 10412 20260 10424
rect 20312 10412 20318 10464
rect 20364 10452 20392 10560
rect 21450 10548 21456 10560
rect 21508 10588 21514 10600
rect 21818 10588 21824 10600
rect 21508 10560 21824 10588
rect 21508 10548 21514 10560
rect 21818 10548 21824 10560
rect 21876 10548 21882 10600
rect 28166 10588 28172 10600
rect 28127 10560 28172 10588
rect 28166 10548 28172 10560
rect 28224 10548 28230 10600
rect 23566 10452 23572 10464
rect 20364 10424 23572 10452
rect 23566 10412 23572 10424
rect 23624 10412 23630 10464
rect 1104 10362 28888 10384
rect 1104 10310 4423 10362
rect 4475 10310 4487 10362
rect 4539 10310 4551 10362
rect 4603 10310 4615 10362
rect 4667 10310 4679 10362
rect 4731 10310 11369 10362
rect 11421 10310 11433 10362
rect 11485 10310 11497 10362
rect 11549 10310 11561 10362
rect 11613 10310 11625 10362
rect 11677 10310 18315 10362
rect 18367 10310 18379 10362
rect 18431 10310 18443 10362
rect 18495 10310 18507 10362
rect 18559 10310 18571 10362
rect 18623 10310 25261 10362
rect 25313 10310 25325 10362
rect 25377 10310 25389 10362
rect 25441 10310 25453 10362
rect 25505 10310 25517 10362
rect 25569 10310 28888 10362
rect 1104 10288 28888 10310
rect 1578 10208 1584 10260
rect 1636 10248 1642 10260
rect 2317 10251 2375 10257
rect 2317 10248 2329 10251
rect 1636 10220 2329 10248
rect 1636 10208 1642 10220
rect 2317 10217 2329 10220
rect 2363 10217 2375 10251
rect 2317 10211 2375 10217
rect 9766 10208 9772 10260
rect 9824 10248 9830 10260
rect 9953 10251 10011 10257
rect 9953 10248 9965 10251
rect 9824 10220 9965 10248
rect 9824 10208 9830 10220
rect 9953 10217 9965 10220
rect 9999 10248 10011 10251
rect 16666 10248 16672 10260
rect 9999 10220 11468 10248
rect 9999 10217 10011 10220
rect 9953 10211 10011 10217
rect 2958 10140 2964 10192
rect 3016 10180 3022 10192
rect 6365 10183 6423 10189
rect 3016 10152 4384 10180
rect 3016 10140 3022 10152
rect 4154 10112 4160 10124
rect 4115 10084 4160 10112
rect 4154 10072 4160 10084
rect 4212 10072 4218 10124
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10044 2467 10047
rect 2774 10044 2780 10056
rect 2455 10016 2780 10044
rect 2455 10013 2467 10016
rect 2409 10007 2467 10013
rect 2774 10004 2780 10016
rect 2832 10004 2838 10056
rect 4246 10044 4252 10056
rect 4159 10016 4252 10044
rect 4246 10004 4252 10016
rect 4304 10004 4310 10056
rect 4356 10044 4384 10152
rect 6365 10149 6377 10183
rect 6411 10180 6423 10183
rect 9306 10180 9312 10192
rect 6411 10152 9312 10180
rect 6411 10149 6423 10152
rect 6365 10143 6423 10149
rect 9306 10140 9312 10152
rect 9364 10140 9370 10192
rect 4982 10112 4988 10124
rect 4943 10084 4988 10112
rect 4982 10072 4988 10084
rect 5040 10072 5046 10124
rect 6086 10112 6092 10124
rect 6047 10084 6092 10112
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 8110 10072 8116 10124
rect 8168 10112 8174 10124
rect 8205 10115 8263 10121
rect 8205 10112 8217 10115
rect 8168 10084 8217 10112
rect 8168 10072 8174 10084
rect 8205 10081 8217 10084
rect 8251 10081 8263 10115
rect 8205 10075 8263 10081
rect 5997 10047 6055 10053
rect 5997 10044 6009 10047
rect 4356 10016 6009 10044
rect 5997 10013 6009 10016
rect 6043 10013 6055 10047
rect 5997 10007 6055 10013
rect 7285 10047 7343 10053
rect 7285 10013 7297 10047
rect 7331 10013 7343 10047
rect 7285 10007 7343 10013
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10013 7527 10047
rect 11333 10047 11391 10053
rect 11333 10044 11345 10047
rect 7469 10007 7527 10013
rect 10888 10016 11345 10044
rect 4264 9908 4292 10004
rect 5534 9936 5540 9988
rect 5592 9976 5598 9988
rect 7300 9976 7328 10007
rect 5592 9948 7328 9976
rect 5592 9936 5598 9948
rect 7484 9908 7512 10007
rect 10888 9988 10916 10016
rect 11333 10013 11345 10016
rect 11379 10013 11391 10047
rect 11440 10044 11468 10220
rect 16500 10220 16672 10248
rect 12342 10112 12348 10124
rect 12255 10084 12348 10112
rect 12342 10072 12348 10084
rect 12400 10112 12406 10124
rect 12618 10112 12624 10124
rect 12400 10084 12624 10112
rect 12400 10072 12406 10084
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 11440 10016 12296 10044
rect 11333 10007 11391 10013
rect 10870 9936 10876 9988
rect 10928 9936 10934 9988
rect 12268 9985 12296 10016
rect 14550 10004 14556 10056
rect 14608 10044 14614 10056
rect 16500 10053 16528 10220
rect 16666 10208 16672 10220
rect 16724 10208 16730 10260
rect 17862 10248 17868 10260
rect 17823 10220 17868 10248
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 18877 10251 18935 10257
rect 18877 10217 18889 10251
rect 18923 10248 18935 10251
rect 19426 10248 19432 10260
rect 18923 10220 19432 10248
rect 18923 10217 18935 10220
rect 18877 10211 18935 10217
rect 19426 10208 19432 10220
rect 19484 10208 19490 10260
rect 20898 10208 20904 10260
rect 20956 10248 20962 10260
rect 22005 10251 22063 10257
rect 22005 10248 22017 10251
rect 20956 10220 22017 10248
rect 20956 10208 20962 10220
rect 22005 10217 22017 10220
rect 22051 10217 22063 10251
rect 22005 10211 22063 10217
rect 17880 10112 17908 10208
rect 26602 10180 26608 10192
rect 23032 10152 26608 10180
rect 18417 10115 18475 10121
rect 18417 10112 18429 10115
rect 17880 10084 18429 10112
rect 18417 10081 18429 10084
rect 18463 10081 18475 10115
rect 20254 10112 20260 10124
rect 20215 10084 20260 10112
rect 18417 10075 18475 10081
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 20530 10112 20536 10124
rect 20491 10084 20536 10112
rect 20530 10072 20536 10084
rect 20588 10072 20594 10124
rect 23032 10056 23060 10152
rect 26602 10140 26608 10152
rect 26660 10140 26666 10192
rect 27614 10180 27620 10192
rect 27575 10152 27620 10180
rect 27614 10140 27620 10152
rect 27672 10140 27678 10192
rect 24029 10115 24087 10121
rect 24029 10081 24041 10115
rect 24075 10112 24087 10115
rect 24118 10112 24124 10124
rect 24075 10084 24124 10112
rect 24075 10081 24087 10084
rect 24029 10075 24087 10081
rect 24118 10072 24124 10084
rect 24176 10072 24182 10124
rect 26510 10072 26516 10124
rect 26568 10112 26574 10124
rect 27157 10115 27215 10121
rect 27157 10112 27169 10115
rect 26568 10084 27169 10112
rect 26568 10072 26574 10084
rect 27157 10081 27169 10084
rect 27203 10081 27215 10115
rect 27157 10075 27215 10081
rect 16758 10053 16764 10056
rect 16485 10047 16543 10053
rect 16485 10044 16497 10047
rect 14608 10016 16497 10044
rect 14608 10004 14614 10016
rect 16485 10013 16497 10016
rect 16531 10013 16543 10047
rect 16752 10044 16764 10053
rect 16719 10016 16764 10044
rect 16485 10007 16543 10013
rect 16752 10007 16764 10016
rect 16758 10004 16764 10007
rect 16816 10004 16822 10056
rect 18506 10044 18512 10056
rect 18467 10016 18512 10044
rect 18506 10004 18512 10016
rect 18564 10004 18570 10056
rect 19797 10047 19855 10053
rect 19797 10013 19809 10047
rect 19843 10013 19855 10047
rect 23014 10044 23020 10056
rect 22975 10016 23020 10044
rect 19797 10007 19855 10013
rect 11088 9979 11146 9985
rect 11088 9945 11100 9979
rect 11134 9976 11146 9979
rect 12253 9979 12311 9985
rect 11134 9948 11836 9976
rect 11134 9945 11146 9948
rect 11088 9939 11146 9945
rect 11808 9917 11836 9948
rect 12253 9945 12265 9979
rect 12299 9945 12311 9979
rect 19812 9976 19840 10007
rect 23014 10004 23020 10016
rect 23072 10004 23078 10056
rect 27249 10047 27307 10053
rect 20806 9976 20812 9988
rect 19812 9948 20812 9976
rect 12253 9939 12311 9945
rect 20806 9936 20812 9948
rect 20864 9936 20870 9988
rect 21266 9936 21272 9988
rect 21324 9936 21330 9988
rect 21818 9936 21824 9988
rect 21876 9976 21882 9988
rect 23124 9976 23152 10030
rect 27249 10013 27261 10047
rect 27295 10044 27307 10047
rect 27614 10044 27620 10056
rect 27295 10016 27620 10044
rect 27295 10013 27307 10016
rect 27249 10007 27307 10013
rect 27614 10004 27620 10016
rect 27672 10004 27678 10056
rect 25958 9976 25964 9988
rect 21876 9948 25964 9976
rect 21876 9936 21882 9948
rect 25958 9936 25964 9948
rect 26016 9936 26022 9988
rect 4264 9880 7512 9908
rect 11793 9911 11851 9917
rect 11793 9877 11805 9911
rect 11839 9877 11851 9911
rect 12158 9908 12164 9920
rect 12119 9880 12164 9908
rect 11793 9871 11851 9877
rect 12158 9868 12164 9880
rect 12216 9868 12222 9920
rect 19334 9868 19340 9920
rect 19392 9908 19398 9920
rect 19705 9911 19763 9917
rect 19705 9908 19717 9911
rect 19392 9880 19717 9908
rect 19392 9868 19398 9880
rect 19705 9877 19717 9880
rect 19751 9877 19763 9911
rect 19705 9871 19763 9877
rect 1104 9818 29048 9840
rect 1104 9766 7896 9818
rect 7948 9766 7960 9818
rect 8012 9766 8024 9818
rect 8076 9766 8088 9818
rect 8140 9766 8152 9818
rect 8204 9766 14842 9818
rect 14894 9766 14906 9818
rect 14958 9766 14970 9818
rect 15022 9766 15034 9818
rect 15086 9766 15098 9818
rect 15150 9766 21788 9818
rect 21840 9766 21852 9818
rect 21904 9766 21916 9818
rect 21968 9766 21980 9818
rect 22032 9766 22044 9818
rect 22096 9766 28734 9818
rect 28786 9766 28798 9818
rect 28850 9766 28862 9818
rect 28914 9766 28926 9818
rect 28978 9766 28990 9818
rect 29042 9766 29048 9818
rect 1104 9744 29048 9766
rect 26510 9704 26516 9716
rect 26471 9676 26516 9704
rect 26510 9664 26516 9676
rect 26568 9664 26574 9716
rect 27614 9704 27620 9716
rect 27575 9676 27620 9704
rect 27614 9664 27620 9676
rect 27672 9664 27678 9716
rect 4338 9596 4344 9648
rect 4396 9636 4402 9648
rect 4617 9639 4675 9645
rect 4617 9636 4629 9639
rect 4396 9608 4629 9636
rect 4396 9596 4402 9608
rect 4617 9605 4629 9608
rect 4663 9605 4675 9639
rect 4617 9599 4675 9605
rect 9677 9639 9735 9645
rect 9677 9605 9689 9639
rect 9723 9636 9735 9639
rect 10594 9636 10600 9648
rect 9723 9608 10364 9636
rect 10555 9608 10600 9636
rect 9723 9605 9735 9608
rect 9677 9599 9735 9605
rect 2774 9528 2780 9580
rect 2832 9568 2838 9580
rect 4062 9568 4068 9580
rect 2832 9540 4068 9568
rect 2832 9528 2838 9540
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 5626 9568 5632 9580
rect 4755 9540 5632 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 9582 9568 9588 9580
rect 9543 9540 9588 9568
rect 9582 9528 9588 9540
rect 9640 9528 9646 9580
rect 9766 9568 9772 9580
rect 9727 9540 9772 9568
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 10226 9568 10232 9580
rect 10187 9540 10232 9568
rect 10226 9528 10232 9540
rect 10284 9528 10290 9580
rect 10336 9577 10364 9608
rect 10594 9596 10600 9608
rect 10652 9596 10658 9648
rect 19245 9639 19303 9645
rect 19245 9605 19257 9639
rect 19291 9636 19303 9639
rect 19334 9636 19340 9648
rect 19291 9608 19340 9636
rect 19291 9605 19303 9608
rect 19245 9599 19303 9605
rect 19334 9596 19340 9608
rect 19392 9596 19398 9648
rect 20622 9596 20628 9648
rect 20680 9636 20686 9648
rect 23014 9636 23020 9648
rect 20680 9608 23020 9636
rect 20680 9596 20686 9608
rect 23014 9596 23020 9608
rect 23072 9596 23078 9648
rect 10322 9571 10380 9577
rect 10322 9537 10334 9571
rect 10368 9537 10380 9571
rect 10322 9531 10380 9537
rect 10502 9528 10508 9580
rect 10560 9568 10566 9580
rect 10735 9571 10793 9577
rect 10560 9540 10605 9568
rect 10560 9528 10566 9540
rect 10735 9537 10747 9571
rect 10781 9568 10793 9571
rect 10870 9568 10876 9580
rect 10781 9540 10876 9568
rect 10781 9537 10793 9540
rect 10735 9531 10793 9537
rect 10870 9528 10876 9540
rect 10928 9528 10934 9580
rect 14642 9528 14648 9580
rect 14700 9568 14706 9580
rect 14921 9571 14979 9577
rect 14921 9568 14933 9571
rect 14700 9540 14933 9568
rect 14700 9528 14706 9540
rect 14921 9537 14933 9540
rect 14967 9568 14979 9571
rect 15102 9568 15108 9580
rect 14967 9540 15108 9568
rect 14967 9537 14979 9540
rect 14921 9531 14979 9537
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 17497 9571 17555 9577
rect 17497 9537 17509 9571
rect 17543 9568 17555 9571
rect 18506 9568 18512 9580
rect 17543 9540 18512 9568
rect 17543 9537 17555 9540
rect 17497 9531 17555 9537
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 20346 9528 20352 9580
rect 20404 9528 20410 9580
rect 4890 9460 4896 9512
rect 4948 9500 4954 9512
rect 4948 9472 12434 9500
rect 4948 9460 4954 9472
rect 10778 9392 10784 9444
rect 10836 9432 10842 9444
rect 10873 9435 10931 9441
rect 10873 9432 10885 9435
rect 10836 9404 10885 9432
rect 10836 9392 10842 9404
rect 10873 9401 10885 9404
rect 10919 9401 10931 9435
rect 12406 9432 12434 9472
rect 18782 9460 18788 9512
rect 18840 9500 18846 9512
rect 18969 9503 19027 9509
rect 18969 9500 18981 9503
rect 18840 9472 18981 9500
rect 18840 9460 18846 9472
rect 18969 9469 18981 9472
rect 19015 9469 19027 9503
rect 18969 9463 19027 9469
rect 19794 9460 19800 9512
rect 19852 9500 19858 9512
rect 20640 9500 20668 9596
rect 26418 9568 26424 9580
rect 26379 9540 26424 9568
rect 26418 9528 26424 9540
rect 26476 9528 26482 9580
rect 26602 9568 26608 9580
rect 26563 9540 26608 9568
rect 26602 9528 26608 9540
rect 26660 9528 26666 9580
rect 19852 9472 20668 9500
rect 20717 9503 20775 9509
rect 19852 9460 19858 9472
rect 20717 9469 20729 9503
rect 20763 9500 20775 9503
rect 20806 9500 20812 9512
rect 20763 9472 20812 9500
rect 20763 9469 20775 9472
rect 20717 9463 20775 9469
rect 20806 9460 20812 9472
rect 20864 9460 20870 9512
rect 27157 9503 27215 9509
rect 27157 9469 27169 9503
rect 27203 9500 27215 9503
rect 27246 9500 27252 9512
rect 27203 9472 27252 9500
rect 27203 9469 27215 9472
rect 27157 9463 27215 9469
rect 27246 9460 27252 9472
rect 27304 9460 27310 9512
rect 27525 9435 27583 9441
rect 12406 9404 19104 9432
rect 10873 9395 10931 9401
rect 2590 9324 2596 9376
rect 2648 9364 2654 9376
rect 2685 9367 2743 9373
rect 2685 9364 2697 9367
rect 2648 9336 2697 9364
rect 2648 9324 2654 9336
rect 2685 9333 2697 9336
rect 2731 9333 2743 9367
rect 2685 9327 2743 9333
rect 14366 9324 14372 9376
rect 14424 9364 14430 9376
rect 14829 9367 14887 9373
rect 14829 9364 14841 9367
rect 14424 9336 14841 9364
rect 14424 9324 14430 9336
rect 14829 9333 14841 9336
rect 14875 9333 14887 9367
rect 14829 9327 14887 9333
rect 17126 9324 17132 9376
rect 17184 9364 17190 9376
rect 17405 9367 17463 9373
rect 17405 9364 17417 9367
rect 17184 9336 17417 9364
rect 17184 9324 17190 9336
rect 17405 9333 17417 9336
rect 17451 9333 17463 9367
rect 19076 9364 19104 9404
rect 27525 9401 27537 9435
rect 27571 9432 27583 9435
rect 27798 9432 27804 9444
rect 27571 9404 27804 9432
rect 27571 9401 27583 9404
rect 27525 9395 27583 9401
rect 27798 9392 27804 9404
rect 27856 9392 27862 9444
rect 20254 9364 20260 9376
rect 19076 9336 20260 9364
rect 17405 9327 17463 9333
rect 20254 9324 20260 9336
rect 20312 9324 20318 9376
rect 1104 9274 28888 9296
rect 1104 9222 4423 9274
rect 4475 9222 4487 9274
rect 4539 9222 4551 9274
rect 4603 9222 4615 9274
rect 4667 9222 4679 9274
rect 4731 9222 11369 9274
rect 11421 9222 11433 9274
rect 11485 9222 11497 9274
rect 11549 9222 11561 9274
rect 11613 9222 11625 9274
rect 11677 9222 18315 9274
rect 18367 9222 18379 9274
rect 18431 9222 18443 9274
rect 18495 9222 18507 9274
rect 18559 9222 18571 9274
rect 18623 9222 25261 9274
rect 25313 9222 25325 9274
rect 25377 9222 25389 9274
rect 25441 9222 25453 9274
rect 25505 9222 25517 9274
rect 25569 9222 28888 9274
rect 1104 9200 28888 9222
rect 10502 9160 10508 9172
rect 10463 9132 10508 9160
rect 10502 9120 10508 9132
rect 10560 9120 10566 9172
rect 18782 9160 18788 9172
rect 18743 9132 18788 9160
rect 18782 9120 18788 9132
rect 18840 9120 18846 9172
rect 26878 9160 26884 9172
rect 26839 9132 26884 9160
rect 26878 9120 26884 9132
rect 26936 9120 26942 9172
rect 9585 9095 9643 9101
rect 9585 9061 9597 9095
rect 9631 9092 9643 9095
rect 10594 9092 10600 9104
rect 9631 9064 10600 9092
rect 9631 9061 9643 9064
rect 9585 9055 9643 9061
rect 10594 9052 10600 9064
rect 10652 9052 10658 9104
rect 25774 9092 25780 9104
rect 12406 9064 25780 9092
rect 2682 9024 2688 9036
rect 2643 8996 2688 9024
rect 2682 8984 2688 8996
rect 2740 9024 2746 9036
rect 4154 9024 4160 9036
rect 2740 8996 4160 9024
rect 2740 8984 2746 8996
rect 4154 8984 4160 8996
rect 4212 9024 4218 9036
rect 5534 9024 5540 9036
rect 4212 8996 5540 9024
rect 4212 8984 4218 8996
rect 5534 8984 5540 8996
rect 5592 8984 5598 9036
rect 7006 9024 7012 9036
rect 6967 8996 7012 9024
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 7282 9024 7288 9036
rect 7243 8996 7288 9024
rect 7282 8984 7288 8996
rect 7340 8984 7346 9036
rect 11514 9024 11520 9036
rect 9692 8996 11520 9024
rect 2498 8916 2504 8968
rect 2556 8956 2562 8968
rect 2593 8959 2651 8965
rect 2593 8956 2605 8959
rect 2556 8928 2605 8956
rect 2556 8916 2562 8928
rect 2593 8925 2605 8928
rect 2639 8956 2651 8959
rect 4246 8956 4252 8968
rect 2639 8928 4252 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 4246 8916 4252 8928
rect 4304 8916 4310 8968
rect 6914 8956 6920 8968
rect 6875 8928 6920 8956
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 9692 8965 9720 8996
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 11698 9024 11704 9036
rect 11659 8996 11704 9024
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 9493 8959 9551 8965
rect 9493 8956 9505 8959
rect 9456 8928 9505 8956
rect 9456 8916 9462 8928
rect 9493 8925 9505 8928
rect 9539 8925 9551 8959
rect 9493 8919 9551 8925
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8925 9735 8959
rect 9677 8919 9735 8925
rect 9766 8916 9772 8968
rect 9824 8956 9830 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9824 8928 10149 8956
rect 9824 8916 9830 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8956 11483 8959
rect 12158 8956 12164 8968
rect 11471 8928 12164 8956
rect 11471 8925 11483 8928
rect 11425 8919 11483 8925
rect 12158 8916 12164 8928
rect 12216 8916 12222 8968
rect 4062 8848 4068 8900
rect 4120 8888 4126 8900
rect 9582 8888 9588 8900
rect 4120 8860 9588 8888
rect 4120 8848 4126 8860
rect 9582 8848 9588 8860
rect 9640 8888 9646 8900
rect 10321 8891 10379 8897
rect 10321 8888 10333 8891
rect 9640 8860 10333 8888
rect 9640 8848 9646 8860
rect 10321 8857 10333 8860
rect 10367 8857 10379 8891
rect 12406 8888 12434 9064
rect 17773 9027 17831 9033
rect 17773 8993 17785 9027
rect 17819 8993 17831 9027
rect 17773 8987 17831 8993
rect 14182 8916 14188 8968
rect 14240 8956 14246 8968
rect 14369 8959 14427 8965
rect 14369 8956 14381 8959
rect 14240 8928 14381 8956
rect 14240 8916 14246 8928
rect 14369 8925 14381 8928
rect 14415 8925 14427 8959
rect 14369 8919 14427 8925
rect 14642 8916 14648 8968
rect 14700 8916 14706 8968
rect 15102 8916 15108 8968
rect 15160 8956 15166 8968
rect 15838 8956 15844 8968
rect 15160 8928 15844 8956
rect 15160 8916 15166 8928
rect 15838 8916 15844 8928
rect 15896 8956 15902 8968
rect 15933 8959 15991 8965
rect 15933 8956 15945 8959
rect 15896 8928 15945 8956
rect 15896 8916 15902 8928
rect 15933 8925 15945 8928
rect 15979 8925 15991 8959
rect 15933 8919 15991 8925
rect 15378 8888 15384 8900
rect 10321 8851 10379 8857
rect 10428 8860 12434 8888
rect 15339 8860 15384 8888
rect 3326 8780 3332 8832
rect 3384 8820 3390 8832
rect 3421 8823 3479 8829
rect 3421 8820 3433 8823
rect 3384 8792 3433 8820
rect 3384 8780 3390 8792
rect 3421 8789 3433 8792
rect 3467 8789 3479 8823
rect 3421 8783 3479 8789
rect 5442 8780 5448 8832
rect 5500 8820 5506 8832
rect 10428 8820 10456 8860
rect 15378 8848 15384 8860
rect 15436 8848 15442 8900
rect 16666 8848 16672 8900
rect 16724 8888 16730 8900
rect 17788 8888 17816 8987
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8956 18291 8959
rect 18524 8956 18552 9064
rect 25774 9052 25780 9064
rect 25832 9052 25838 9104
rect 27430 9052 27436 9104
rect 27488 9092 27494 9104
rect 27985 9095 28043 9101
rect 27985 9092 27997 9095
rect 27488 9064 27997 9092
rect 27488 9052 27494 9064
rect 27985 9061 27997 9064
rect 28031 9061 28043 9095
rect 27985 9055 28043 9061
rect 19705 9027 19763 9033
rect 19705 9024 19717 9027
rect 19536 8996 19717 9024
rect 18690 8956 18696 8968
rect 18279 8928 18552 8956
rect 18651 8928 18696 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 18690 8916 18696 8928
rect 18748 8916 18754 8968
rect 19536 8888 19564 8996
rect 19705 8993 19717 8996
rect 19751 9024 19763 9027
rect 19794 9024 19800 9036
rect 19751 8996 19800 9024
rect 19751 8993 19763 8996
rect 19705 8987 19763 8993
rect 19794 8984 19800 8996
rect 19852 8984 19858 9036
rect 20346 8984 20352 9036
rect 20404 9024 20410 9036
rect 20441 9027 20499 9033
rect 20441 9024 20453 9027
rect 20404 8996 20453 9024
rect 20404 8984 20410 8996
rect 20441 8993 20453 8996
rect 20487 8993 20499 9027
rect 20441 8987 20499 8993
rect 22278 8984 22284 9036
rect 22336 9024 22342 9036
rect 22738 9024 22744 9036
rect 22336 8996 22744 9024
rect 22336 8984 22342 8996
rect 22738 8984 22744 8996
rect 22796 9024 22802 9036
rect 23842 9024 23848 9036
rect 22796 8996 22876 9024
rect 23803 8996 23848 9024
rect 22796 8984 22802 8996
rect 20168 8968 20220 8974
rect 20254 8916 20260 8968
rect 20312 8956 20318 8968
rect 22848 8965 22876 8996
rect 23842 8984 23848 8996
rect 23900 8984 23906 9036
rect 26602 8984 26608 9036
rect 26660 9024 26666 9036
rect 27893 9027 27951 9033
rect 27893 9024 27905 9027
rect 26660 8996 27905 9024
rect 26660 8984 26666 8996
rect 22649 8959 22707 8965
rect 22649 8956 22661 8959
rect 20312 8928 22661 8956
rect 20312 8916 20318 8928
rect 22649 8925 22661 8928
rect 22695 8925 22707 8959
rect 22649 8919 22707 8925
rect 22833 8959 22891 8965
rect 22833 8925 22845 8959
rect 22879 8925 22891 8959
rect 23658 8956 23664 8968
rect 23619 8928 23664 8956
rect 22833 8919 22891 8925
rect 23658 8916 23664 8928
rect 23716 8916 23722 8968
rect 26418 8916 26424 8968
rect 26476 8956 26482 8968
rect 27172 8965 27200 8996
rect 27893 8993 27905 8996
rect 27939 8993 27951 9027
rect 27893 8987 27951 8993
rect 27065 8959 27123 8965
rect 27065 8956 27077 8959
rect 26476 8928 27077 8956
rect 26476 8916 26482 8928
rect 27065 8925 27077 8928
rect 27111 8925 27123 8959
rect 27065 8919 27123 8925
rect 27157 8959 27215 8965
rect 27157 8925 27169 8959
rect 27203 8925 27215 8959
rect 27157 8919 27215 8925
rect 27246 8916 27252 8968
rect 27304 8956 27310 8968
rect 27377 8959 27435 8965
rect 27304 8928 27349 8956
rect 27304 8916 27310 8928
rect 27377 8925 27389 8959
rect 27423 8956 27435 8959
rect 27798 8956 27804 8968
rect 27423 8928 27804 8956
rect 27423 8925 27435 8928
rect 27377 8919 27435 8925
rect 27798 8916 27804 8928
rect 27856 8916 27862 8968
rect 20168 8910 20220 8916
rect 28350 8888 28356 8900
rect 16724 8860 19564 8888
rect 28311 8860 28356 8888
rect 16724 8848 16730 8860
rect 28350 8848 28356 8860
rect 28408 8848 28414 8900
rect 11054 8820 11060 8832
rect 5500 8792 10456 8820
rect 11015 8792 11060 8820
rect 5500 8780 5506 8792
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 11514 8780 11520 8832
rect 11572 8820 11578 8832
rect 12158 8820 12164 8832
rect 11572 8792 12164 8820
rect 11572 8780 11578 8792
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 16025 8823 16083 8829
rect 16025 8789 16037 8823
rect 16071 8820 16083 8823
rect 16850 8820 16856 8832
rect 16071 8792 16856 8820
rect 16071 8789 16083 8792
rect 16025 8783 16083 8789
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 22830 8820 22836 8832
rect 22791 8792 22836 8820
rect 22830 8780 22836 8792
rect 22888 8780 22894 8832
rect 23106 8780 23112 8832
rect 23164 8820 23170 8832
rect 23293 8823 23351 8829
rect 23293 8820 23305 8823
rect 23164 8792 23305 8820
rect 23164 8780 23170 8792
rect 23293 8789 23305 8792
rect 23339 8789 23351 8823
rect 23293 8783 23351 8789
rect 23753 8823 23811 8829
rect 23753 8789 23765 8823
rect 23799 8820 23811 8823
rect 25130 8820 25136 8832
rect 23799 8792 25136 8820
rect 23799 8789 23811 8792
rect 23753 8783 23811 8789
rect 25130 8780 25136 8792
rect 25188 8780 25194 8832
rect 1104 8730 29048 8752
rect 1104 8678 7896 8730
rect 7948 8678 7960 8730
rect 8012 8678 8024 8730
rect 8076 8678 8088 8730
rect 8140 8678 8152 8730
rect 8204 8678 14842 8730
rect 14894 8678 14906 8730
rect 14958 8678 14970 8730
rect 15022 8678 15034 8730
rect 15086 8678 15098 8730
rect 15150 8678 21788 8730
rect 21840 8678 21852 8730
rect 21904 8678 21916 8730
rect 21968 8678 21980 8730
rect 22032 8678 22044 8730
rect 22096 8678 28734 8730
rect 28786 8678 28798 8730
rect 28850 8678 28862 8730
rect 28914 8678 28926 8730
rect 28978 8678 28990 8730
rect 29042 8678 29048 8730
rect 1104 8656 29048 8678
rect 4062 8616 4068 8628
rect 4023 8588 4068 8616
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 7006 8576 7012 8628
rect 7064 8616 7070 8628
rect 7742 8616 7748 8628
rect 7064 8588 7748 8616
rect 7064 8576 7070 8588
rect 7742 8576 7748 8588
rect 7800 8616 7806 8628
rect 8113 8619 8171 8625
rect 8113 8616 8125 8619
rect 7800 8588 8125 8616
rect 7800 8576 7806 8588
rect 8113 8585 8125 8588
rect 8159 8585 8171 8619
rect 10870 8616 10876 8628
rect 10831 8588 10876 8616
rect 8113 8579 8171 8585
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 15838 8616 15844 8628
rect 15799 8588 15844 8616
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 18601 8619 18659 8625
rect 18601 8585 18613 8619
rect 18647 8616 18659 8619
rect 18690 8616 18696 8628
rect 18647 8588 18696 8616
rect 18647 8585 18659 8588
rect 18601 8579 18659 8585
rect 18690 8576 18696 8588
rect 18748 8576 18754 8628
rect 22830 8576 22836 8628
rect 22888 8616 22894 8628
rect 24581 8619 24639 8625
rect 22888 8588 23520 8616
rect 22888 8576 22894 8588
rect 2590 8548 2596 8560
rect 2551 8520 2596 8548
rect 2590 8508 2596 8520
rect 2648 8508 2654 8560
rect 3326 8508 3332 8560
rect 3384 8508 3390 8560
rect 10505 8551 10563 8557
rect 10505 8517 10517 8551
rect 10551 8548 10563 8551
rect 11514 8548 11520 8560
rect 10551 8520 11520 8548
rect 10551 8517 10563 8520
rect 10505 8511 10563 8517
rect 11514 8508 11520 8520
rect 11572 8508 11578 8560
rect 14366 8548 14372 8560
rect 14327 8520 14372 8548
rect 14366 8508 14372 8520
rect 14424 8508 14430 8560
rect 15378 8508 15384 8560
rect 15436 8508 15442 8560
rect 17126 8548 17132 8560
rect 17087 8520 17132 8548
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 18138 8508 18144 8560
rect 18196 8508 18202 8560
rect 23106 8548 23112 8560
rect 23067 8520 23112 8548
rect 23106 8508 23112 8520
rect 23164 8508 23170 8560
rect 23492 8548 23520 8588
rect 24581 8585 24593 8619
rect 24627 8616 24639 8619
rect 25130 8616 25136 8628
rect 24627 8588 25136 8616
rect 24627 8585 24639 8588
rect 24581 8579 24639 8585
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 27709 8619 27767 8625
rect 27709 8585 27721 8619
rect 27755 8616 27767 8619
rect 27890 8616 27896 8628
rect 27755 8588 27896 8616
rect 27755 8585 27767 8588
rect 27709 8579 27767 8585
rect 27890 8576 27896 8588
rect 27948 8576 27954 8628
rect 23492 8520 23598 8548
rect 4982 8440 4988 8492
rect 5040 8480 5046 8492
rect 5718 8480 5724 8492
rect 5040 8452 5724 8480
rect 5040 8440 5046 8452
rect 5718 8440 5724 8452
rect 5776 8480 5782 8492
rect 6733 8483 6791 8489
rect 6733 8480 6745 8483
rect 5776 8452 6745 8480
rect 5776 8440 5782 8452
rect 6733 8449 6745 8452
rect 6779 8449 6791 8483
rect 6733 8443 6791 8449
rect 7000 8483 7058 8489
rect 7000 8449 7012 8483
rect 7046 8480 7058 8483
rect 7374 8480 7380 8492
rect 7046 8452 7380 8480
rect 7046 8449 7058 8452
rect 7000 8443 7058 8449
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 9398 8440 9404 8492
rect 9456 8480 9462 8492
rect 10689 8483 10747 8489
rect 10689 8480 10701 8483
rect 9456 8452 10701 8480
rect 9456 8440 9462 8452
rect 10689 8449 10701 8452
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 10778 8440 10784 8492
rect 10836 8480 10842 8492
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 10836 8452 11713 8480
rect 10836 8440 10842 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 11790 8440 11796 8492
rect 11848 8480 11854 8492
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 11848 8452 11897 8480
rect 11848 8440 11854 8452
rect 11885 8449 11897 8452
rect 11931 8449 11943 8483
rect 13630 8480 13636 8492
rect 13591 8452 13636 8480
rect 11885 8443 11943 8449
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 16850 8480 16856 8492
rect 16811 8452 16856 8480
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 22738 8440 22744 8492
rect 22796 8480 22802 8492
rect 22833 8483 22891 8489
rect 22833 8480 22845 8483
rect 22796 8452 22845 8480
rect 22796 8440 22802 8452
rect 22833 8449 22845 8452
rect 22879 8449 22891 8483
rect 22833 8443 22891 8449
rect 27341 8483 27399 8489
rect 27341 8449 27353 8483
rect 27387 8480 27399 8483
rect 27522 8480 27528 8492
rect 27387 8452 27528 8480
rect 27387 8449 27399 8452
rect 27341 8443 27399 8449
rect 27522 8440 27528 8452
rect 27580 8480 27586 8492
rect 28350 8480 28356 8492
rect 27580 8452 28356 8480
rect 27580 8440 27586 8452
rect 28350 8440 28356 8452
rect 28408 8440 28414 8492
rect 2314 8412 2320 8424
rect 2275 8384 2320 8412
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 13541 8415 13599 8421
rect 13541 8381 13553 8415
rect 13587 8412 13599 8415
rect 14093 8415 14151 8421
rect 14093 8412 14105 8415
rect 13587 8384 14105 8412
rect 13587 8381 13599 8384
rect 13541 8375 13599 8381
rect 14093 8381 14105 8384
rect 14139 8381 14151 8415
rect 27430 8412 27436 8424
rect 27391 8384 27436 8412
rect 14093 8375 14151 8381
rect 27430 8372 27436 8384
rect 27488 8372 27494 8424
rect 11882 8344 11888 8356
rect 11843 8316 11888 8344
rect 11882 8304 11888 8316
rect 11940 8304 11946 8356
rect 1104 8186 28888 8208
rect 1104 8134 4423 8186
rect 4475 8134 4487 8186
rect 4539 8134 4551 8186
rect 4603 8134 4615 8186
rect 4667 8134 4679 8186
rect 4731 8134 11369 8186
rect 11421 8134 11433 8186
rect 11485 8134 11497 8186
rect 11549 8134 11561 8186
rect 11613 8134 11625 8186
rect 11677 8134 18315 8186
rect 18367 8134 18379 8186
rect 18431 8134 18443 8186
rect 18495 8134 18507 8186
rect 18559 8134 18571 8186
rect 18623 8134 25261 8186
rect 25313 8134 25325 8186
rect 25377 8134 25389 8186
rect 25441 8134 25453 8186
rect 25505 8134 25517 8186
rect 25569 8134 28888 8186
rect 1104 8112 28888 8134
rect 2314 8032 2320 8084
rect 2372 8072 2378 8084
rect 2593 8075 2651 8081
rect 2593 8072 2605 8075
rect 2372 8044 2605 8072
rect 2372 8032 2378 8044
rect 2593 8041 2605 8044
rect 2639 8041 2651 8075
rect 2593 8035 2651 8041
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 5813 8075 5871 8081
rect 5813 8072 5825 8075
rect 5592 8044 5825 8072
rect 5592 8032 5598 8044
rect 5813 8041 5825 8044
rect 5859 8041 5871 8075
rect 9306 8072 9312 8084
rect 9267 8044 9312 8072
rect 5813 8035 5871 8041
rect 9306 8032 9312 8044
rect 9364 8032 9370 8084
rect 12158 8072 12164 8084
rect 12119 8044 12164 8072
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 13630 8032 13636 8084
rect 13688 8072 13694 8084
rect 15654 8072 15660 8084
rect 13688 8044 15660 8072
rect 13688 8032 13694 8044
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7936 9551 7939
rect 10686 7936 10692 7948
rect 9539 7908 10692 7936
rect 9539 7905 9551 7908
rect 9493 7899 9551 7905
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7868 2743 7871
rect 3326 7868 3332 7880
rect 2731 7840 3332 7868
rect 2731 7837 2743 7840
rect 2685 7831 2743 7837
rect 3326 7828 3332 7840
rect 3384 7828 3390 7880
rect 8478 7868 8484 7880
rect 8439 7840 8484 7868
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9309 7871 9367 7877
rect 9309 7868 9321 7871
rect 9088 7840 9321 7868
rect 9088 7828 9094 7840
rect 9309 7837 9321 7840
rect 9355 7837 9367 7871
rect 9309 7831 9367 7837
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7868 10839 7871
rect 10870 7868 10876 7880
rect 10827 7840 10876 7868
rect 10827 7837 10839 7840
rect 10781 7831 10839 7837
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 11054 7877 11060 7880
rect 11048 7868 11060 7877
rect 11015 7840 11060 7868
rect 11048 7831 11060 7840
rect 11054 7828 11060 7831
rect 11112 7828 11118 7880
rect 13740 7877 13768 8044
rect 15654 8032 15660 8044
rect 15712 8072 15718 8084
rect 16025 8075 16083 8081
rect 16025 8072 16037 8075
rect 15712 8044 16037 8072
rect 15712 8032 15718 8044
rect 16025 8041 16037 8044
rect 16071 8041 16083 8075
rect 16025 8035 16083 8041
rect 26789 8075 26847 8081
rect 26789 8041 26801 8075
rect 26835 8072 26847 8075
rect 27246 8072 27252 8084
rect 26835 8044 27252 8072
rect 26835 8041 26847 8044
rect 26789 8035 26847 8041
rect 27246 8032 27252 8044
rect 27304 8032 27310 8084
rect 27798 8072 27804 8084
rect 27759 8044 27804 8072
rect 27798 8032 27804 8044
rect 27856 8032 27862 8084
rect 14642 7896 14648 7948
rect 14700 7936 14706 7948
rect 17681 7939 17739 7945
rect 14700 7908 17356 7936
rect 14700 7896 14706 7908
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 13964 7840 14289 7868
rect 13964 7828 13970 7840
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 16666 7868 16672 7880
rect 16627 7840 16672 7868
rect 14277 7831 14335 7837
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 17328 7868 17356 7908
rect 17681 7905 17693 7939
rect 17727 7936 17739 7939
rect 18138 7936 18144 7948
rect 17727 7908 18144 7936
rect 17727 7905 17739 7908
rect 17681 7899 17739 7905
rect 18138 7896 18144 7908
rect 18196 7896 18202 7948
rect 19978 7896 19984 7948
rect 20036 7936 20042 7948
rect 20257 7939 20315 7945
rect 20257 7936 20269 7939
rect 20036 7908 20269 7936
rect 20036 7896 20042 7908
rect 20257 7905 20269 7908
rect 20303 7905 20315 7939
rect 20257 7899 20315 7905
rect 21634 7896 21640 7948
rect 21692 7936 21698 7948
rect 22186 7936 22192 7948
rect 21692 7908 22192 7936
rect 21692 7896 21698 7908
rect 22186 7896 22192 7908
rect 22244 7936 22250 7948
rect 22244 7908 24624 7936
rect 22244 7896 22250 7908
rect 19334 7868 19340 7880
rect 17328 7854 19340 7868
rect 17342 7840 19340 7854
rect 19334 7828 19340 7840
rect 19392 7828 19398 7880
rect 24596 7877 24624 7908
rect 26252 7908 27292 7936
rect 24581 7871 24639 7877
rect 24581 7837 24593 7871
rect 24627 7837 24639 7871
rect 24762 7868 24768 7880
rect 24723 7840 24768 7868
rect 24581 7831 24639 7837
rect 24762 7828 24768 7840
rect 24820 7828 24826 7880
rect 4525 7803 4583 7809
rect 4525 7769 4537 7803
rect 4571 7800 4583 7803
rect 6914 7800 6920 7812
rect 4571 7772 6920 7800
rect 4571 7769 4583 7772
rect 4525 7763 4583 7769
rect 6914 7760 6920 7772
rect 6972 7760 6978 7812
rect 9582 7800 9588 7812
rect 9543 7772 9588 7800
rect 9582 7760 9588 7772
rect 9640 7760 9646 7812
rect 13633 7803 13691 7809
rect 13633 7769 13645 7803
rect 13679 7800 13691 7803
rect 14553 7803 14611 7809
rect 14553 7800 14565 7803
rect 13679 7772 14565 7800
rect 13679 7769 13691 7772
rect 13633 7763 13691 7769
rect 14553 7769 14565 7772
rect 14599 7769 14611 7803
rect 14553 7763 14611 7769
rect 15194 7760 15200 7812
rect 15252 7760 15258 7812
rect 20524 7803 20582 7809
rect 20524 7769 20536 7803
rect 20570 7800 20582 7803
rect 21174 7800 21180 7812
rect 20570 7772 21180 7800
rect 20570 7769 20582 7772
rect 20524 7763 20582 7769
rect 21174 7760 21180 7772
rect 21232 7760 21238 7812
rect 22462 7800 22468 7812
rect 22423 7772 22468 7800
rect 22462 7760 22468 7772
rect 22520 7760 22526 7812
rect 24673 7803 24731 7809
rect 24673 7800 24685 7803
rect 23690 7772 24685 7800
rect 24673 7769 24685 7772
rect 24719 7769 24731 7803
rect 24673 7763 24731 7769
rect 25958 7760 25964 7812
rect 26016 7800 26022 7812
rect 26252 7809 26280 7908
rect 27264 7877 27292 7908
rect 27356 7908 27660 7936
rect 27249 7871 27307 7877
rect 27249 7837 27261 7871
rect 27295 7837 27307 7871
rect 27249 7831 27307 7837
rect 26237 7803 26295 7809
rect 26237 7800 26249 7803
rect 26016 7772 26249 7800
rect 26016 7760 26022 7772
rect 26237 7769 26249 7772
rect 26283 7769 26295 7803
rect 26237 7763 26295 7769
rect 26513 7803 26571 7809
rect 26513 7769 26525 7803
rect 26559 7800 26571 7803
rect 27356 7800 27384 7908
rect 27632 7877 27660 7908
rect 27617 7871 27675 7877
rect 27617 7837 27629 7871
rect 27663 7868 27675 7871
rect 27982 7868 27988 7880
rect 27663 7840 27988 7868
rect 27663 7837 27675 7840
rect 27617 7831 27675 7837
rect 27982 7828 27988 7840
rect 28040 7828 28046 7880
rect 26559 7772 27384 7800
rect 27433 7803 27491 7809
rect 26559 7769 26571 7772
rect 26513 7763 26571 7769
rect 27433 7769 27445 7803
rect 27479 7769 27491 7803
rect 27433 7763 27491 7769
rect 27525 7803 27583 7809
rect 27525 7769 27537 7803
rect 27571 7769 27583 7803
rect 27525 7763 27583 7769
rect 2406 7692 2412 7744
rect 2464 7732 2470 7744
rect 3237 7735 3295 7741
rect 3237 7732 3249 7735
rect 2464 7704 3249 7732
rect 2464 7692 2470 7704
rect 3237 7701 3249 7704
rect 3283 7701 3295 7735
rect 9122 7732 9128 7744
rect 9083 7704 9128 7732
rect 3237 7695 3295 7701
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 21637 7735 21695 7741
rect 21637 7701 21649 7735
rect 21683 7732 21695 7735
rect 22186 7732 22192 7744
rect 21683 7704 22192 7732
rect 21683 7701 21695 7704
rect 21637 7695 21695 7701
rect 22186 7692 22192 7704
rect 22244 7692 22250 7744
rect 23937 7735 23995 7741
rect 23937 7701 23949 7735
rect 23983 7732 23995 7735
rect 25406 7732 25412 7744
rect 23983 7704 25412 7732
rect 23983 7701 23995 7704
rect 23937 7695 23995 7701
rect 25406 7692 25412 7704
rect 25464 7732 25470 7744
rect 25682 7732 25688 7744
rect 25464 7704 25688 7732
rect 25464 7692 25470 7704
rect 25682 7692 25688 7704
rect 25740 7732 25746 7744
rect 26418 7732 26424 7744
rect 25740 7704 26424 7732
rect 25740 7692 25746 7704
rect 26418 7692 26424 7704
rect 26476 7692 26482 7744
rect 26602 7732 26608 7744
rect 26563 7704 26608 7732
rect 26602 7692 26608 7704
rect 26660 7732 26666 7744
rect 27448 7732 27476 7763
rect 26660 7704 27476 7732
rect 27540 7732 27568 7763
rect 27614 7732 27620 7744
rect 27540 7704 27620 7732
rect 26660 7692 26666 7704
rect 27614 7692 27620 7704
rect 27672 7692 27678 7744
rect 1104 7642 29048 7664
rect 1104 7590 7896 7642
rect 7948 7590 7960 7642
rect 8012 7590 8024 7642
rect 8076 7590 8088 7642
rect 8140 7590 8152 7642
rect 8204 7590 14842 7642
rect 14894 7590 14906 7642
rect 14958 7590 14970 7642
rect 15022 7590 15034 7642
rect 15086 7590 15098 7642
rect 15150 7590 21788 7642
rect 21840 7590 21852 7642
rect 21904 7590 21916 7642
rect 21968 7590 21980 7642
rect 22032 7590 22044 7642
rect 22096 7590 28734 7642
rect 28786 7590 28798 7642
rect 28850 7590 28862 7642
rect 28914 7590 28926 7642
rect 28978 7590 28990 7642
rect 29042 7590 29048 7642
rect 1104 7568 29048 7590
rect 3326 7488 3332 7540
rect 3384 7528 3390 7540
rect 3881 7531 3939 7537
rect 3881 7528 3893 7531
rect 3384 7500 3893 7528
rect 3384 7488 3390 7500
rect 3881 7497 3893 7500
rect 3927 7528 3939 7531
rect 7006 7528 7012 7540
rect 3927 7500 7012 7528
rect 3927 7497 3939 7500
rect 3881 7491 3939 7497
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 7374 7528 7380 7540
rect 7335 7500 7380 7528
rect 7374 7488 7380 7500
rect 7432 7488 7438 7540
rect 7742 7488 7748 7540
rect 7800 7528 7806 7540
rect 7837 7531 7895 7537
rect 7837 7528 7849 7531
rect 7800 7500 7849 7528
rect 7800 7488 7806 7500
rect 7837 7497 7849 7500
rect 7883 7497 7895 7531
rect 7837 7491 7895 7497
rect 9490 7488 9496 7540
rect 9548 7528 9554 7540
rect 10321 7531 10379 7537
rect 10321 7528 10333 7531
rect 9548 7500 10333 7528
rect 9548 7488 9554 7500
rect 10321 7497 10333 7500
rect 10367 7497 10379 7531
rect 10321 7491 10379 7497
rect 18693 7531 18751 7537
rect 18693 7497 18705 7531
rect 18739 7528 18751 7531
rect 19334 7528 19340 7540
rect 18739 7500 19340 7528
rect 18739 7497 18751 7500
rect 18693 7491 18751 7497
rect 19334 7488 19340 7500
rect 19392 7528 19398 7540
rect 20162 7528 20168 7540
rect 19392 7500 20168 7528
rect 19392 7488 19398 7500
rect 20162 7488 20168 7500
rect 20220 7488 20226 7540
rect 21174 7528 21180 7540
rect 21135 7500 21180 7528
rect 21174 7488 21180 7500
rect 21232 7488 21238 7540
rect 22462 7488 22468 7540
rect 22520 7528 22526 7540
rect 23201 7531 23259 7537
rect 23201 7528 23213 7531
rect 22520 7500 23213 7528
rect 22520 7488 22526 7500
rect 23201 7497 23213 7500
rect 23247 7497 23259 7531
rect 23566 7528 23572 7540
rect 23527 7500 23572 7528
rect 23201 7491 23259 7497
rect 23566 7488 23572 7500
rect 23624 7488 23630 7540
rect 23661 7531 23719 7537
rect 23661 7497 23673 7531
rect 23707 7528 23719 7531
rect 25406 7528 25412 7540
rect 23707 7500 25412 7528
rect 23707 7497 23719 7500
rect 23661 7491 23719 7497
rect 25406 7488 25412 7500
rect 25464 7488 25470 7540
rect 26329 7531 26387 7537
rect 26329 7497 26341 7531
rect 26375 7528 26387 7531
rect 26418 7528 26424 7540
rect 26375 7500 26424 7528
rect 26375 7497 26387 7500
rect 26329 7491 26387 7497
rect 2406 7460 2412 7472
rect 2367 7432 2412 7460
rect 2406 7420 2412 7432
rect 2464 7420 2470 7472
rect 3418 7420 3424 7472
rect 3476 7420 3482 7472
rect 4700 7463 4758 7469
rect 4700 7429 4712 7463
rect 4746 7460 4758 7463
rect 4890 7460 4896 7472
rect 4746 7432 4896 7460
rect 4746 7429 4758 7432
rect 4700 7423 4758 7429
rect 4890 7420 4896 7432
rect 4948 7420 4954 7472
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7392 4491 7395
rect 4982 7392 4988 7404
rect 4479 7364 4988 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7392 7803 7395
rect 9508 7392 9536 7488
rect 15013 7463 15071 7469
rect 15013 7429 15025 7463
rect 15059 7460 15071 7463
rect 15194 7460 15200 7472
rect 15059 7432 15200 7460
rect 15059 7429 15071 7432
rect 15013 7423 15071 7429
rect 15194 7420 15200 7432
rect 15252 7420 15258 7472
rect 19702 7420 19708 7472
rect 19760 7460 19766 7472
rect 19981 7463 20039 7469
rect 19981 7460 19993 7463
rect 19760 7432 19993 7460
rect 19760 7420 19766 7432
rect 19981 7429 19993 7432
rect 20027 7429 20039 7463
rect 19981 7423 20039 7429
rect 25038 7420 25044 7472
rect 25096 7460 25102 7472
rect 25317 7463 25375 7469
rect 25317 7460 25329 7463
rect 25096 7432 25329 7460
rect 25096 7420 25102 7432
rect 25317 7429 25329 7432
rect 25363 7429 25375 7463
rect 26344 7460 26372 7491
rect 26418 7488 26424 7500
rect 26476 7488 26482 7540
rect 26510 7488 26516 7540
rect 26568 7528 26574 7540
rect 26605 7531 26663 7537
rect 26605 7528 26617 7531
rect 26568 7500 26617 7528
rect 26568 7488 26574 7500
rect 26605 7497 26617 7500
rect 26651 7528 26663 7531
rect 27522 7528 27528 7540
rect 26651 7500 27384 7528
rect 27483 7500 27528 7528
rect 26651 7497 26663 7500
rect 26605 7491 26663 7497
rect 27356 7469 27384 7500
rect 27522 7488 27528 7500
rect 27580 7488 27586 7540
rect 25317 7423 25375 7429
rect 25700 7432 26372 7460
rect 27341 7463 27399 7469
rect 7791 7364 9536 7392
rect 14648 7404 14700 7410
rect 7791 7361 7803 7364
rect 7745 7355 7803 7361
rect 21269 7395 21327 7401
rect 21269 7361 21281 7395
rect 21315 7392 21327 7395
rect 22186 7392 22192 7404
rect 21315 7364 22192 7392
rect 21315 7361 21327 7364
rect 21269 7355 21327 7361
rect 22186 7352 22192 7364
rect 22244 7392 22250 7404
rect 22646 7392 22652 7404
rect 22244 7364 22652 7392
rect 22244 7352 22250 7364
rect 22646 7352 22652 7364
rect 22704 7352 22710 7404
rect 25130 7392 25136 7404
rect 25043 7364 25136 7392
rect 25130 7352 25136 7364
rect 25188 7352 25194 7404
rect 25406 7392 25412 7404
rect 25367 7364 25412 7392
rect 25406 7352 25412 7364
rect 25464 7352 25470 7404
rect 25537 7401 25595 7407
rect 25537 7367 25549 7401
rect 25583 7398 25595 7401
rect 25700 7398 25728 7432
rect 27341 7429 27353 7463
rect 27387 7429 27399 7463
rect 27341 7423 27399 7429
rect 25583 7370 25728 7398
rect 26237 7395 26295 7401
rect 25583 7367 25595 7370
rect 25537 7361 25595 7367
rect 26237 7361 26249 7395
rect 26283 7392 26295 7395
rect 26326 7392 26332 7404
rect 26283 7364 26332 7392
rect 26283 7361 26295 7364
rect 26237 7355 26295 7361
rect 26326 7352 26332 7364
rect 26384 7352 26390 7404
rect 26421 7395 26479 7401
rect 26421 7361 26433 7395
rect 26467 7392 26479 7395
rect 26510 7392 26516 7404
rect 26467 7364 26516 7392
rect 26467 7361 26479 7364
rect 26421 7355 26479 7361
rect 26510 7352 26516 7364
rect 26568 7352 26574 7404
rect 27157 7395 27215 7401
rect 27157 7361 27169 7395
rect 27203 7361 27215 7395
rect 27982 7392 27988 7404
rect 27943 7364 27988 7392
rect 27157 7355 27215 7361
rect 14648 7346 14700 7352
rect 2130 7324 2136 7336
rect 2091 7296 2136 7324
rect 2130 7284 2136 7296
rect 2188 7284 2194 7336
rect 8021 7327 8079 7333
rect 8021 7293 8033 7327
rect 8067 7293 8079 7327
rect 8021 7287 8079 7293
rect 7006 7216 7012 7268
rect 7064 7256 7070 7268
rect 8036 7256 8064 7287
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 10413 7327 10471 7333
rect 10413 7324 10425 7327
rect 9548 7296 10425 7324
rect 9548 7284 9554 7296
rect 10413 7293 10425 7296
rect 10459 7293 10471 7327
rect 10413 7287 10471 7293
rect 10502 7284 10508 7336
rect 10560 7324 10566 7336
rect 10597 7327 10655 7333
rect 10597 7324 10609 7327
rect 10560 7296 10609 7324
rect 10560 7284 10566 7296
rect 10597 7293 10609 7296
rect 10643 7324 10655 7327
rect 11698 7324 11704 7336
rect 10643 7296 11704 7324
rect 10643 7293 10655 7296
rect 10597 7287 10655 7293
rect 11698 7284 11704 7296
rect 11756 7284 11762 7336
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 14182 7324 14188 7336
rect 13872 7296 14188 7324
rect 13872 7284 13878 7296
rect 14182 7284 14188 7296
rect 14240 7284 14246 7336
rect 23842 7324 23848 7336
rect 23803 7296 23848 7324
rect 23842 7284 23848 7296
rect 23900 7284 23906 7336
rect 12342 7256 12348 7268
rect 7064 7228 12348 7256
rect 7064 7216 7070 7228
rect 12342 7216 12348 7228
rect 12400 7216 12406 7268
rect 25148 7256 25176 7352
rect 25225 7327 25283 7333
rect 25225 7293 25237 7327
rect 25271 7324 25283 7327
rect 27172 7324 27200 7355
rect 27982 7352 27988 7364
rect 28040 7352 28046 7404
rect 25271 7296 27200 7324
rect 25271 7293 25283 7296
rect 25225 7287 25283 7293
rect 25958 7256 25964 7268
rect 25148 7228 25964 7256
rect 25958 7216 25964 7228
rect 26016 7256 26022 7268
rect 26053 7259 26111 7265
rect 26053 7256 26065 7259
rect 26016 7228 26065 7256
rect 26016 7216 26022 7228
rect 26053 7225 26065 7228
rect 26099 7225 26111 7259
rect 26053 7219 26111 7225
rect 5810 7188 5816 7200
rect 5771 7160 5816 7188
rect 5810 7148 5816 7160
rect 5868 7148 5874 7200
rect 9953 7191 10011 7197
rect 9953 7157 9965 7191
rect 9999 7188 10011 7191
rect 10594 7188 10600 7200
rect 9999 7160 10600 7188
rect 9999 7157 10011 7160
rect 9953 7151 10011 7157
rect 10594 7148 10600 7160
rect 10652 7148 10658 7200
rect 25038 7148 25044 7200
rect 25096 7188 25102 7200
rect 26510 7188 26516 7200
rect 25096 7160 26516 7188
rect 25096 7148 25102 7160
rect 26510 7148 26516 7160
rect 26568 7148 26574 7200
rect 28074 7188 28080 7200
rect 28035 7160 28080 7188
rect 28074 7148 28080 7160
rect 28132 7148 28138 7200
rect 1104 7098 28888 7120
rect 1104 7046 4423 7098
rect 4475 7046 4487 7098
rect 4539 7046 4551 7098
rect 4603 7046 4615 7098
rect 4667 7046 4679 7098
rect 4731 7046 11369 7098
rect 11421 7046 11433 7098
rect 11485 7046 11497 7098
rect 11549 7046 11561 7098
rect 11613 7046 11625 7098
rect 11677 7046 18315 7098
rect 18367 7046 18379 7098
rect 18431 7046 18443 7098
rect 18495 7046 18507 7098
rect 18559 7046 18571 7098
rect 18623 7046 25261 7098
rect 25313 7046 25325 7098
rect 25377 7046 25389 7098
rect 25441 7046 25453 7098
rect 25505 7046 25517 7098
rect 25569 7046 28888 7098
rect 1104 7024 28888 7046
rect 4890 6984 4896 6996
rect 4851 6956 4896 6984
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 7653 6987 7711 6993
rect 7653 6984 7665 6987
rect 7340 6956 7665 6984
rect 7340 6944 7346 6956
rect 7653 6953 7665 6956
rect 7699 6953 7711 6987
rect 7653 6947 7711 6953
rect 27709 6987 27767 6993
rect 27709 6953 27721 6987
rect 27755 6984 27767 6987
rect 27982 6984 27988 6996
rect 27755 6956 27988 6984
rect 27755 6953 27767 6956
rect 27709 6947 27767 6953
rect 27982 6944 27988 6956
rect 28040 6944 28046 6996
rect 12728 6888 12940 6916
rect 12728 6860 12756 6888
rect 2682 6848 2688 6860
rect 2643 6820 2688 6848
rect 2682 6808 2688 6820
rect 2740 6808 2746 6860
rect 3418 6848 3424 6860
rect 3379 6820 3424 6848
rect 3418 6808 3424 6820
rect 3476 6808 3482 6860
rect 5537 6851 5595 6857
rect 5537 6817 5549 6851
rect 5583 6848 5595 6851
rect 6641 6851 6699 6857
rect 6641 6848 6653 6851
rect 5583 6820 6653 6848
rect 5583 6817 5595 6820
rect 5537 6811 5595 6817
rect 6641 6817 6653 6820
rect 6687 6817 6699 6851
rect 6641 6811 6699 6817
rect 2498 6740 2504 6792
rect 2556 6780 2562 6792
rect 2593 6783 2651 6789
rect 2593 6780 2605 6783
rect 2556 6752 2605 6780
rect 2556 6740 2562 6752
rect 2593 6749 2605 6752
rect 2639 6749 2651 6783
rect 2593 6743 2651 6749
rect 5353 6783 5411 6789
rect 5353 6749 5365 6783
rect 5399 6780 5411 6783
rect 5810 6780 5816 6792
rect 5399 6752 5816 6780
rect 5399 6749 5411 6752
rect 5353 6743 5411 6749
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 6656 6780 6684 6811
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 6788 6820 7757 6848
rect 6788 6808 6794 6820
rect 7745 6817 7757 6820
rect 7791 6817 7803 6851
rect 9122 6848 9128 6860
rect 7745 6811 7803 6817
rect 7852 6820 9128 6848
rect 7006 6780 7012 6792
rect 6656 6752 7012 6780
rect 7006 6740 7012 6752
rect 7064 6740 7070 6792
rect 7653 6783 7711 6789
rect 7653 6749 7665 6783
rect 7699 6780 7711 6783
rect 7852 6780 7880 6820
rect 9122 6808 9128 6820
rect 9180 6808 9186 6860
rect 10870 6848 10876 6860
rect 10831 6820 10876 6848
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 12710 6808 12716 6860
rect 12768 6808 12774 6860
rect 12805 6851 12863 6857
rect 12805 6817 12817 6851
rect 12851 6817 12863 6851
rect 12912 6848 12940 6888
rect 13998 6848 14004 6860
rect 12912 6820 14004 6848
rect 12805 6811 12863 6817
rect 7699 6752 7880 6780
rect 7929 6783 7987 6789
rect 7699 6749 7711 6752
rect 7653 6743 7711 6749
rect 7929 6749 7941 6783
rect 7975 6749 7987 6783
rect 9674 6780 9680 6792
rect 7929 6743 7987 6749
rect 8036 6752 9680 6780
rect 5261 6715 5319 6721
rect 5261 6681 5273 6715
rect 5307 6712 5319 6715
rect 5307 6684 7696 6712
rect 5307 6681 5319 6684
rect 5261 6675 5319 6681
rect 6086 6644 6092 6656
rect 6047 6616 6092 6644
rect 6086 6604 6092 6616
rect 6144 6604 6150 6656
rect 6454 6644 6460 6656
rect 6415 6616 6460 6644
rect 6454 6604 6460 6616
rect 6512 6604 6518 6656
rect 6546 6604 6552 6656
rect 6604 6644 6610 6656
rect 7668 6644 7696 6684
rect 7742 6672 7748 6724
rect 7800 6712 7806 6724
rect 7944 6712 7972 6743
rect 7800 6684 7972 6712
rect 7800 6672 7806 6684
rect 8036 6644 8064 6752
rect 9674 6740 9680 6752
rect 9732 6780 9738 6792
rect 10226 6780 10232 6792
rect 9732 6752 10232 6780
rect 9732 6740 9738 6752
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 10594 6740 10600 6792
rect 10652 6789 10658 6792
rect 10652 6780 10664 6789
rect 10652 6752 10697 6780
rect 10652 6743 10664 6752
rect 10652 6740 10658 6743
rect 11698 6740 11704 6792
rect 11756 6780 11762 6792
rect 12820 6780 12848 6811
rect 13998 6808 14004 6820
rect 14056 6808 14062 6860
rect 17126 6848 17132 6860
rect 17039 6820 17132 6848
rect 17126 6808 17132 6820
rect 17184 6848 17190 6860
rect 17184 6820 22784 6848
rect 17184 6808 17190 6820
rect 11756 6752 12848 6780
rect 11756 6740 11762 6752
rect 13078 6740 13084 6792
rect 13136 6780 13142 6792
rect 16853 6783 16911 6789
rect 16853 6780 16865 6783
rect 13136 6752 16865 6780
rect 13136 6740 13142 6752
rect 16853 6749 16865 6752
rect 16899 6749 16911 6783
rect 19426 6780 19432 6792
rect 19387 6752 19432 6780
rect 16853 6743 16911 6749
rect 11790 6712 11796 6724
rect 8128 6684 11796 6712
rect 8128 6653 8156 6684
rect 11790 6672 11796 6684
rect 11848 6672 11854 6724
rect 6604 6616 6649 6644
rect 7668 6616 8064 6644
rect 8113 6647 8171 6653
rect 6604 6604 6610 6616
rect 8113 6613 8125 6647
rect 8159 6613 8171 6647
rect 9490 6644 9496 6656
rect 9451 6616 9496 6644
rect 8113 6607 8171 6613
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 12250 6644 12256 6656
rect 12211 6616 12256 6644
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 12618 6644 12624 6656
rect 12579 6616 12624 6644
rect 12618 6604 12624 6616
rect 12676 6604 12682 6656
rect 12710 6604 12716 6656
rect 12768 6644 12774 6656
rect 16868 6644 16896 6743
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 19613 6783 19671 6789
rect 19613 6749 19625 6783
rect 19659 6780 19671 6783
rect 20714 6780 20720 6792
rect 19659 6752 20720 6780
rect 19659 6749 19671 6752
rect 19613 6743 19671 6749
rect 20714 6740 20720 6752
rect 20772 6780 20778 6792
rect 21634 6780 21640 6792
rect 20772 6752 21640 6780
rect 20772 6740 20778 6752
rect 21634 6740 21640 6752
rect 21692 6740 21698 6792
rect 22646 6780 22652 6792
rect 22607 6752 22652 6780
rect 22646 6740 22652 6752
rect 22704 6740 22710 6792
rect 22756 6780 22784 6820
rect 22905 6783 22963 6789
rect 22905 6780 22917 6783
rect 22756 6752 22917 6780
rect 22905 6749 22917 6752
rect 22951 6749 22963 6783
rect 22905 6743 22963 6749
rect 25685 6783 25743 6789
rect 25685 6749 25697 6783
rect 25731 6749 25743 6783
rect 25685 6743 25743 6749
rect 25777 6783 25835 6789
rect 25777 6749 25789 6783
rect 25823 6780 25835 6783
rect 26329 6783 26387 6789
rect 26329 6780 26341 6783
rect 25823 6752 26341 6780
rect 25823 6749 25835 6752
rect 25777 6743 25835 6749
rect 26329 6749 26341 6752
rect 26375 6749 26387 6783
rect 26329 6743 26387 6749
rect 26596 6783 26654 6789
rect 26596 6749 26608 6783
rect 26642 6780 26654 6783
rect 28074 6780 28080 6792
rect 26642 6752 28080 6780
rect 26642 6749 26654 6752
rect 26596 6743 26654 6749
rect 17586 6672 17592 6724
rect 17644 6672 17650 6724
rect 25700 6712 25728 6743
rect 28074 6740 28080 6752
rect 28132 6740 28138 6792
rect 26418 6712 26424 6724
rect 25700 6684 26424 6712
rect 26418 6672 26424 6684
rect 26476 6672 26482 6724
rect 18138 6644 18144 6656
rect 12768 6616 12813 6644
rect 16868 6616 18144 6644
rect 12768 6604 12774 6616
rect 18138 6604 18144 6616
rect 18196 6604 18202 6656
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 18601 6647 18659 6653
rect 18601 6644 18613 6647
rect 18564 6616 18613 6644
rect 18564 6604 18570 6616
rect 18601 6613 18613 6616
rect 18647 6613 18659 6647
rect 19518 6644 19524 6656
rect 19479 6616 19524 6644
rect 18601 6607 18659 6613
rect 19518 6604 19524 6616
rect 19576 6604 19582 6656
rect 24029 6647 24087 6653
rect 24029 6613 24041 6647
rect 24075 6644 24087 6647
rect 26602 6644 26608 6656
rect 24075 6616 26608 6644
rect 24075 6613 24087 6616
rect 24029 6607 24087 6613
rect 26602 6604 26608 6616
rect 26660 6604 26666 6656
rect 1104 6554 29048 6576
rect 1104 6502 7896 6554
rect 7948 6502 7960 6554
rect 8012 6502 8024 6554
rect 8076 6502 8088 6554
rect 8140 6502 8152 6554
rect 8204 6502 14842 6554
rect 14894 6502 14906 6554
rect 14958 6502 14970 6554
rect 15022 6502 15034 6554
rect 15086 6502 15098 6554
rect 15150 6502 21788 6554
rect 21840 6502 21852 6554
rect 21904 6502 21916 6554
rect 21968 6502 21980 6554
rect 22032 6502 22044 6554
rect 22096 6502 28734 6554
rect 28786 6502 28798 6554
rect 28850 6502 28862 6554
rect 28914 6502 28926 6554
rect 28978 6502 28990 6554
rect 29042 6502 29048 6554
rect 1104 6480 29048 6502
rect 2130 6400 2136 6452
rect 2188 6440 2194 6452
rect 2593 6443 2651 6449
rect 2593 6440 2605 6443
rect 2188 6412 2605 6440
rect 2188 6400 2194 6412
rect 2593 6409 2605 6412
rect 2639 6409 2651 6443
rect 2593 6403 2651 6409
rect 6454 6400 6460 6452
rect 6512 6440 6518 6452
rect 12618 6440 12624 6452
rect 6512 6412 12624 6440
rect 6512 6400 6518 6412
rect 12618 6400 12624 6412
rect 12676 6400 12682 6452
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 13265 6443 13323 6449
rect 13265 6440 13277 6443
rect 12768 6412 13277 6440
rect 12768 6400 12774 6412
rect 13265 6409 13277 6412
rect 13311 6409 13323 6443
rect 17586 6440 17592 6452
rect 17547 6412 17592 6440
rect 13265 6403 13323 6409
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 19426 6440 19432 6452
rect 17696 6412 19432 6440
rect 6546 6332 6552 6384
rect 6604 6372 6610 6384
rect 6641 6375 6699 6381
rect 6641 6372 6653 6375
rect 6604 6344 6653 6372
rect 6604 6332 6610 6344
rect 6641 6341 6653 6344
rect 6687 6341 6699 6375
rect 6641 6335 6699 6341
rect 12152 6375 12210 6381
rect 12152 6341 12164 6375
rect 12198 6372 12210 6375
rect 12250 6372 12256 6384
rect 12198 6344 12256 6372
rect 12198 6341 12210 6344
rect 12152 6335 12210 6341
rect 12250 6332 12256 6344
rect 12308 6332 12314 6384
rect 17696 6372 17724 6412
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 24305 6443 24363 6449
rect 24305 6409 24317 6443
rect 24351 6440 24363 6443
rect 25038 6440 25044 6452
rect 24351 6412 25044 6440
rect 24351 6409 24363 6412
rect 24305 6403 24363 6409
rect 25038 6400 25044 6412
rect 25096 6400 25102 6452
rect 17512 6344 17724 6372
rect 2590 6264 2596 6316
rect 2648 6304 2654 6316
rect 2685 6307 2743 6313
rect 2685 6304 2697 6307
rect 2648 6276 2697 6304
rect 2648 6264 2654 6276
rect 2685 6273 2697 6276
rect 2731 6304 2743 6307
rect 3145 6307 3203 6313
rect 3145 6304 3157 6307
rect 2731 6276 3157 6304
rect 2731 6273 2743 6276
rect 2685 6267 2743 6273
rect 3145 6273 3157 6276
rect 3191 6304 3203 6307
rect 5077 6307 5135 6313
rect 5077 6304 5089 6307
rect 3191 6276 5089 6304
rect 3191 6273 3203 6276
rect 3145 6267 3203 6273
rect 5077 6273 5089 6276
rect 5123 6273 5135 6307
rect 6822 6304 6828 6316
rect 6783 6276 6828 6304
rect 5077 6267 5135 6273
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 7098 6264 7104 6316
rect 7156 6304 7162 6316
rect 7653 6307 7711 6313
rect 7653 6304 7665 6307
rect 7156 6276 7665 6304
rect 7156 6264 7162 6276
rect 7653 6273 7665 6276
rect 7699 6273 7711 6307
rect 9490 6304 9496 6316
rect 7653 6267 7711 6273
rect 7760 6276 9496 6304
rect 5169 6239 5227 6245
rect 5169 6205 5181 6239
rect 5215 6236 5227 6239
rect 5810 6236 5816 6248
rect 5215 6208 5816 6236
rect 5215 6205 5227 6208
rect 5169 6199 5227 6205
rect 5810 6196 5816 6208
rect 5868 6196 5874 6248
rect 7760 6245 7788 6276
rect 9490 6264 9496 6276
rect 9548 6264 9554 6316
rect 9950 6264 9956 6316
rect 10008 6304 10014 6316
rect 10514 6307 10572 6313
rect 10514 6304 10526 6307
rect 10008 6276 10526 6304
rect 10008 6264 10014 6276
rect 10514 6273 10526 6276
rect 10560 6273 10572 6307
rect 10514 6267 10572 6273
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6304 10839 6307
rect 10870 6304 10876 6316
rect 10827 6276 10876 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 10870 6264 10876 6276
rect 10928 6304 10934 6316
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 10928 6276 11897 6304
rect 10928 6264 10934 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 17034 6264 17040 6316
rect 17092 6304 17098 6316
rect 17512 6313 17540 6344
rect 19518 6332 19524 6384
rect 19576 6332 19582 6384
rect 17497 6307 17555 6313
rect 17497 6304 17509 6307
rect 17092 6276 17509 6304
rect 17092 6264 17098 6276
rect 17497 6273 17509 6276
rect 17543 6273 17555 6307
rect 17497 6267 17555 6273
rect 17681 6307 17739 6313
rect 17681 6273 17693 6307
rect 17727 6273 17739 6307
rect 18506 6304 18512 6316
rect 18467 6276 18512 6304
rect 17681 6267 17739 6273
rect 7745 6239 7803 6245
rect 7745 6205 7757 6239
rect 7791 6205 7803 6239
rect 7745 6199 7803 6205
rect 8021 6239 8079 6245
rect 8021 6205 8033 6239
rect 8067 6236 8079 6239
rect 9582 6236 9588 6248
rect 8067 6208 9588 6236
rect 8067 6205 8079 6208
rect 8021 6199 8079 6205
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 16850 6196 16856 6248
rect 16908 6236 16914 6248
rect 17696 6236 17724 6267
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 19426 6264 19432 6316
rect 19484 6304 19490 6316
rect 20441 6307 20499 6313
rect 20441 6304 20453 6307
rect 19484 6276 20453 6304
rect 19484 6264 19490 6276
rect 20441 6273 20453 6276
rect 20487 6273 20499 6307
rect 20441 6267 20499 6273
rect 20625 6307 20683 6313
rect 20625 6273 20637 6307
rect 20671 6304 20683 6307
rect 20714 6304 20720 6316
rect 20671 6276 20720 6304
rect 20671 6273 20683 6276
rect 20625 6267 20683 6273
rect 18138 6236 18144 6248
rect 16908 6208 17724 6236
rect 18051 6208 18144 6236
rect 16908 6196 16914 6208
rect 18138 6196 18144 6208
rect 18196 6236 18202 6248
rect 19518 6236 19524 6248
rect 18196 6208 19524 6236
rect 18196 6196 18202 6208
rect 19518 6196 19524 6208
rect 19576 6196 19582 6248
rect 20456 6236 20484 6267
rect 20714 6264 20720 6276
rect 20772 6264 20778 6316
rect 21266 6264 21272 6316
rect 21324 6304 21330 6316
rect 23181 6307 23239 6313
rect 23181 6304 23193 6307
rect 21324 6276 23193 6304
rect 21324 6264 21330 6276
rect 23181 6273 23193 6276
rect 23227 6273 23239 6307
rect 27890 6304 27896 6316
rect 27851 6276 27896 6304
rect 23181 6267 23239 6273
rect 27890 6264 27896 6276
rect 27948 6264 27954 6316
rect 20456 6208 22094 6236
rect 5445 6171 5503 6177
rect 5445 6137 5457 6171
rect 5491 6168 5503 6171
rect 6730 6168 6736 6180
rect 5491 6140 6736 6168
rect 5491 6137 5503 6140
rect 5445 6131 5503 6137
rect 6730 6128 6736 6140
rect 6788 6128 6794 6180
rect 22066 6112 22094 6208
rect 22646 6196 22652 6248
rect 22704 6236 22710 6248
rect 22925 6239 22983 6245
rect 22925 6236 22937 6239
rect 22704 6208 22937 6236
rect 22704 6196 22710 6208
rect 22925 6205 22937 6208
rect 22971 6205 22983 6239
rect 28166 6236 28172 6248
rect 28127 6208 28172 6236
rect 22925 6199 22983 6205
rect 28166 6196 28172 6208
rect 28224 6196 28230 6248
rect 3237 6103 3295 6109
rect 3237 6069 3249 6103
rect 3283 6100 3295 6103
rect 4062 6100 4068 6112
rect 3283 6072 4068 6100
rect 3283 6069 3295 6072
rect 3237 6063 3295 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 7009 6103 7067 6109
rect 7009 6069 7021 6103
rect 7055 6100 7067 6103
rect 7650 6100 7656 6112
rect 7055 6072 7656 6100
rect 7055 6069 7067 6072
rect 7009 6063 7067 6069
rect 7650 6060 7656 6072
rect 7708 6060 7714 6112
rect 8478 6060 8484 6112
rect 8536 6100 8542 6112
rect 9401 6103 9459 6109
rect 9401 6100 9413 6103
rect 8536 6072 9413 6100
rect 8536 6060 8542 6072
rect 9401 6069 9413 6072
rect 9447 6069 9459 6103
rect 9401 6063 9459 6069
rect 19794 6060 19800 6112
rect 19852 6100 19858 6112
rect 19935 6103 19993 6109
rect 19935 6100 19947 6103
rect 19852 6072 19947 6100
rect 19852 6060 19858 6072
rect 19935 6069 19947 6072
rect 19981 6069 19993 6103
rect 20530 6100 20536 6112
rect 20491 6072 20536 6100
rect 19935 6063 19993 6069
rect 20530 6060 20536 6072
rect 20588 6060 20594 6112
rect 22066 6072 22100 6112
rect 22094 6060 22100 6072
rect 22152 6100 22158 6112
rect 24762 6100 24768 6112
rect 22152 6072 24768 6100
rect 22152 6060 22158 6072
rect 24762 6060 24768 6072
rect 24820 6060 24826 6112
rect 1104 6010 28888 6032
rect 1104 5958 4423 6010
rect 4475 5958 4487 6010
rect 4539 5958 4551 6010
rect 4603 5958 4615 6010
rect 4667 5958 4679 6010
rect 4731 5958 11369 6010
rect 11421 5958 11433 6010
rect 11485 5958 11497 6010
rect 11549 5958 11561 6010
rect 11613 5958 11625 6010
rect 11677 5958 18315 6010
rect 18367 5958 18379 6010
rect 18431 5958 18443 6010
rect 18495 5958 18507 6010
rect 18559 5958 18571 6010
rect 18623 5958 25261 6010
rect 25313 5958 25325 6010
rect 25377 5958 25389 6010
rect 25441 5958 25453 6010
rect 25505 5958 25517 6010
rect 25569 5958 28888 6010
rect 1104 5936 28888 5958
rect 4798 5856 4804 5908
rect 4856 5896 4862 5908
rect 4856 5868 6408 5896
rect 4856 5856 4862 5868
rect 6380 5828 6408 5868
rect 6546 5856 6552 5908
rect 6604 5896 6610 5908
rect 6825 5899 6883 5905
rect 6825 5896 6837 5899
rect 6604 5868 6837 5896
rect 6604 5856 6610 5868
rect 6825 5865 6837 5868
rect 6871 5865 6883 5899
rect 6825 5859 6883 5865
rect 7742 5856 7748 5908
rect 7800 5896 7806 5908
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 7800 5868 7849 5896
rect 7800 5856 7806 5868
rect 7837 5865 7849 5868
rect 7883 5865 7895 5899
rect 7837 5859 7895 5865
rect 9861 5899 9919 5905
rect 9861 5865 9873 5899
rect 9907 5896 9919 5899
rect 9950 5896 9956 5908
rect 9907 5868 9956 5896
rect 9907 5865 9919 5868
rect 9861 5859 9919 5865
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 10686 5856 10692 5908
rect 10744 5896 10750 5908
rect 11793 5899 11851 5905
rect 11793 5896 11805 5899
rect 10744 5868 11805 5896
rect 10744 5856 10750 5868
rect 11793 5865 11805 5868
rect 11839 5865 11851 5899
rect 11793 5859 11851 5865
rect 13906 5856 13912 5908
rect 13964 5896 13970 5908
rect 15102 5896 15108 5908
rect 13964 5868 15108 5896
rect 13964 5856 13970 5868
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 17126 5856 17132 5908
rect 17184 5905 17190 5908
rect 17184 5899 17233 5905
rect 17184 5865 17187 5899
rect 17221 5865 17233 5899
rect 21266 5896 21272 5908
rect 21227 5868 21272 5896
rect 17184 5859 17233 5865
rect 17184 5856 17190 5859
rect 21266 5856 21272 5868
rect 21324 5856 21330 5908
rect 6380 5800 12848 5828
rect 4982 5720 4988 5772
rect 5040 5760 5046 5772
rect 5445 5763 5503 5769
rect 5445 5760 5457 5763
rect 5040 5732 5457 5760
rect 5040 5720 5046 5732
rect 5445 5729 5457 5732
rect 5491 5729 5503 5763
rect 10502 5760 10508 5772
rect 10463 5732 10508 5760
rect 5445 5723 5503 5729
rect 10502 5720 10508 5732
rect 10560 5720 10566 5772
rect 12253 5763 12311 5769
rect 12253 5729 12265 5763
rect 12299 5760 12311 5763
rect 12710 5760 12716 5772
rect 12299 5732 12716 5760
rect 12299 5729 12311 5732
rect 12253 5723 12311 5729
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 2498 5652 2504 5704
rect 2556 5692 2562 5704
rect 2593 5695 2651 5701
rect 2593 5692 2605 5695
rect 2556 5664 2605 5692
rect 2556 5652 2562 5664
rect 2593 5661 2605 5664
rect 2639 5661 2651 5695
rect 2593 5655 2651 5661
rect 3053 5695 3111 5701
rect 3053 5661 3065 5695
rect 3099 5661 3111 5695
rect 3053 5655 3111 5661
rect 3068 5624 3096 5655
rect 3326 5652 3332 5704
rect 3384 5692 3390 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3384 5664 3985 5692
rect 3384 5652 3390 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 5712 5695 5770 5701
rect 5712 5661 5724 5695
rect 5758 5692 5770 5695
rect 6086 5692 6092 5704
rect 5758 5664 6092 5692
rect 5758 5661 5770 5664
rect 5712 5655 5770 5661
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 7282 5692 7288 5704
rect 7243 5664 7288 5692
rect 7282 5652 7288 5664
rect 7340 5652 7346 5704
rect 7650 5692 7656 5704
rect 7611 5664 7656 5692
rect 7650 5652 7656 5664
rect 7708 5652 7714 5704
rect 8294 5692 8300 5704
rect 8255 5664 8300 5692
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 8478 5692 8484 5704
rect 8439 5664 8484 5692
rect 8478 5652 8484 5664
rect 8536 5692 8542 5704
rect 10321 5695 10379 5701
rect 10321 5692 10333 5695
rect 8536 5664 10333 5692
rect 8536 5652 8542 5664
rect 10321 5661 10333 5664
rect 10367 5661 10379 5695
rect 12158 5692 12164 5704
rect 12119 5664 12164 5692
rect 10321 5655 10379 5661
rect 12158 5652 12164 5664
rect 12216 5652 12222 5704
rect 12820 5692 12848 5800
rect 14476 5800 15056 5828
rect 14476 5692 14504 5800
rect 14550 5720 14556 5772
rect 14608 5760 14614 5772
rect 15028 5760 15056 5800
rect 17034 5760 17040 5772
rect 14608 5732 14964 5760
rect 15028 5732 17040 5760
rect 14608 5720 14614 5732
rect 14936 5701 14964 5732
rect 17034 5720 17040 5732
rect 17092 5720 17098 5772
rect 19794 5760 19800 5772
rect 19755 5732 19800 5760
rect 19794 5720 19800 5732
rect 19852 5720 19858 5772
rect 14737 5695 14795 5701
rect 14737 5692 14749 5695
rect 12820 5664 14749 5692
rect 14737 5661 14749 5664
rect 14783 5661 14795 5695
rect 14737 5655 14795 5661
rect 14921 5695 14979 5701
rect 14921 5661 14933 5695
rect 14967 5661 14979 5695
rect 14921 5655 14979 5661
rect 4154 5624 4160 5636
rect 3068 5596 4160 5624
rect 4154 5584 4160 5596
rect 4212 5584 4218 5636
rect 7469 5627 7527 5633
rect 7469 5593 7481 5627
rect 7515 5593 7527 5627
rect 7469 5587 7527 5593
rect 3418 5556 3424 5568
rect 3379 5528 3424 5556
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 4065 5559 4123 5565
rect 4065 5525 4077 5559
rect 4111 5556 4123 5559
rect 4338 5556 4344 5568
rect 4111 5528 4344 5556
rect 4111 5525 4123 5528
rect 4065 5519 4123 5525
rect 4338 5516 4344 5528
rect 4396 5516 4402 5568
rect 7484 5556 7512 5587
rect 7558 5584 7564 5636
rect 7616 5624 7622 5636
rect 10226 5624 10232 5636
rect 7616 5596 7661 5624
rect 10187 5596 10232 5624
rect 7616 5584 7622 5596
rect 10226 5584 10232 5596
rect 10284 5584 10290 5636
rect 14936 5624 14964 5655
rect 15102 5652 15108 5704
rect 15160 5692 15166 5704
rect 15381 5695 15439 5701
rect 15381 5692 15393 5695
rect 15160 5664 15393 5692
rect 15160 5652 15166 5664
rect 15381 5661 15393 5664
rect 15427 5661 15439 5695
rect 15746 5692 15752 5704
rect 15707 5664 15752 5692
rect 15381 5655 15439 5661
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 19518 5692 19524 5704
rect 19479 5664 19524 5692
rect 19518 5652 19524 5664
rect 19576 5652 19582 5704
rect 21634 5652 21640 5704
rect 21692 5692 21698 5704
rect 21729 5695 21787 5701
rect 21729 5692 21741 5695
rect 21692 5664 21741 5692
rect 21692 5652 21698 5664
rect 21729 5661 21741 5664
rect 21775 5661 21787 5695
rect 21729 5655 21787 5661
rect 21913 5695 21971 5701
rect 21913 5661 21925 5695
rect 21959 5692 21971 5695
rect 22094 5692 22100 5704
rect 21959 5664 22100 5692
rect 21959 5661 21971 5664
rect 21913 5655 21971 5661
rect 22094 5652 22100 5664
rect 22152 5652 22158 5704
rect 27798 5692 27804 5704
rect 27759 5664 27804 5692
rect 27798 5652 27804 5664
rect 27856 5652 27862 5704
rect 14936 5596 15424 5624
rect 8297 5559 8355 5565
rect 8297 5556 8309 5559
rect 7484 5528 8309 5556
rect 8297 5525 8309 5528
rect 8343 5525 8355 5559
rect 8297 5519 8355 5525
rect 14921 5559 14979 5565
rect 14921 5525 14933 5559
rect 14967 5556 14979 5559
rect 15286 5556 15292 5568
rect 14967 5528 15292 5556
rect 14967 5525 14979 5528
rect 14921 5519 14979 5525
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 15396 5556 15424 5596
rect 16758 5584 16764 5636
rect 16816 5584 16822 5636
rect 20530 5584 20536 5636
rect 20588 5584 20594 5636
rect 27246 5584 27252 5636
rect 27304 5624 27310 5636
rect 27534 5627 27592 5633
rect 27534 5624 27546 5627
rect 27304 5596 27546 5624
rect 27304 5584 27310 5596
rect 27534 5593 27546 5596
rect 27580 5593 27592 5627
rect 27534 5587 27592 5593
rect 16942 5556 16948 5568
rect 15396 5528 16948 5556
rect 16942 5516 16948 5528
rect 17000 5516 17006 5568
rect 21634 5516 21640 5568
rect 21692 5556 21698 5568
rect 21729 5559 21787 5565
rect 21729 5556 21741 5559
rect 21692 5528 21741 5556
rect 21692 5516 21698 5528
rect 21729 5525 21741 5528
rect 21775 5525 21787 5559
rect 26418 5556 26424 5568
rect 26379 5528 26424 5556
rect 21729 5519 21787 5525
rect 26418 5516 26424 5528
rect 26476 5516 26482 5568
rect 1104 5466 29048 5488
rect 1104 5414 7896 5466
rect 7948 5414 7960 5466
rect 8012 5414 8024 5466
rect 8076 5414 8088 5466
rect 8140 5414 8152 5466
rect 8204 5414 14842 5466
rect 14894 5414 14906 5466
rect 14958 5414 14970 5466
rect 15022 5414 15034 5466
rect 15086 5414 15098 5466
rect 15150 5414 21788 5466
rect 21840 5414 21852 5466
rect 21904 5414 21916 5466
rect 21968 5414 21980 5466
rect 22032 5414 22044 5466
rect 22096 5414 28734 5466
rect 28786 5414 28798 5466
rect 28850 5414 28862 5466
rect 28914 5414 28926 5466
rect 28978 5414 28990 5466
rect 29042 5414 29048 5466
rect 1104 5392 29048 5414
rect 2590 5352 2596 5364
rect 2551 5324 2596 5352
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 7282 5312 7288 5364
rect 7340 5352 7346 5364
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 7340 5324 7389 5352
rect 7340 5312 7346 5324
rect 7377 5321 7389 5324
rect 7423 5321 7435 5355
rect 7377 5315 7435 5321
rect 7558 5312 7564 5364
rect 7616 5312 7622 5364
rect 15746 5352 15752 5364
rect 15707 5324 15752 5352
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 16758 5312 16764 5364
rect 16816 5352 16822 5364
rect 16853 5355 16911 5361
rect 16853 5352 16865 5355
rect 16816 5324 16865 5352
rect 16816 5312 16822 5324
rect 16853 5321 16865 5324
rect 16899 5321 16911 5355
rect 16853 5315 16911 5321
rect 25682 5312 25688 5364
rect 25740 5352 25746 5364
rect 26145 5355 26203 5361
rect 26145 5352 26157 5355
rect 25740 5324 26157 5352
rect 25740 5312 25746 5324
rect 26145 5321 26157 5324
rect 26191 5321 26203 5355
rect 27246 5352 27252 5364
rect 27207 5324 27252 5352
rect 26145 5315 26203 5321
rect 27246 5312 27252 5324
rect 27304 5312 27310 5364
rect 27798 5312 27804 5364
rect 27856 5352 27862 5364
rect 27893 5355 27951 5361
rect 27893 5352 27905 5355
rect 27856 5324 27905 5352
rect 27856 5312 27862 5324
rect 27893 5321 27905 5324
rect 27939 5321 27951 5355
rect 27893 5315 27951 5321
rect 3418 5244 3424 5296
rect 3476 5244 3482 5296
rect 4062 5284 4068 5296
rect 4023 5256 4068 5284
rect 4062 5244 4068 5256
rect 4120 5244 4126 5296
rect 6825 5287 6883 5293
rect 6825 5253 6837 5287
rect 6871 5284 6883 5287
rect 7576 5284 7604 5312
rect 6871 5256 7604 5284
rect 7745 5287 7803 5293
rect 6871 5253 6883 5256
rect 6825 5247 6883 5253
rect 7745 5253 7757 5287
rect 7791 5284 7803 5287
rect 8478 5284 8484 5296
rect 7791 5256 8484 5284
rect 7791 5253 7803 5256
rect 7745 5247 7803 5253
rect 8478 5244 8484 5256
rect 8536 5244 8542 5296
rect 15286 5244 15292 5296
rect 15344 5244 15350 5296
rect 22020 5256 22876 5284
rect 4338 5176 4344 5228
rect 4396 5216 4402 5228
rect 4396 5188 4441 5216
rect 4396 5176 4402 5188
rect 6546 5176 6552 5228
rect 6604 5216 6610 5228
rect 6733 5219 6791 5225
rect 6733 5216 6745 5219
rect 6604 5188 6745 5216
rect 6604 5176 6610 5188
rect 6733 5185 6745 5188
rect 6779 5185 6791 5219
rect 6733 5179 6791 5185
rect 6917 5219 6975 5225
rect 6917 5185 6929 5219
rect 6963 5185 6975 5219
rect 6917 5179 6975 5185
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 8294 5216 8300 5228
rect 7607 5188 8300 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 5534 5108 5540 5160
rect 5592 5148 5598 5160
rect 6822 5148 6828 5160
rect 5592 5120 6828 5148
rect 5592 5108 5598 5120
rect 6822 5108 6828 5120
rect 6880 5148 6886 5160
rect 6932 5148 6960 5179
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 16850 5216 16856 5228
rect 16811 5188 16856 5216
rect 16850 5176 16856 5188
rect 16908 5176 16914 5228
rect 17034 5216 17040 5228
rect 16995 5188 17040 5216
rect 17034 5176 17040 5188
rect 17092 5176 17098 5228
rect 21542 5176 21548 5228
rect 21600 5216 21606 5228
rect 22020 5225 22048 5256
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 21600 5188 22017 5216
rect 21600 5176 21606 5188
rect 22005 5185 22017 5188
rect 22051 5185 22063 5219
rect 22186 5216 22192 5228
rect 22147 5188 22192 5216
rect 22005 5179 22063 5185
rect 22186 5176 22192 5188
rect 22244 5216 22250 5228
rect 22848 5225 22876 5256
rect 26418 5244 26424 5296
rect 26476 5284 26482 5296
rect 26476 5256 27200 5284
rect 26476 5244 26482 5256
rect 22649 5219 22707 5225
rect 22649 5216 22661 5219
rect 22244 5188 22661 5216
rect 22244 5176 22250 5188
rect 22649 5185 22661 5188
rect 22695 5185 22707 5219
rect 22649 5179 22707 5185
rect 22833 5219 22891 5225
rect 22833 5185 22845 5219
rect 22879 5185 22891 5219
rect 22833 5179 22891 5185
rect 26142 5176 26148 5228
rect 26200 5216 26206 5228
rect 26237 5219 26295 5225
rect 26237 5216 26249 5219
rect 26200 5188 26249 5216
rect 26200 5176 26206 5188
rect 26237 5185 26249 5188
rect 26283 5185 26295 5219
rect 26237 5179 26295 5185
rect 26326 5176 26332 5228
rect 26384 5216 26390 5228
rect 27172 5225 27200 5256
rect 27157 5219 27215 5225
rect 26384 5188 26429 5216
rect 26384 5176 26390 5188
rect 27157 5185 27169 5219
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 27522 5176 27528 5228
rect 27580 5216 27586 5228
rect 27801 5219 27859 5225
rect 27801 5216 27813 5219
rect 27580 5188 27813 5216
rect 27580 5176 27586 5188
rect 27801 5185 27813 5188
rect 27847 5185 27859 5219
rect 27801 5179 27859 5185
rect 6880 5120 6960 5148
rect 6880 5108 6886 5120
rect 13906 5108 13912 5160
rect 13964 5148 13970 5160
rect 14001 5151 14059 5157
rect 14001 5148 14013 5151
rect 13964 5120 14013 5148
rect 13964 5108 13970 5120
rect 14001 5117 14013 5120
rect 14047 5117 14059 5151
rect 14274 5148 14280 5160
rect 14235 5120 14280 5148
rect 14001 5111 14059 5117
rect 14274 5108 14280 5120
rect 14332 5108 14338 5160
rect 25958 5148 25964 5160
rect 25919 5120 25964 5148
rect 25958 5108 25964 5120
rect 26016 5108 26022 5160
rect 22097 5015 22155 5021
rect 22097 4981 22109 5015
rect 22143 5012 22155 5015
rect 22278 5012 22284 5024
rect 22143 4984 22284 5012
rect 22143 4981 22155 4984
rect 22097 4975 22155 4981
rect 22278 4972 22284 4984
rect 22336 4972 22342 5024
rect 22738 5012 22744 5024
rect 22699 4984 22744 5012
rect 22738 4972 22744 4984
rect 22796 4972 22802 5024
rect 26237 5015 26295 5021
rect 26237 4981 26249 5015
rect 26283 5012 26295 5015
rect 26694 5012 26700 5024
rect 26283 4984 26700 5012
rect 26283 4981 26295 4984
rect 26237 4975 26295 4981
rect 26694 4972 26700 4984
rect 26752 4972 26758 5024
rect 1104 4922 28888 4944
rect 1104 4870 4423 4922
rect 4475 4870 4487 4922
rect 4539 4870 4551 4922
rect 4603 4870 4615 4922
rect 4667 4870 4679 4922
rect 4731 4870 11369 4922
rect 11421 4870 11433 4922
rect 11485 4870 11497 4922
rect 11549 4870 11561 4922
rect 11613 4870 11625 4922
rect 11677 4870 18315 4922
rect 18367 4870 18379 4922
rect 18431 4870 18443 4922
rect 18495 4870 18507 4922
rect 18559 4870 18571 4922
rect 18623 4870 25261 4922
rect 25313 4870 25325 4922
rect 25377 4870 25389 4922
rect 25441 4870 25453 4922
rect 25505 4870 25517 4922
rect 25569 4870 28888 4922
rect 1104 4848 28888 4870
rect 24029 4811 24087 4817
rect 24029 4777 24041 4811
rect 24075 4808 24087 4811
rect 26326 4808 26332 4820
rect 24075 4780 26332 4808
rect 24075 4777 24087 4780
rect 24029 4771 24087 4777
rect 26326 4768 26332 4780
rect 26384 4808 26390 4820
rect 27246 4808 27252 4820
rect 26384 4780 27252 4808
rect 26384 4768 26390 4780
rect 27246 4768 27252 4780
rect 27304 4768 27310 4820
rect 27341 4811 27399 4817
rect 27341 4777 27353 4811
rect 27387 4808 27399 4811
rect 27430 4808 27436 4820
rect 27387 4780 27436 4808
rect 27387 4777 27399 4780
rect 27341 4771 27399 4777
rect 27430 4768 27436 4780
rect 27488 4768 27494 4820
rect 27890 4808 27896 4820
rect 27851 4780 27896 4808
rect 27890 4768 27896 4780
rect 27948 4768 27954 4820
rect 4154 4632 4160 4684
rect 4212 4672 4218 4684
rect 6457 4675 6515 4681
rect 6457 4672 6469 4675
rect 4212 4644 6469 4672
rect 4212 4632 4218 4644
rect 6457 4641 6469 4644
rect 6503 4672 6515 4675
rect 6822 4672 6828 4684
rect 6503 4644 6828 4672
rect 6503 4641 6515 4644
rect 6457 4635 6515 4641
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 11054 4672 11060 4684
rect 9968 4644 11060 4672
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4573 4767 4607
rect 6730 4604 6736 4616
rect 6691 4576 6736 4604
rect 4709 4567 4767 4573
rect 4724 4536 4752 4567
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4604 7895 4607
rect 8294 4604 8300 4616
rect 7883 4576 8300 4604
rect 7883 4573 7895 4576
rect 7837 4567 7895 4573
rect 8294 4564 8300 4576
rect 8352 4604 8358 4616
rect 9968 4613 9996 4644
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 20717 4675 20775 4681
rect 20717 4641 20729 4675
rect 20763 4672 20775 4675
rect 21266 4672 21272 4684
rect 20763 4644 21272 4672
rect 20763 4641 20775 4644
rect 20717 4635 20775 4641
rect 21266 4632 21272 4644
rect 21324 4632 21330 4684
rect 28258 4672 28264 4684
rect 28219 4644 28264 4672
rect 28258 4632 28264 4644
rect 28316 4632 28322 4684
rect 9953 4607 10011 4613
rect 9953 4604 9965 4607
rect 8352 4576 9965 4604
rect 8352 4564 8358 4576
rect 9953 4573 9965 4576
rect 9999 4573 10011 4607
rect 9953 4567 10011 4573
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4573 10563 4607
rect 10686 4604 10692 4616
rect 10647 4576 10692 4604
rect 10505 4567 10563 4573
rect 6638 4536 6644 4548
rect 4724 4508 6644 4536
rect 6638 4496 6644 4508
rect 6696 4496 6702 4548
rect 9766 4496 9772 4548
rect 9824 4536 9830 4548
rect 10520 4536 10548 4567
rect 10686 4564 10692 4576
rect 10744 4604 10750 4616
rect 13814 4604 13820 4616
rect 10744 4576 13820 4604
rect 10744 4564 10750 4576
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 19518 4564 19524 4616
rect 19576 4604 19582 4616
rect 20349 4607 20407 4613
rect 20349 4604 20361 4607
rect 19576 4576 20361 4604
rect 19576 4564 19582 4576
rect 20349 4573 20361 4576
rect 20395 4604 20407 4607
rect 20622 4604 20628 4616
rect 20395 4576 20628 4604
rect 20395 4573 20407 4576
rect 20349 4567 20407 4573
rect 20622 4564 20628 4576
rect 20680 4564 20686 4616
rect 22646 4604 22652 4616
rect 22559 4576 22652 4604
rect 22646 4564 22652 4576
rect 22704 4604 22710 4616
rect 23290 4604 23296 4616
rect 22704 4576 23296 4604
rect 22704 4564 22710 4576
rect 23290 4564 23296 4576
rect 23348 4564 23354 4616
rect 25501 4607 25559 4613
rect 25501 4573 25513 4607
rect 25547 4604 25559 4607
rect 25958 4604 25964 4616
rect 25547 4576 25964 4604
rect 25547 4573 25559 4576
rect 25501 4567 25559 4573
rect 25958 4564 25964 4576
rect 26016 4604 26022 4616
rect 26234 4604 26240 4616
rect 26016 4576 26240 4604
rect 26016 4564 26022 4576
rect 26234 4564 26240 4576
rect 26292 4564 26298 4616
rect 27065 4607 27123 4613
rect 27065 4573 27077 4607
rect 27111 4573 27123 4607
rect 27065 4567 27123 4573
rect 27157 4607 27215 4613
rect 27157 4573 27169 4607
rect 27203 4604 27215 4607
rect 27706 4604 27712 4616
rect 27203 4576 27712 4604
rect 27203 4573 27215 4576
rect 27157 4567 27215 4573
rect 9824 4508 10548 4536
rect 9824 4496 9830 4508
rect 10594 4496 10600 4548
rect 10652 4536 10658 4548
rect 13630 4536 13636 4548
rect 10652 4508 13636 4536
rect 10652 4496 10658 4508
rect 13630 4496 13636 4508
rect 13688 4496 13694 4548
rect 21634 4496 21640 4548
rect 21692 4496 21698 4548
rect 22922 4545 22928 4548
rect 22916 4499 22928 4545
rect 22980 4536 22986 4548
rect 22980 4508 23016 4536
rect 22922 4496 22928 4499
rect 22980 4496 22986 4508
rect 25590 4496 25596 4548
rect 25648 4536 25654 4548
rect 25777 4539 25835 4545
rect 25777 4536 25789 4539
rect 25648 4508 25789 4536
rect 25648 4496 25654 4508
rect 25777 4505 25789 4508
rect 25823 4505 25835 4539
rect 25777 4499 25835 4505
rect 26053 4539 26111 4545
rect 26053 4505 26065 4539
rect 26099 4536 26111 4539
rect 27080 4536 27108 4567
rect 27706 4564 27712 4576
rect 27764 4564 27770 4616
rect 28169 4607 28227 4613
rect 28169 4573 28181 4607
rect 28215 4573 28227 4607
rect 28169 4567 28227 4573
rect 27430 4536 27436 4548
rect 26099 4508 27436 4536
rect 26099 4505 26111 4508
rect 26053 4499 26111 4505
rect 27430 4496 27436 4508
rect 27488 4536 27494 4548
rect 28184 4536 28212 4567
rect 27488 4508 28212 4536
rect 27488 4496 27494 4508
rect 4338 4428 4344 4480
rect 4396 4468 4402 4480
rect 4617 4471 4675 4477
rect 4617 4468 4629 4471
rect 4396 4440 4629 4468
rect 4396 4428 4402 4440
rect 4617 4437 4629 4440
rect 4663 4437 4675 4471
rect 7374 4468 7380 4480
rect 7335 4440 7380 4468
rect 4617 4431 4675 4437
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 7929 4471 7987 4477
rect 7929 4437 7941 4471
rect 7975 4468 7987 4471
rect 8386 4468 8392 4480
rect 7975 4440 8392 4468
rect 7975 4437 7987 4440
rect 7929 4431 7987 4437
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 9861 4471 9919 4477
rect 9861 4468 9873 4471
rect 9732 4440 9873 4468
rect 9732 4428 9738 4440
rect 9861 4437 9873 4440
rect 9907 4437 9919 4471
rect 9861 4431 9919 4437
rect 11517 4471 11575 4477
rect 11517 4437 11529 4471
rect 11563 4468 11575 4471
rect 11698 4468 11704 4480
rect 11563 4440 11704 4468
rect 11563 4437 11575 4440
rect 11517 4431 11575 4437
rect 11698 4428 11704 4440
rect 11756 4428 11762 4480
rect 22186 4477 22192 4480
rect 22143 4471 22192 4477
rect 22143 4437 22155 4471
rect 22189 4437 22192 4471
rect 22143 4431 22192 4437
rect 22186 4428 22192 4431
rect 22244 4428 22250 4480
rect 25682 4468 25688 4480
rect 25643 4440 25688 4468
rect 25682 4428 25688 4440
rect 25740 4428 25746 4480
rect 25869 4471 25927 4477
rect 25869 4437 25881 4471
rect 25915 4468 25927 4471
rect 25958 4468 25964 4480
rect 25915 4440 25964 4468
rect 25915 4437 25927 4440
rect 25869 4431 25927 4437
rect 25958 4428 25964 4440
rect 26016 4428 26022 4480
rect 26694 4468 26700 4480
rect 26607 4440 26700 4468
rect 26694 4428 26700 4440
rect 26752 4468 26758 4480
rect 28350 4468 28356 4480
rect 26752 4440 28356 4468
rect 26752 4428 26758 4440
rect 28350 4428 28356 4440
rect 28408 4428 28414 4480
rect 1104 4378 29048 4400
rect 1104 4326 7896 4378
rect 7948 4326 7960 4378
rect 8012 4326 8024 4378
rect 8076 4326 8088 4378
rect 8140 4326 8152 4378
rect 8204 4326 14842 4378
rect 14894 4326 14906 4378
rect 14958 4326 14970 4378
rect 15022 4326 15034 4378
rect 15086 4326 15098 4378
rect 15150 4326 21788 4378
rect 21840 4326 21852 4378
rect 21904 4326 21916 4378
rect 21968 4326 21980 4378
rect 22032 4326 22044 4378
rect 22096 4326 28734 4378
rect 28786 4326 28798 4378
rect 28850 4326 28862 4378
rect 28914 4326 28926 4378
rect 28978 4326 28990 4378
rect 29042 4326 29048 4378
rect 1104 4304 29048 4326
rect 6730 4224 6736 4276
rect 6788 4264 6794 4276
rect 10594 4264 10600 4276
rect 6788 4236 10600 4264
rect 6788 4224 6794 4236
rect 4338 4196 4344 4208
rect 3804 4168 4344 4196
rect 3326 4128 3332 4140
rect 3287 4100 3332 4128
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 3804 4137 3832 4168
rect 4338 4156 4344 4168
rect 4396 4156 4402 4208
rect 5074 4156 5080 4208
rect 5132 4156 5138 4208
rect 3789 4131 3847 4137
rect 3789 4097 3801 4131
rect 3835 4097 3847 4131
rect 6638 4128 6644 4140
rect 6599 4100 6644 4128
rect 3789 4091 3847 4097
rect 6638 4088 6644 4100
rect 6696 4088 6702 4140
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 6880 4100 7389 4128
rect 6880 4088 6886 4100
rect 7377 4097 7389 4100
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 7745 4131 7803 4137
rect 7745 4097 7757 4131
rect 7791 4128 7803 4131
rect 7852 4128 7880 4236
rect 10594 4224 10600 4236
rect 10652 4224 10658 4276
rect 11054 4264 11060 4276
rect 11015 4236 11060 4264
rect 11054 4224 11060 4236
rect 11112 4224 11118 4276
rect 27706 4264 27712 4276
rect 25884 4236 26234 4264
rect 27667 4236 27712 4264
rect 10870 4196 10876 4208
rect 10810 4168 10876 4196
rect 10870 4156 10876 4168
rect 10928 4156 10934 4208
rect 13630 4156 13636 4208
rect 13688 4156 13694 4208
rect 25682 4156 25688 4208
rect 25740 4196 25746 4208
rect 25884 4196 25912 4236
rect 25740 4168 25912 4196
rect 26206 4196 26234 4236
rect 27706 4224 27712 4236
rect 27764 4224 27770 4276
rect 28258 4264 28264 4276
rect 28219 4236 28264 4264
rect 28258 4224 28264 4236
rect 28316 4224 28322 4276
rect 27433 4199 27491 4205
rect 27433 4196 27445 4199
rect 26206 4168 27445 4196
rect 25740 4156 25746 4168
rect 7791 4100 7880 4128
rect 7791 4097 7803 4100
rect 7745 4091 7803 4097
rect 4065 4063 4123 4069
rect 4065 4060 4077 4063
rect 3896 4032 4077 4060
rect 3237 3995 3295 4001
rect 3237 3961 3249 3995
rect 3283 3992 3295 3995
rect 3896 3992 3924 4032
rect 4065 4029 4077 4032
rect 4111 4029 4123 4063
rect 4065 4023 4123 4029
rect 3283 3964 3924 3992
rect 7392 3992 7420 4091
rect 11054 4088 11060 4140
rect 11112 4128 11118 4140
rect 11701 4131 11759 4137
rect 11701 4128 11713 4131
rect 11112 4100 11713 4128
rect 11112 4088 11118 4100
rect 11701 4097 11713 4100
rect 11747 4128 11759 4131
rect 12158 4128 12164 4140
rect 11747 4100 12164 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 17218 4128 17224 4140
rect 17179 4100 17224 4128
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 19817 4131 19875 4137
rect 19817 4097 19829 4131
rect 19863 4128 19875 4131
rect 19978 4128 19984 4140
rect 19863 4100 19984 4128
rect 19863 4097 19875 4100
rect 19817 4091 19875 4097
rect 19978 4088 19984 4100
rect 20036 4088 20042 4140
rect 23376 4131 23434 4137
rect 23376 4097 23388 4131
rect 23422 4128 23434 4131
rect 24670 4128 24676 4140
rect 23422 4100 24676 4128
rect 23422 4097 23434 4100
rect 23376 4091 23434 4097
rect 24670 4088 24676 4100
rect 24728 4088 24734 4140
rect 25590 4128 25596 4140
rect 25551 4100 25596 4128
rect 25590 4088 25596 4100
rect 25648 4088 25654 4140
rect 25792 4137 25820 4168
rect 27433 4165 27445 4168
rect 27479 4165 27491 4199
rect 27433 4159 27491 4165
rect 25777 4131 25835 4137
rect 25777 4097 25789 4131
rect 25823 4128 25835 4131
rect 25823 4100 25857 4128
rect 25823 4097 25835 4100
rect 25777 4091 25835 4097
rect 25958 4088 25964 4140
rect 26016 4128 26022 4140
rect 26234 4128 26240 4140
rect 26016 4100 26061 4128
rect 26147 4100 26240 4128
rect 26016 4088 26022 4100
rect 26234 4088 26240 4100
rect 26292 4128 26298 4140
rect 27157 4131 27215 4137
rect 27157 4128 27169 4131
rect 26292 4100 27169 4128
rect 26292 4088 26298 4100
rect 27157 4097 27169 4100
rect 27203 4097 27215 4131
rect 27157 4091 27215 4097
rect 27246 4088 27252 4140
rect 27304 4128 27310 4140
rect 27341 4131 27399 4137
rect 27341 4128 27353 4131
rect 27304 4100 27353 4128
rect 27304 4088 27310 4100
rect 27341 4097 27353 4100
rect 27387 4097 27399 4131
rect 27341 4091 27399 4097
rect 27522 4088 27528 4140
rect 27580 4128 27586 4140
rect 27724 4128 27752 4224
rect 28169 4131 28227 4137
rect 28169 4128 28181 4131
rect 27580 4100 27673 4128
rect 27724 4100 28181 4128
rect 27580 4088 27586 4100
rect 28169 4097 28181 4100
rect 28215 4097 28227 4131
rect 28350 4128 28356 4140
rect 28311 4100 28356 4128
rect 28169 4091 28227 4097
rect 28350 4088 28356 4100
rect 28408 4088 28414 4140
rect 8294 4060 8300 4072
rect 8255 4032 8300 4060
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 9306 4060 9312 4072
rect 9267 4032 9312 4060
rect 9306 4020 9312 4032
rect 9364 4020 9370 4072
rect 9585 4063 9643 4069
rect 9585 4029 9597 4063
rect 9631 4060 9643 4063
rect 9674 4060 9680 4072
rect 9631 4032 9680 4060
rect 9631 4029 9643 4032
rect 9585 4023 9643 4029
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 12618 4020 12624 4072
rect 12676 4060 12682 4072
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12676 4032 12909 4060
rect 12676 4020 12682 4032
rect 12897 4029 12909 4032
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 13998 4060 14004 4072
rect 13311 4032 14004 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 14274 4020 14280 4072
rect 14332 4060 14338 4072
rect 14691 4063 14749 4069
rect 14691 4060 14703 4063
rect 14332 4032 14703 4060
rect 14332 4020 14338 4032
rect 14691 4029 14703 4032
rect 14737 4029 14749 4063
rect 14691 4023 14749 4029
rect 16114 4020 16120 4072
rect 16172 4060 16178 4072
rect 17129 4063 17187 4069
rect 17129 4060 17141 4063
rect 16172 4032 17141 4060
rect 16172 4020 16178 4032
rect 17129 4029 17141 4032
rect 17175 4029 17187 4063
rect 17129 4023 17187 4029
rect 20073 4063 20131 4069
rect 20073 4029 20085 4063
rect 20119 4060 20131 4063
rect 20622 4060 20628 4072
rect 20119 4032 20628 4060
rect 20119 4029 20131 4032
rect 20073 4023 20131 4029
rect 20622 4020 20628 4032
rect 20680 4020 20686 4072
rect 23109 4063 23167 4069
rect 23109 4060 23121 4063
rect 22066 4032 23121 4060
rect 7392 3964 8156 3992
rect 3283 3961 3295 3964
rect 3237 3955 3295 3961
rect 3326 3884 3332 3936
rect 3384 3924 3390 3936
rect 5534 3924 5540 3936
rect 3384 3896 5540 3924
rect 3384 3884 3390 3896
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 6733 3927 6791 3933
rect 6733 3893 6745 3927
rect 6779 3924 6791 3927
rect 7006 3924 7012 3936
rect 6779 3896 7012 3924
rect 6779 3893 6791 3896
rect 6733 3887 6791 3893
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 8128 3924 8156 3964
rect 9766 3924 9772 3936
rect 8128 3896 9772 3924
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 11793 3927 11851 3933
rect 11793 3893 11805 3927
rect 11839 3924 11851 3927
rect 12250 3924 12256 3936
rect 11839 3896 12256 3924
rect 11839 3893 11851 3896
rect 11793 3887 11851 3893
rect 12250 3884 12256 3896
rect 12308 3884 12314 3936
rect 14642 3884 14648 3936
rect 14700 3924 14706 3936
rect 16853 3927 16911 3933
rect 16853 3924 16865 3927
rect 14700 3896 16865 3924
rect 14700 3884 14706 3896
rect 16853 3893 16865 3896
rect 16899 3893 16911 3927
rect 16853 3887 16911 3893
rect 18693 3927 18751 3933
rect 18693 3893 18705 3927
rect 18739 3924 18751 3927
rect 19702 3924 19708 3936
rect 18739 3896 19708 3924
rect 18739 3893 18751 3896
rect 18693 3887 18751 3893
rect 19702 3884 19708 3896
rect 19760 3884 19766 3936
rect 19794 3884 19800 3936
rect 19852 3924 19858 3936
rect 22066 3924 22094 4032
rect 23109 4029 23121 4032
rect 23155 4029 23167 4063
rect 23109 4023 23167 4029
rect 26142 4020 26148 4072
rect 26200 4060 26206 4072
rect 27540 4060 27568 4088
rect 26200 4032 27568 4060
rect 26200 4020 26206 4032
rect 19852 3896 22094 3924
rect 24489 3927 24547 3933
rect 19852 3884 19858 3896
rect 24489 3893 24501 3927
rect 24535 3924 24547 3927
rect 25590 3924 25596 3936
rect 24535 3896 25596 3924
rect 24535 3893 24547 3896
rect 24489 3887 24547 3893
rect 25590 3884 25596 3896
rect 25648 3884 25654 3936
rect 26237 3927 26295 3933
rect 26237 3893 26249 3927
rect 26283 3924 26295 3927
rect 27154 3924 27160 3936
rect 26283 3896 27160 3924
rect 26283 3893 26295 3896
rect 26237 3887 26295 3893
rect 27154 3884 27160 3896
rect 27212 3884 27218 3936
rect 1104 3834 28888 3856
rect 1104 3782 4423 3834
rect 4475 3782 4487 3834
rect 4539 3782 4551 3834
rect 4603 3782 4615 3834
rect 4667 3782 4679 3834
rect 4731 3782 11369 3834
rect 11421 3782 11433 3834
rect 11485 3782 11497 3834
rect 11549 3782 11561 3834
rect 11613 3782 11625 3834
rect 11677 3782 18315 3834
rect 18367 3782 18379 3834
rect 18431 3782 18443 3834
rect 18495 3782 18507 3834
rect 18559 3782 18571 3834
rect 18623 3782 25261 3834
rect 25313 3782 25325 3834
rect 25377 3782 25389 3834
rect 25441 3782 25453 3834
rect 25505 3782 25517 3834
rect 25569 3782 28888 3834
rect 1104 3760 28888 3782
rect 6638 3680 6644 3732
rect 6696 3720 6702 3732
rect 6696 3692 8524 3720
rect 6696 3680 6702 3692
rect 6730 3652 6736 3664
rect 4448 3624 6736 3652
rect 4154 3584 4160 3596
rect 4115 3556 4160 3584
rect 4154 3544 4160 3556
rect 4212 3544 4218 3596
rect 2498 3476 2504 3528
rect 2556 3516 2562 3528
rect 4448 3525 4476 3624
rect 6730 3612 6736 3624
rect 6788 3612 6794 3664
rect 8496 3661 8524 3692
rect 9306 3680 9312 3732
rect 9364 3720 9370 3732
rect 10137 3723 10195 3729
rect 10137 3720 10149 3723
rect 9364 3692 10149 3720
rect 9364 3680 9370 3692
rect 10137 3689 10149 3692
rect 10183 3689 10195 3723
rect 10137 3683 10195 3689
rect 10781 3723 10839 3729
rect 10781 3689 10793 3723
rect 10827 3720 10839 3723
rect 11054 3720 11060 3732
rect 10827 3692 11060 3720
rect 10827 3689 10839 3692
rect 10781 3683 10839 3689
rect 8481 3655 8539 3661
rect 8481 3621 8493 3655
rect 8527 3652 8539 3655
rect 9398 3652 9404 3664
rect 8527 3624 9404 3652
rect 8527 3621 8539 3624
rect 8481 3615 8539 3621
rect 9398 3612 9404 3624
rect 9456 3612 9462 3664
rect 5074 3584 5080 3596
rect 5035 3556 5080 3584
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 7006 3584 7012 3596
rect 6967 3556 7012 3584
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 4433 3519 4491 3525
rect 4433 3516 4445 3519
rect 2556 3488 4445 3516
rect 2556 3476 2562 3488
rect 4433 3485 4445 3488
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 6273 3519 6331 3525
rect 6273 3485 6285 3519
rect 6319 3485 6331 3519
rect 6273 3479 6331 3485
rect 6733 3519 6791 3525
rect 6733 3485 6745 3519
rect 6779 3485 6791 3519
rect 8294 3516 8300 3528
rect 8142 3488 8300 3516
rect 6733 3479 6791 3485
rect 6178 3380 6184 3392
rect 6139 3352 6184 3380
rect 6178 3340 6184 3352
rect 6236 3340 6242 3392
rect 6288 3380 6316 3479
rect 6748 3448 6776 3479
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 10229 3519 10287 3525
rect 10229 3485 10241 3519
rect 10275 3516 10287 3519
rect 10796 3516 10824 3683
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 11882 3680 11888 3732
rect 11940 3720 11946 3732
rect 16114 3720 16120 3732
rect 11940 3692 15700 3720
rect 16075 3692 16120 3720
rect 11940 3680 11946 3692
rect 15672 3652 15700 3692
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 19794 3720 19800 3732
rect 16546 3692 19800 3720
rect 16546 3652 16574 3692
rect 19794 3680 19800 3692
rect 19852 3680 19858 3732
rect 19978 3720 19984 3732
rect 19939 3692 19984 3720
rect 19978 3680 19984 3692
rect 20036 3680 20042 3732
rect 22787 3723 22845 3729
rect 22787 3689 22799 3723
rect 22833 3720 22845 3723
rect 22922 3720 22928 3732
rect 22833 3692 22928 3720
rect 22833 3689 22845 3692
rect 22787 3683 22845 3689
rect 22922 3680 22928 3692
rect 22980 3680 22986 3732
rect 24670 3720 24676 3732
rect 24631 3692 24676 3720
rect 24670 3680 24676 3692
rect 24728 3680 24734 3732
rect 25869 3723 25927 3729
rect 25869 3689 25881 3723
rect 25915 3720 25927 3723
rect 26142 3720 26148 3732
rect 25915 3692 26148 3720
rect 25915 3689 25927 3692
rect 25869 3683 25927 3689
rect 26142 3680 26148 3692
rect 26200 3680 26206 3732
rect 15672 3624 16574 3652
rect 12250 3584 12256 3596
rect 12211 3556 12256 3584
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 16574 3544 16580 3596
rect 16632 3584 16638 3596
rect 19518 3584 19524 3596
rect 16632 3556 16677 3584
rect 19479 3556 19524 3584
rect 16632 3544 16638 3556
rect 19518 3544 19524 3556
rect 19576 3544 19582 3596
rect 21361 3587 21419 3593
rect 21361 3553 21373 3587
rect 21407 3584 21419 3587
rect 22186 3584 22192 3596
rect 21407 3556 22192 3584
rect 21407 3553 21419 3556
rect 21361 3547 21419 3553
rect 22186 3544 22192 3556
rect 22244 3544 22250 3596
rect 10275 3488 10824 3516
rect 12529 3519 12587 3525
rect 10275 3485 10287 3488
rect 10229 3479 10287 3485
rect 12529 3485 12541 3519
rect 12575 3516 12587 3519
rect 12618 3516 12624 3528
rect 12575 3488 12624 3516
rect 12575 3485 12587 3488
rect 12529 3479 12587 3485
rect 12618 3476 12624 3488
rect 12676 3516 12682 3528
rect 13722 3516 13728 3528
rect 12676 3488 13728 3516
rect 12676 3476 12682 3488
rect 13722 3476 13728 3488
rect 13780 3516 13786 3528
rect 13906 3516 13912 3528
rect 13780 3488 13912 3516
rect 13780 3476 13786 3488
rect 13906 3476 13912 3488
rect 13964 3516 13970 3528
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 13964 3488 14749 3516
rect 13964 3476 13970 3488
rect 14737 3485 14749 3488
rect 14783 3516 14795 3519
rect 16298 3516 16304 3528
rect 14783 3488 16304 3516
rect 14783 3485 14795 3488
rect 14737 3479 14795 3485
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 16844 3519 16902 3525
rect 16844 3485 16856 3519
rect 16890 3516 16902 3519
rect 17218 3516 17224 3528
rect 16890 3488 17224 3516
rect 16890 3485 16902 3488
rect 16844 3479 16902 3485
rect 17218 3476 17224 3488
rect 17276 3516 17282 3528
rect 19610 3516 19616 3528
rect 17276 3488 19616 3516
rect 17276 3476 17282 3488
rect 19610 3476 19616 3488
rect 19668 3476 19674 3528
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 20993 3519 21051 3525
rect 20993 3516 21005 3519
rect 20680 3488 21005 3516
rect 20680 3476 20686 3488
rect 20993 3485 21005 3488
rect 21039 3485 21051 3519
rect 20993 3479 21051 3485
rect 24765 3519 24823 3525
rect 24765 3485 24777 3519
rect 24811 3516 24823 3519
rect 25590 3516 25596 3528
rect 24811 3488 25596 3516
rect 24811 3485 24823 3488
rect 24765 3479 24823 3485
rect 25590 3476 25596 3488
rect 25648 3476 25654 3528
rect 27246 3516 27252 3528
rect 27207 3488 27252 3516
rect 27246 3476 27252 3488
rect 27304 3476 27310 3528
rect 27522 3476 27528 3528
rect 27580 3516 27586 3528
rect 27709 3519 27767 3525
rect 27709 3516 27721 3519
rect 27580 3488 27721 3516
rect 27580 3476 27586 3488
rect 27709 3485 27721 3488
rect 27755 3485 27767 3519
rect 27709 3479 27767 3485
rect 7282 3448 7288 3460
rect 6748 3420 7288 3448
rect 7282 3408 7288 3420
rect 7340 3408 7346 3460
rect 11698 3408 11704 3460
rect 11756 3408 11762 3460
rect 14982 3451 15040 3457
rect 14982 3448 14994 3451
rect 14752 3420 14994 3448
rect 14752 3392 14780 3420
rect 14982 3417 14994 3420
rect 15028 3417 15040 3451
rect 14982 3411 15040 3417
rect 22278 3408 22284 3460
rect 22336 3408 22342 3460
rect 27004 3451 27062 3457
rect 27004 3417 27016 3451
rect 27050 3448 27062 3451
rect 27801 3451 27859 3457
rect 27801 3448 27813 3451
rect 27050 3420 27813 3448
rect 27050 3417 27062 3420
rect 27004 3411 27062 3417
rect 27801 3417 27813 3420
rect 27847 3417 27859 3451
rect 27801 3411 27859 3417
rect 7098 3380 7104 3392
rect 6288 3352 7104 3380
rect 7098 3340 7104 3352
rect 7156 3340 7162 3392
rect 14734 3340 14740 3392
rect 14792 3340 14798 3392
rect 17954 3380 17960 3392
rect 17915 3352 17960 3380
rect 17954 3340 17960 3352
rect 18012 3340 18018 3392
rect 1104 3290 29048 3312
rect 1104 3238 7896 3290
rect 7948 3238 7960 3290
rect 8012 3238 8024 3290
rect 8076 3238 8088 3290
rect 8140 3238 8152 3290
rect 8204 3238 14842 3290
rect 14894 3238 14906 3290
rect 14958 3238 14970 3290
rect 15022 3238 15034 3290
rect 15086 3238 15098 3290
rect 15150 3238 21788 3290
rect 21840 3238 21852 3290
rect 21904 3238 21916 3290
rect 21968 3238 21980 3290
rect 22032 3238 22044 3290
rect 22096 3238 28734 3290
rect 28786 3238 28798 3290
rect 28850 3238 28862 3290
rect 28914 3238 28926 3290
rect 28978 3238 28990 3290
rect 29042 3238 29048 3290
rect 1104 3216 29048 3238
rect 6178 3136 6184 3188
rect 6236 3176 6242 3188
rect 10870 3176 10876 3188
rect 6236 3148 8156 3176
rect 10831 3148 10876 3176
rect 6236 3136 6242 3148
rect 4154 3068 4160 3120
rect 4212 3108 4218 3120
rect 4249 3111 4307 3117
rect 4249 3108 4261 3111
rect 4212 3080 4261 3108
rect 4212 3068 4218 3080
rect 4249 3077 4261 3080
rect 4295 3077 4307 3111
rect 4249 3071 4307 3077
rect 7374 3068 7380 3120
rect 7432 3068 7438 3120
rect 8128 3117 8156 3148
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 13998 3176 14004 3188
rect 13959 3148 14004 3176
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 14734 3136 14740 3188
rect 14792 3176 14798 3188
rect 14921 3179 14979 3185
rect 14921 3176 14933 3179
rect 14792 3148 14933 3176
rect 14792 3136 14798 3148
rect 14921 3145 14933 3148
rect 14967 3145 14979 3179
rect 14921 3139 14979 3145
rect 18969 3179 19027 3185
rect 18969 3145 18981 3179
rect 19015 3176 19027 3179
rect 19518 3176 19524 3188
rect 19015 3148 19524 3176
rect 19015 3145 19027 3148
rect 18969 3139 19027 3145
rect 19518 3136 19524 3148
rect 19576 3136 19582 3188
rect 19610 3136 19616 3188
rect 19668 3176 19674 3188
rect 23753 3179 23811 3185
rect 23753 3176 23765 3179
rect 19668 3148 23765 3176
rect 19668 3136 19674 3148
rect 8113 3111 8171 3117
rect 8113 3077 8125 3111
rect 8159 3077 8171 3111
rect 8113 3071 8171 3077
rect 17856 3111 17914 3117
rect 17856 3077 17868 3111
rect 17902 3108 17914 3111
rect 17954 3108 17960 3120
rect 17902 3080 17960 3108
rect 17902 3077 17914 3080
rect 17856 3071 17914 3077
rect 17954 3068 17960 3080
rect 18012 3068 18018 3120
rect 5997 3043 6055 3049
rect 5997 3009 6009 3043
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 6012 2972 6040 3003
rect 8386 3000 8392 3052
rect 8444 3040 8450 3052
rect 8444 3012 8489 3040
rect 8444 3000 8450 3012
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 9824 3012 9873 3040
rect 9824 3000 9830 3012
rect 9861 3009 9873 3012
rect 9907 3009 9919 3043
rect 9861 3003 9919 3009
rect 10229 3043 10287 3049
rect 10229 3009 10241 3043
rect 10275 3040 10287 3043
rect 10686 3040 10692 3052
rect 10275 3012 10692 3040
rect 10275 3009 10287 3012
rect 10229 3003 10287 3009
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 19812 3049 19840 3148
rect 23753 3145 23765 3148
rect 23799 3145 23811 3179
rect 23753 3139 23811 3145
rect 25685 3179 25743 3185
rect 25685 3145 25697 3179
rect 25731 3176 25743 3179
rect 25958 3176 25964 3188
rect 25731 3148 25964 3176
rect 25731 3145 25743 3148
rect 25685 3139 25743 3145
rect 22738 3068 22744 3120
rect 22796 3068 22802 3120
rect 23768 3108 23796 3139
rect 25958 3136 25964 3148
rect 26016 3136 26022 3188
rect 26237 3179 26295 3185
rect 26237 3145 26249 3179
rect 26283 3176 26295 3179
rect 27246 3176 27252 3188
rect 26283 3148 27252 3176
rect 26283 3145 26295 3148
rect 26237 3139 26295 3145
rect 27246 3136 27252 3148
rect 27304 3136 27310 3188
rect 24550 3111 24608 3117
rect 24550 3108 24562 3111
rect 23768 3080 24562 3108
rect 24550 3077 24562 3080
rect 24596 3077 24608 3111
rect 24550 3071 24608 3077
rect 12877 3043 12935 3049
rect 12877 3040 12889 3043
rect 12492 3012 12889 3040
rect 12492 3000 12498 3012
rect 12877 3009 12889 3012
rect 12923 3009 12935 3043
rect 12877 3003 12935 3009
rect 16045 3043 16103 3049
rect 16045 3009 16057 3043
rect 16091 3040 16103 3043
rect 19797 3043 19855 3049
rect 16091 3012 19472 3040
rect 16091 3009 16103 3012
rect 16045 3003 16103 3009
rect 6914 2972 6920 2984
rect 6012 2944 6920 2972
rect 6914 2932 6920 2944
rect 6972 2932 6978 2984
rect 12618 2972 12624 2984
rect 12579 2944 12624 2972
rect 12618 2932 12624 2944
rect 12676 2932 12682 2984
rect 16298 2972 16304 2984
rect 16259 2944 16304 2972
rect 16298 2932 16304 2944
rect 16356 2932 16362 2984
rect 19444 2981 19472 3012
rect 19797 3009 19809 3043
rect 19843 3009 19855 3043
rect 19797 3003 19855 3009
rect 20622 3000 20628 3052
rect 20680 3040 20686 3052
rect 22005 3043 22063 3049
rect 22005 3040 22017 3043
rect 20680 3012 22017 3040
rect 20680 3000 20686 3012
rect 22005 3009 22017 3012
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 25590 3000 25596 3052
rect 25648 3040 25654 3052
rect 26145 3043 26203 3049
rect 26145 3040 26157 3043
rect 25648 3012 26157 3040
rect 25648 3000 25654 3012
rect 26145 3009 26157 3012
rect 26191 3009 26203 3043
rect 27154 3040 27160 3052
rect 27115 3012 27160 3040
rect 26145 3003 26203 3009
rect 27154 3000 27160 3012
rect 27212 3000 27218 3052
rect 27341 3043 27399 3049
rect 27341 3009 27353 3043
rect 27387 3040 27399 3043
rect 27430 3040 27436 3052
rect 27387 3012 27436 3040
rect 27387 3009 27399 3012
rect 27341 3003 27399 3009
rect 27430 3000 27436 3012
rect 27488 3000 27494 3052
rect 17589 2975 17647 2981
rect 17589 2941 17601 2975
rect 17635 2941 17647 2975
rect 17589 2935 17647 2941
rect 19429 2975 19487 2981
rect 19429 2941 19441 2975
rect 19475 2941 19487 2975
rect 19702 2972 19708 2984
rect 19663 2944 19708 2972
rect 19429 2935 19487 2941
rect 6641 2907 6699 2913
rect 6641 2873 6653 2907
rect 6687 2904 6699 2907
rect 7098 2904 7104 2916
rect 6687 2876 7104 2904
rect 6687 2873 6699 2876
rect 6641 2867 6699 2873
rect 7098 2864 7104 2876
rect 7156 2864 7162 2916
rect 17604 2836 17632 2935
rect 19702 2932 19708 2944
rect 19760 2932 19766 2984
rect 22281 2975 22339 2981
rect 22281 2941 22293 2975
rect 22327 2972 22339 2975
rect 22922 2972 22928 2984
rect 22327 2944 22928 2972
rect 22327 2941 22339 2944
rect 22281 2935 22339 2941
rect 22922 2932 22928 2944
rect 22980 2932 22986 2984
rect 23290 2932 23296 2984
rect 23348 2972 23354 2984
rect 24305 2975 24363 2981
rect 24305 2972 24317 2975
rect 23348 2944 24317 2972
rect 23348 2932 23354 2944
rect 24305 2941 24317 2944
rect 24351 2941 24363 2975
rect 24305 2935 24363 2941
rect 20622 2836 20628 2848
rect 17604 2808 20628 2836
rect 20622 2796 20628 2808
rect 20680 2796 20686 2848
rect 27157 2839 27215 2845
rect 27157 2805 27169 2839
rect 27203 2836 27215 2839
rect 27890 2836 27896 2848
rect 27203 2808 27896 2836
rect 27203 2805 27215 2808
rect 27157 2799 27215 2805
rect 27890 2796 27896 2808
rect 27948 2796 27954 2848
rect 1104 2746 28888 2768
rect 1104 2694 4423 2746
rect 4475 2694 4487 2746
rect 4539 2694 4551 2746
rect 4603 2694 4615 2746
rect 4667 2694 4679 2746
rect 4731 2694 11369 2746
rect 11421 2694 11433 2746
rect 11485 2694 11497 2746
rect 11549 2694 11561 2746
rect 11613 2694 11625 2746
rect 11677 2694 18315 2746
rect 18367 2694 18379 2746
rect 18431 2694 18443 2746
rect 18495 2694 18507 2746
rect 18559 2694 18571 2746
rect 18623 2694 25261 2746
rect 25313 2694 25325 2746
rect 25377 2694 25389 2746
rect 25441 2694 25453 2746
rect 25505 2694 25517 2746
rect 25569 2694 28888 2746
rect 1104 2672 28888 2694
rect 7282 2632 7288 2644
rect 7243 2604 7288 2632
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 12345 2635 12403 2641
rect 12345 2601 12357 2635
rect 12391 2632 12403 2635
rect 12434 2632 12440 2644
rect 12391 2604 12440 2632
rect 12391 2601 12403 2604
rect 12345 2595 12403 2601
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 13722 2496 13728 2508
rect 13683 2468 13728 2496
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7156 2400 7389 2428
rect 7156 2388 7162 2400
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 27890 2428 27896 2440
rect 27851 2400 27896 2428
rect 7377 2391 7435 2397
rect 27890 2388 27896 2400
rect 27948 2388 27954 2440
rect 13480 2363 13538 2369
rect 13480 2329 13492 2363
rect 13526 2360 13538 2363
rect 14642 2360 14648 2372
rect 13526 2332 14648 2360
rect 13526 2329 13538 2332
rect 13480 2323 13538 2329
rect 14642 2320 14648 2332
rect 14700 2320 14706 2372
rect 28166 2360 28172 2372
rect 28127 2332 28172 2360
rect 28166 2320 28172 2332
rect 28224 2320 28230 2372
rect 1104 2202 29048 2224
rect 1104 2150 7896 2202
rect 7948 2150 7960 2202
rect 8012 2150 8024 2202
rect 8076 2150 8088 2202
rect 8140 2150 8152 2202
rect 8204 2150 14842 2202
rect 14894 2150 14906 2202
rect 14958 2150 14970 2202
rect 15022 2150 15034 2202
rect 15086 2150 15098 2202
rect 15150 2150 21788 2202
rect 21840 2150 21852 2202
rect 21904 2150 21916 2202
rect 21968 2150 21980 2202
rect 22032 2150 22044 2202
rect 22096 2150 28734 2202
rect 28786 2150 28798 2202
rect 28850 2150 28862 2202
rect 28914 2150 28926 2202
rect 28978 2150 28990 2202
rect 29042 2150 29048 2202
rect 1104 2128 29048 2150
<< via1 >>
rect 4423 27718 4475 27770
rect 4487 27718 4539 27770
rect 4551 27718 4603 27770
rect 4615 27718 4667 27770
rect 4679 27718 4731 27770
rect 11369 27718 11421 27770
rect 11433 27718 11485 27770
rect 11497 27718 11549 27770
rect 11561 27718 11613 27770
rect 11625 27718 11677 27770
rect 18315 27718 18367 27770
rect 18379 27718 18431 27770
rect 18443 27718 18495 27770
rect 18507 27718 18559 27770
rect 18571 27718 18623 27770
rect 25261 27718 25313 27770
rect 25325 27718 25377 27770
rect 25389 27718 25441 27770
rect 25453 27718 25505 27770
rect 25517 27718 25569 27770
rect 17684 27480 17736 27532
rect 27896 27480 27948 27532
rect 3332 27412 3384 27464
rect 5724 27412 5776 27464
rect 9588 27455 9640 27464
rect 9588 27421 9597 27455
rect 9597 27421 9631 27455
rect 9631 27421 9640 27455
rect 9588 27412 9640 27421
rect 13084 27455 13136 27464
rect 13084 27421 13093 27455
rect 13093 27421 13127 27455
rect 13127 27421 13136 27455
rect 13084 27412 13136 27421
rect 17040 27455 17092 27464
rect 17040 27421 17049 27455
rect 17049 27421 17083 27455
rect 17083 27421 17092 27455
rect 17040 27412 17092 27421
rect 20628 27455 20680 27464
rect 20628 27421 20637 27455
rect 20637 27421 20671 27455
rect 20671 27421 20680 27455
rect 20628 27412 20680 27421
rect 22284 27412 22336 27464
rect 24124 27412 24176 27464
rect 27712 27455 27764 27464
rect 27712 27421 27721 27455
rect 27721 27421 27755 27455
rect 27755 27421 27764 27455
rect 27712 27412 27764 27421
rect 4528 27344 4580 27396
rect 12624 27344 12676 27396
rect 13728 27344 13780 27396
rect 28080 27387 28132 27396
rect 28080 27353 28089 27387
rect 28089 27353 28123 27387
rect 28123 27353 28132 27387
rect 28080 27344 28132 27353
rect 3148 27319 3200 27328
rect 3148 27285 3157 27319
rect 3157 27285 3191 27319
rect 3191 27285 3200 27319
rect 3148 27276 3200 27285
rect 6920 27319 6972 27328
rect 6920 27285 6929 27319
rect 6929 27285 6963 27319
rect 6963 27285 6972 27319
rect 16948 27319 17000 27328
rect 6920 27276 6972 27285
rect 16948 27285 16957 27319
rect 16957 27285 16991 27319
rect 16991 27285 17000 27319
rect 16948 27276 17000 27285
rect 20904 27319 20956 27328
rect 20904 27285 20913 27319
rect 20913 27285 20947 27319
rect 20947 27285 20956 27319
rect 20904 27276 20956 27285
rect 22192 27276 22244 27328
rect 24952 27319 25004 27328
rect 24952 27285 24961 27319
rect 24961 27285 24995 27319
rect 24995 27285 25004 27319
rect 24952 27276 25004 27285
rect 7896 27174 7948 27226
rect 7960 27174 8012 27226
rect 8024 27174 8076 27226
rect 8088 27174 8140 27226
rect 8152 27174 8204 27226
rect 14842 27174 14894 27226
rect 14906 27174 14958 27226
rect 14970 27174 15022 27226
rect 15034 27174 15086 27226
rect 15098 27174 15150 27226
rect 21788 27174 21840 27226
rect 21852 27174 21904 27226
rect 21916 27174 21968 27226
rect 21980 27174 22032 27226
rect 22044 27174 22096 27226
rect 28734 27174 28786 27226
rect 28798 27174 28850 27226
rect 28862 27174 28914 27226
rect 28926 27174 28978 27226
rect 28990 27174 29042 27226
rect 3424 27004 3476 27056
rect 4528 27047 4580 27056
rect 4528 27013 4537 27047
rect 4537 27013 4571 27047
rect 4571 27013 4580 27047
rect 4528 27004 4580 27013
rect 5264 27004 5316 27056
rect 16948 27047 17000 27056
rect 16948 27013 16957 27047
rect 16957 27013 16991 27047
rect 16991 27013 17000 27047
rect 16948 27004 17000 27013
rect 2872 26979 2924 26988
rect 2872 26945 2906 26979
rect 2906 26945 2924 26979
rect 2872 26936 2924 26945
rect 6920 26936 6972 26988
rect 8300 26936 8352 26988
rect 9496 26936 9548 26988
rect 10416 26979 10468 26988
rect 10416 26945 10425 26979
rect 10425 26945 10459 26979
rect 10459 26945 10468 26979
rect 10416 26936 10468 26945
rect 12256 26936 12308 26988
rect 15292 26936 15344 26988
rect 19800 26979 19852 26988
rect 19800 26945 19809 26979
rect 19809 26945 19843 26979
rect 19843 26945 19852 26979
rect 19800 26936 19852 26945
rect 19984 26979 20036 26988
rect 19984 26945 19993 26979
rect 19993 26945 20027 26979
rect 20027 26945 20036 26979
rect 19984 26936 20036 26945
rect 22836 27004 22888 27056
rect 22284 26936 22336 26988
rect 23020 26979 23072 26988
rect 23020 26945 23029 26979
rect 23029 26945 23063 26979
rect 23063 26945 23072 26979
rect 23020 26936 23072 26945
rect 25780 26979 25832 26988
rect 25780 26945 25789 26979
rect 25789 26945 25823 26979
rect 25823 26945 25832 26979
rect 25780 26936 25832 26945
rect 27528 27004 27580 27056
rect 27712 26936 27764 26988
rect 27896 26979 27948 26988
rect 27896 26945 27905 26979
rect 27905 26945 27939 26979
rect 27939 26945 27948 26979
rect 27896 26936 27948 26945
rect 8760 26911 8812 26920
rect 8760 26877 8769 26911
rect 8769 26877 8803 26911
rect 8803 26877 8812 26911
rect 8760 26868 8812 26877
rect 9680 26868 9732 26920
rect 12532 26911 12584 26920
rect 12532 26877 12541 26911
rect 12541 26877 12575 26911
rect 12575 26877 12584 26911
rect 12532 26868 12584 26877
rect 12808 26911 12860 26920
rect 12808 26877 12817 26911
rect 12817 26877 12851 26911
rect 12851 26877 12860 26911
rect 12808 26868 12860 26877
rect 20352 26911 20404 26920
rect 20352 26877 20361 26911
rect 20361 26877 20395 26911
rect 20395 26877 20404 26911
rect 20352 26868 20404 26877
rect 20904 26868 20956 26920
rect 22928 26911 22980 26920
rect 16764 26800 16816 26852
rect 22376 26800 22428 26852
rect 22928 26877 22937 26911
rect 22937 26877 22971 26911
rect 22971 26877 22980 26911
rect 22928 26868 22980 26877
rect 26056 26911 26108 26920
rect 26056 26877 26065 26911
rect 26065 26877 26099 26911
rect 26099 26877 26108 26911
rect 26056 26868 26108 26877
rect 26700 26868 26752 26920
rect 23940 26800 23992 26852
rect 4160 26732 4212 26784
rect 6552 26732 6604 26784
rect 8392 26732 8444 26784
rect 10508 26775 10560 26784
rect 10508 26741 10517 26775
rect 10517 26741 10551 26775
rect 10551 26741 10560 26775
rect 10508 26732 10560 26741
rect 10784 26732 10836 26784
rect 13176 26732 13228 26784
rect 21732 26732 21784 26784
rect 23388 26775 23440 26784
rect 23388 26741 23397 26775
rect 23397 26741 23431 26775
rect 23431 26741 23440 26775
rect 23388 26732 23440 26741
rect 27252 26775 27304 26784
rect 27252 26741 27261 26775
rect 27261 26741 27295 26775
rect 27295 26741 27304 26775
rect 27252 26732 27304 26741
rect 4423 26630 4475 26682
rect 4487 26630 4539 26682
rect 4551 26630 4603 26682
rect 4615 26630 4667 26682
rect 4679 26630 4731 26682
rect 11369 26630 11421 26682
rect 11433 26630 11485 26682
rect 11497 26630 11549 26682
rect 11561 26630 11613 26682
rect 11625 26630 11677 26682
rect 18315 26630 18367 26682
rect 18379 26630 18431 26682
rect 18443 26630 18495 26682
rect 18507 26630 18559 26682
rect 18571 26630 18623 26682
rect 25261 26630 25313 26682
rect 25325 26630 25377 26682
rect 25389 26630 25441 26682
rect 25453 26630 25505 26682
rect 25517 26630 25569 26682
rect 4160 26571 4212 26580
rect 4160 26537 4169 26571
rect 4169 26537 4203 26571
rect 4203 26537 4212 26571
rect 4160 26528 4212 26537
rect 8760 26528 8812 26580
rect 9864 26528 9916 26580
rect 4988 26460 5040 26512
rect 3424 26435 3476 26444
rect 3424 26401 3433 26435
rect 3433 26401 3467 26435
rect 3467 26401 3476 26435
rect 3424 26392 3476 26401
rect 6552 26435 6604 26444
rect 6552 26401 6561 26435
rect 6561 26401 6595 26435
rect 6595 26401 6604 26435
rect 6552 26392 6604 26401
rect 8300 26392 8352 26444
rect 9312 26392 9364 26444
rect 10508 26435 10560 26444
rect 10508 26401 10517 26435
rect 10517 26401 10551 26435
rect 10551 26401 10560 26435
rect 10508 26392 10560 26401
rect 10784 26435 10836 26444
rect 10784 26401 10793 26435
rect 10793 26401 10827 26435
rect 10827 26401 10836 26435
rect 10784 26392 10836 26401
rect 12808 26528 12860 26580
rect 17684 26571 17736 26580
rect 17684 26537 17693 26571
rect 17693 26537 17727 26571
rect 17727 26537 17736 26571
rect 17684 26528 17736 26537
rect 19800 26528 19852 26580
rect 22468 26528 22520 26580
rect 23020 26528 23072 26580
rect 27712 26571 27764 26580
rect 27712 26537 27721 26571
rect 27721 26537 27755 26571
rect 27755 26537 27764 26571
rect 27712 26528 27764 26537
rect 15292 26435 15344 26444
rect 2872 26324 2924 26376
rect 15292 26401 15301 26435
rect 15301 26401 15335 26435
rect 15335 26401 15344 26435
rect 15292 26392 15344 26401
rect 21732 26435 21784 26444
rect 21732 26401 21741 26435
rect 21741 26401 21775 26435
rect 21775 26401 21784 26435
rect 21732 26392 21784 26401
rect 22100 26392 22152 26444
rect 27252 26392 27304 26444
rect 5080 26367 5132 26376
rect 3148 26299 3200 26308
rect 3148 26265 3166 26299
rect 3166 26265 3200 26299
rect 3148 26256 3200 26265
rect 3332 26256 3384 26308
rect 4436 26256 4488 26308
rect 2136 26188 2188 26240
rect 5080 26333 5089 26367
rect 5089 26333 5123 26367
rect 5123 26333 5132 26367
rect 5080 26324 5132 26333
rect 6276 26367 6328 26376
rect 6276 26333 6285 26367
rect 6285 26333 6319 26367
rect 6319 26333 6328 26367
rect 6276 26324 6328 26333
rect 7656 26324 7708 26376
rect 10140 26324 10192 26376
rect 10416 26324 10468 26376
rect 13176 26324 13228 26376
rect 14372 26367 14424 26376
rect 14372 26333 14381 26367
rect 14381 26333 14415 26367
rect 14415 26333 14424 26367
rect 14372 26324 14424 26333
rect 14556 26324 14608 26376
rect 16304 26367 16356 26376
rect 16304 26333 16313 26367
rect 16313 26333 16347 26367
rect 16347 26333 16356 26367
rect 16304 26324 16356 26333
rect 18144 26367 18196 26376
rect 18144 26333 18153 26367
rect 18153 26333 18187 26367
rect 18187 26333 18196 26367
rect 18144 26324 18196 26333
rect 21272 26367 21324 26376
rect 21272 26333 21281 26367
rect 21281 26333 21315 26367
rect 21315 26333 21324 26367
rect 21272 26324 21324 26333
rect 23112 26324 23164 26376
rect 11796 26256 11848 26308
rect 16764 26256 16816 26308
rect 20352 26256 20404 26308
rect 20720 26256 20772 26308
rect 26148 26256 26200 26308
rect 26700 26256 26752 26308
rect 4344 26231 4396 26240
rect 4344 26197 4353 26231
rect 4353 26197 4387 26231
rect 4387 26197 4396 26231
rect 4344 26188 4396 26197
rect 4896 26188 4948 26240
rect 8668 26188 8720 26240
rect 12072 26188 12124 26240
rect 12256 26231 12308 26240
rect 12256 26197 12265 26231
rect 12265 26197 12299 26231
rect 12299 26197 12308 26231
rect 12256 26188 12308 26197
rect 18788 26188 18840 26240
rect 19708 26188 19760 26240
rect 7896 26086 7948 26138
rect 7960 26086 8012 26138
rect 8024 26086 8076 26138
rect 8088 26086 8140 26138
rect 8152 26086 8204 26138
rect 14842 26086 14894 26138
rect 14906 26086 14958 26138
rect 14970 26086 15022 26138
rect 15034 26086 15086 26138
rect 15098 26086 15150 26138
rect 21788 26086 21840 26138
rect 21852 26086 21904 26138
rect 21916 26086 21968 26138
rect 21980 26086 22032 26138
rect 22044 26086 22096 26138
rect 28734 26086 28786 26138
rect 28798 26086 28850 26138
rect 28862 26086 28914 26138
rect 28926 26086 28978 26138
rect 28990 26086 29042 26138
rect 2780 25984 2832 26036
rect 4436 26027 4488 26036
rect 4436 25993 4445 26027
rect 4445 25993 4479 26027
rect 4479 25993 4488 26027
rect 4436 25984 4488 25993
rect 2136 25891 2188 25900
rect 2136 25857 2145 25891
rect 2145 25857 2179 25891
rect 2179 25857 2188 25891
rect 2136 25848 2188 25857
rect 2872 25780 2924 25832
rect 4344 25848 4396 25900
rect 4988 25891 5040 25900
rect 4988 25857 4997 25891
rect 4997 25857 5031 25891
rect 5031 25857 5040 25891
rect 9496 25984 9548 26036
rect 10140 26027 10192 26036
rect 10140 25993 10149 26027
rect 10149 25993 10183 26027
rect 10183 25993 10192 26027
rect 10140 25984 10192 25993
rect 12532 25984 12584 26036
rect 18144 25984 18196 26036
rect 20720 25984 20772 26036
rect 21272 25984 21324 26036
rect 22284 25984 22336 26036
rect 23112 26027 23164 26036
rect 23112 25993 23121 26027
rect 23121 25993 23155 26027
rect 23155 25993 23164 26027
rect 23112 25984 23164 25993
rect 23940 26027 23992 26036
rect 23940 25993 23949 26027
rect 23949 25993 23983 26027
rect 23983 25993 23992 26027
rect 23940 25984 23992 25993
rect 7656 25959 7708 25968
rect 7656 25925 7665 25959
rect 7665 25925 7699 25959
rect 7699 25925 7708 25959
rect 7656 25916 7708 25925
rect 8668 25959 8720 25968
rect 8668 25925 8677 25959
rect 8677 25925 8711 25959
rect 8711 25925 8720 25959
rect 8668 25916 8720 25925
rect 9680 25916 9732 25968
rect 15384 25916 15436 25968
rect 18236 25916 18288 25968
rect 18788 25959 18840 25968
rect 18788 25925 18797 25959
rect 18797 25925 18831 25959
rect 18831 25925 18840 25959
rect 18788 25916 18840 25925
rect 8392 25891 8444 25900
rect 4988 25848 5040 25857
rect 8392 25857 8401 25891
rect 8401 25857 8435 25891
rect 8435 25857 8444 25891
rect 8392 25848 8444 25857
rect 12072 25848 12124 25900
rect 19708 25891 19760 25900
rect 4804 25780 4856 25832
rect 5264 25780 5316 25832
rect 6644 25780 6696 25832
rect 8760 25780 8812 25832
rect 4160 25644 4212 25696
rect 19708 25857 19717 25891
rect 19717 25857 19751 25891
rect 19751 25857 19760 25891
rect 19708 25848 19760 25857
rect 22468 25891 22520 25900
rect 22468 25857 22477 25891
rect 22477 25857 22511 25891
rect 22511 25857 22520 25891
rect 25780 25891 25832 25900
rect 22468 25848 22520 25857
rect 25780 25857 25789 25891
rect 25789 25857 25823 25891
rect 25823 25857 25832 25891
rect 25780 25848 25832 25857
rect 26148 25848 26200 25900
rect 14096 25823 14148 25832
rect 14096 25789 14105 25823
rect 14105 25789 14139 25823
rect 14139 25789 14148 25823
rect 14096 25780 14148 25789
rect 19984 25780 20036 25832
rect 24032 25823 24084 25832
rect 24032 25789 24041 25823
rect 24041 25789 24075 25823
rect 24075 25789 24084 25823
rect 24032 25780 24084 25789
rect 23664 25712 23716 25764
rect 26056 25823 26108 25832
rect 26056 25789 26065 25823
rect 26065 25789 26099 25823
rect 26099 25789 26108 25823
rect 26056 25780 26108 25789
rect 26516 25823 26568 25832
rect 26516 25789 26525 25823
rect 26525 25789 26559 25823
rect 26559 25789 26568 25823
rect 26516 25780 26568 25789
rect 27436 25712 27488 25764
rect 15660 25644 15712 25696
rect 23572 25687 23624 25696
rect 23572 25653 23581 25687
rect 23581 25653 23615 25687
rect 23615 25653 23624 25687
rect 23572 25644 23624 25653
rect 27528 25644 27580 25696
rect 4423 25542 4475 25594
rect 4487 25542 4539 25594
rect 4551 25542 4603 25594
rect 4615 25542 4667 25594
rect 4679 25542 4731 25594
rect 11369 25542 11421 25594
rect 11433 25542 11485 25594
rect 11497 25542 11549 25594
rect 11561 25542 11613 25594
rect 11625 25542 11677 25594
rect 18315 25542 18367 25594
rect 18379 25542 18431 25594
rect 18443 25542 18495 25594
rect 18507 25542 18559 25594
rect 18571 25542 18623 25594
rect 25261 25542 25313 25594
rect 25325 25542 25377 25594
rect 25389 25542 25441 25594
rect 25453 25542 25505 25594
rect 25517 25542 25569 25594
rect 4252 25440 4304 25492
rect 4804 25440 4856 25492
rect 6276 25440 6328 25492
rect 14096 25440 14148 25492
rect 22928 25440 22980 25492
rect 5080 25304 5132 25356
rect 7748 25304 7800 25356
rect 11244 25304 11296 25356
rect 11796 25347 11848 25356
rect 11796 25313 11805 25347
rect 11805 25313 11839 25347
rect 11839 25313 11848 25347
rect 11796 25304 11848 25313
rect 3148 25279 3200 25288
rect 3148 25245 3157 25279
rect 3157 25245 3191 25279
rect 3191 25245 3200 25279
rect 3148 25236 3200 25245
rect 4160 25279 4212 25288
rect 4160 25245 4169 25279
rect 4169 25245 4203 25279
rect 4203 25245 4212 25279
rect 4160 25236 4212 25245
rect 4344 25236 4396 25288
rect 6368 25236 6420 25288
rect 9312 25279 9364 25288
rect 2964 25143 3016 25152
rect 2964 25109 2973 25143
rect 2973 25109 3007 25143
rect 3007 25109 3016 25143
rect 2964 25100 3016 25109
rect 4068 25100 4120 25152
rect 4252 25100 4304 25152
rect 4896 25168 4948 25220
rect 5264 25211 5316 25220
rect 5264 25177 5273 25211
rect 5273 25177 5307 25211
rect 5307 25177 5316 25211
rect 5264 25168 5316 25177
rect 9312 25245 9321 25279
rect 9321 25245 9355 25279
rect 9355 25245 9364 25279
rect 9312 25236 9364 25245
rect 9956 25236 10008 25288
rect 7472 25168 7524 25220
rect 9496 25168 9548 25220
rect 13176 25236 13228 25288
rect 14372 25279 14424 25288
rect 14372 25245 14381 25279
rect 14381 25245 14415 25279
rect 14415 25245 14424 25279
rect 14372 25236 14424 25245
rect 14556 25304 14608 25356
rect 15384 25347 15436 25356
rect 15384 25313 15393 25347
rect 15393 25313 15427 25347
rect 15427 25313 15436 25347
rect 15384 25304 15436 25313
rect 19800 25372 19852 25424
rect 18236 25304 18288 25356
rect 23664 25347 23716 25356
rect 23664 25313 23673 25347
rect 23673 25313 23707 25347
rect 23707 25313 23716 25347
rect 23664 25304 23716 25313
rect 24032 25304 24084 25356
rect 25044 25304 25096 25356
rect 19800 25236 19852 25288
rect 19984 25236 20036 25288
rect 22744 25236 22796 25288
rect 26148 25304 26200 25356
rect 27528 25347 27580 25356
rect 27528 25313 27537 25347
rect 27537 25313 27571 25347
rect 27571 25313 27580 25347
rect 27528 25304 27580 25313
rect 7104 25100 7156 25152
rect 26516 25168 26568 25220
rect 27252 25168 27304 25220
rect 23480 25143 23532 25152
rect 23480 25109 23489 25143
rect 23489 25109 23523 25143
rect 23523 25109 23532 25143
rect 23480 25100 23532 25109
rect 23756 25100 23808 25152
rect 28080 25100 28132 25152
rect 7896 24998 7948 25050
rect 7960 24998 8012 25050
rect 8024 24998 8076 25050
rect 8088 24998 8140 25050
rect 8152 24998 8204 25050
rect 14842 24998 14894 25050
rect 14906 24998 14958 25050
rect 14970 24998 15022 25050
rect 15034 24998 15086 25050
rect 15098 24998 15150 25050
rect 21788 24998 21840 25050
rect 21852 24998 21904 25050
rect 21916 24998 21968 25050
rect 21980 24998 22032 25050
rect 22044 24998 22096 25050
rect 28734 24998 28786 25050
rect 28798 24998 28850 25050
rect 28862 24998 28914 25050
rect 28926 24998 28978 25050
rect 28990 24998 29042 25050
rect 4160 24896 4212 24948
rect 7472 24939 7524 24948
rect 7472 24905 7481 24939
rect 7481 24905 7515 24939
rect 7515 24905 7524 24939
rect 7472 24896 7524 24905
rect 7748 24896 7800 24948
rect 23480 24896 23532 24948
rect 24032 24896 24084 24948
rect 2044 24828 2096 24880
rect 3976 24828 4028 24880
rect 9496 24828 9548 24880
rect 14280 24828 14332 24880
rect 23388 24828 23440 24880
rect 2964 24760 3016 24812
rect 12072 24760 12124 24812
rect 15660 24760 15712 24812
rect 17132 24803 17184 24812
rect 17132 24769 17166 24803
rect 17166 24769 17184 24803
rect 17132 24760 17184 24769
rect 18144 24760 18196 24812
rect 23572 24760 23624 24812
rect 25136 24803 25188 24812
rect 2872 24735 2924 24744
rect 2872 24701 2881 24735
rect 2881 24701 2915 24735
rect 2915 24701 2924 24735
rect 2872 24692 2924 24701
rect 7748 24692 7800 24744
rect 11796 24692 11848 24744
rect 12348 24735 12400 24744
rect 12348 24701 12357 24735
rect 12357 24701 12391 24735
rect 12391 24701 12400 24735
rect 12348 24692 12400 24701
rect 14740 24735 14792 24744
rect 14740 24701 14749 24735
rect 14749 24701 14783 24735
rect 14783 24701 14792 24735
rect 14740 24692 14792 24701
rect 15016 24692 15068 24744
rect 16856 24735 16908 24744
rect 16856 24701 16865 24735
rect 16865 24701 16899 24735
rect 16899 24701 16908 24735
rect 16856 24692 16908 24701
rect 12440 24624 12492 24676
rect 11704 24599 11756 24608
rect 11704 24565 11713 24599
rect 11713 24565 11747 24599
rect 11747 24565 11756 24599
rect 11704 24556 11756 24565
rect 12716 24556 12768 24608
rect 17500 24556 17552 24608
rect 22744 24692 22796 24744
rect 25136 24769 25145 24803
rect 25145 24769 25179 24803
rect 25179 24769 25188 24803
rect 25136 24760 25188 24769
rect 26148 24803 26200 24812
rect 26148 24769 26157 24803
rect 26157 24769 26191 24803
rect 26191 24769 26200 24803
rect 26148 24760 26200 24769
rect 27252 24692 27304 24744
rect 24676 24599 24728 24608
rect 24676 24565 24685 24599
rect 24685 24565 24719 24599
rect 24719 24565 24728 24599
rect 24676 24556 24728 24565
rect 25044 24599 25096 24608
rect 25044 24565 25053 24599
rect 25053 24565 25087 24599
rect 25087 24565 25096 24599
rect 25044 24556 25096 24565
rect 4423 24454 4475 24506
rect 4487 24454 4539 24506
rect 4551 24454 4603 24506
rect 4615 24454 4667 24506
rect 4679 24454 4731 24506
rect 11369 24454 11421 24506
rect 11433 24454 11485 24506
rect 11497 24454 11549 24506
rect 11561 24454 11613 24506
rect 11625 24454 11677 24506
rect 18315 24454 18367 24506
rect 18379 24454 18431 24506
rect 18443 24454 18495 24506
rect 18507 24454 18559 24506
rect 18571 24454 18623 24506
rect 25261 24454 25313 24506
rect 25325 24454 25377 24506
rect 25389 24454 25441 24506
rect 25453 24454 25505 24506
rect 25517 24454 25569 24506
rect 3148 24352 3200 24404
rect 11796 24395 11848 24404
rect 11796 24361 11805 24395
rect 11805 24361 11839 24395
rect 11839 24361 11848 24395
rect 11796 24352 11848 24361
rect 12716 24395 12768 24404
rect 12716 24361 12725 24395
rect 12725 24361 12759 24395
rect 12759 24361 12768 24395
rect 12716 24352 12768 24361
rect 15016 24352 15068 24404
rect 17132 24352 17184 24404
rect 2780 24148 2832 24200
rect 4068 24148 4120 24200
rect 5264 24216 5316 24268
rect 17500 24259 17552 24268
rect 17500 24225 17509 24259
rect 17509 24225 17543 24259
rect 17543 24225 17552 24259
rect 17500 24216 17552 24225
rect 17684 24259 17736 24268
rect 17684 24225 17693 24259
rect 17693 24225 17727 24259
rect 17727 24225 17736 24259
rect 17684 24216 17736 24225
rect 22468 24216 22520 24268
rect 23664 24216 23716 24268
rect 6368 24191 6420 24200
rect 6368 24157 6377 24191
rect 6377 24157 6411 24191
rect 6411 24157 6420 24191
rect 6368 24148 6420 24157
rect 9404 24148 9456 24200
rect 11704 24148 11756 24200
rect 12440 24191 12492 24200
rect 12440 24157 12449 24191
rect 12449 24157 12483 24191
rect 12483 24157 12492 24191
rect 12440 24148 12492 24157
rect 12532 24191 12584 24200
rect 12532 24157 12541 24191
rect 12541 24157 12575 24191
rect 12575 24157 12584 24191
rect 12532 24148 12584 24157
rect 16856 24148 16908 24200
rect 18144 24148 18196 24200
rect 19616 24191 19668 24200
rect 19616 24157 19625 24191
rect 19625 24157 19659 24191
rect 19659 24157 19668 24191
rect 19616 24148 19668 24157
rect 22376 24191 22428 24200
rect 22376 24157 22385 24191
rect 22385 24157 22419 24191
rect 22419 24157 22428 24191
rect 22376 24148 22428 24157
rect 27620 24148 27672 24200
rect 4252 24080 4304 24132
rect 11244 24080 11296 24132
rect 14372 24080 14424 24132
rect 3884 24012 3936 24064
rect 6828 24012 6880 24064
rect 12164 24012 12216 24064
rect 14280 24012 14332 24064
rect 20904 24080 20956 24132
rect 28172 24123 28224 24132
rect 28172 24089 28181 24123
rect 28181 24089 28215 24123
rect 28215 24089 28224 24123
rect 28172 24080 28224 24089
rect 18604 24055 18656 24064
rect 18604 24021 18613 24055
rect 18613 24021 18647 24055
rect 18647 24021 18656 24055
rect 18604 24012 18656 24021
rect 18880 24012 18932 24064
rect 22284 24012 22336 24064
rect 23480 24012 23532 24064
rect 7896 23910 7948 23962
rect 7960 23910 8012 23962
rect 8024 23910 8076 23962
rect 8088 23910 8140 23962
rect 8152 23910 8204 23962
rect 14842 23910 14894 23962
rect 14906 23910 14958 23962
rect 14970 23910 15022 23962
rect 15034 23910 15086 23962
rect 15098 23910 15150 23962
rect 21788 23910 21840 23962
rect 21852 23910 21904 23962
rect 21916 23910 21968 23962
rect 21980 23910 22032 23962
rect 22044 23910 22096 23962
rect 28734 23910 28786 23962
rect 28798 23910 28850 23962
rect 28862 23910 28914 23962
rect 28926 23910 28978 23962
rect 28990 23910 29042 23962
rect 2872 23851 2924 23860
rect 2872 23817 2881 23851
rect 2881 23817 2915 23851
rect 2915 23817 2924 23851
rect 2872 23808 2924 23817
rect 6368 23808 6420 23860
rect 7840 23808 7892 23860
rect 23480 23808 23532 23860
rect 6828 23783 6880 23792
rect 6828 23749 6837 23783
rect 6837 23749 6871 23783
rect 6871 23749 6880 23783
rect 6828 23740 6880 23749
rect 7288 23740 7340 23792
rect 18880 23783 18932 23792
rect 18880 23749 18889 23783
rect 18889 23749 18923 23783
rect 18923 23749 18932 23783
rect 18880 23740 18932 23749
rect 19432 23740 19484 23792
rect 22284 23783 22336 23792
rect 22284 23749 22318 23783
rect 22318 23749 22336 23783
rect 22284 23740 22336 23749
rect 26056 23740 26108 23792
rect 4344 23715 4396 23724
rect 4344 23681 4353 23715
rect 4353 23681 4387 23715
rect 4387 23681 4396 23715
rect 4344 23672 4396 23681
rect 14280 23672 14332 23724
rect 18604 23715 18656 23724
rect 18604 23681 18613 23715
rect 18613 23681 18647 23715
rect 18647 23681 18656 23715
rect 18604 23672 18656 23681
rect 20536 23672 20588 23724
rect 26148 23672 26200 23724
rect 27436 23715 27488 23724
rect 27436 23681 27445 23715
rect 27445 23681 27479 23715
rect 27479 23681 27488 23715
rect 27436 23672 27488 23681
rect 6552 23647 6604 23656
rect 6552 23613 6561 23647
rect 6561 23613 6595 23647
rect 6595 23613 6604 23647
rect 6552 23604 6604 23613
rect 14556 23647 14608 23656
rect 14556 23613 14565 23647
rect 14565 23613 14599 23647
rect 14599 23613 14608 23647
rect 14556 23604 14608 23613
rect 19616 23604 19668 23656
rect 27344 23647 27396 23656
rect 27344 23613 27353 23647
rect 27353 23613 27387 23647
rect 27387 23613 27396 23647
rect 27344 23604 27396 23613
rect 27988 23604 28040 23656
rect 26700 23468 26752 23520
rect 4423 23366 4475 23418
rect 4487 23366 4539 23418
rect 4551 23366 4603 23418
rect 4615 23366 4667 23418
rect 4679 23366 4731 23418
rect 11369 23366 11421 23418
rect 11433 23366 11485 23418
rect 11497 23366 11549 23418
rect 11561 23366 11613 23418
rect 11625 23366 11677 23418
rect 18315 23366 18367 23418
rect 18379 23366 18431 23418
rect 18443 23366 18495 23418
rect 18507 23366 18559 23418
rect 18571 23366 18623 23418
rect 25261 23366 25313 23418
rect 25325 23366 25377 23418
rect 25389 23366 25441 23418
rect 25453 23366 25505 23418
rect 25517 23366 25569 23418
rect 4068 23264 4120 23316
rect 12532 23264 12584 23316
rect 14372 23264 14424 23316
rect 25136 23307 25188 23316
rect 25136 23273 25145 23307
rect 25145 23273 25179 23307
rect 25179 23273 25188 23307
rect 25136 23264 25188 23273
rect 26148 23264 26200 23316
rect 2228 23060 2280 23112
rect 2780 23196 2832 23248
rect 23664 23196 23716 23248
rect 3056 23060 3108 23112
rect 3424 23103 3476 23112
rect 3424 23069 3433 23103
rect 3433 23069 3467 23103
rect 3467 23069 3476 23103
rect 3976 23103 4028 23112
rect 3424 23060 3476 23069
rect 3976 23069 3985 23103
rect 3985 23069 4019 23103
rect 4019 23069 4028 23103
rect 3976 23060 4028 23069
rect 5816 23060 5868 23112
rect 6644 23128 6696 23180
rect 7288 23171 7340 23180
rect 7288 23137 7297 23171
rect 7297 23137 7331 23171
rect 7331 23137 7340 23171
rect 7288 23128 7340 23137
rect 8208 23128 8260 23180
rect 9772 23128 9824 23180
rect 10508 23128 10560 23180
rect 6460 23060 6512 23112
rect 7840 23060 7892 23112
rect 12624 23128 12676 23180
rect 13176 23128 13228 23180
rect 14740 23171 14792 23180
rect 14740 23137 14749 23171
rect 14749 23137 14783 23171
rect 14783 23137 14792 23171
rect 14740 23128 14792 23137
rect 2780 22924 2832 22976
rect 4344 22924 4396 22976
rect 6368 22924 6420 22976
rect 6736 22924 6788 22976
rect 12808 23060 12860 23112
rect 14648 23060 14700 23112
rect 23572 23128 23624 23180
rect 15660 23103 15712 23112
rect 15660 23069 15669 23103
rect 15669 23069 15703 23103
rect 15703 23069 15712 23103
rect 15660 23060 15712 23069
rect 24032 23128 24084 23180
rect 26700 23171 26752 23180
rect 26700 23137 26709 23171
rect 26709 23137 26743 23171
rect 26743 23137 26752 23171
rect 26700 23128 26752 23137
rect 26240 23060 26292 23112
rect 26424 23103 26476 23112
rect 26424 23069 26433 23103
rect 26433 23069 26467 23103
rect 26467 23069 26476 23103
rect 26424 23060 26476 23069
rect 19800 22992 19852 23044
rect 22560 23035 22612 23044
rect 22560 23001 22569 23035
rect 22569 23001 22603 23035
rect 22603 23001 22612 23035
rect 22560 22992 22612 23001
rect 27988 22992 28040 23044
rect 12256 22967 12308 22976
rect 12256 22933 12265 22967
rect 12265 22933 12299 22967
rect 12299 22933 12308 22967
rect 12256 22924 12308 22933
rect 14096 22924 14148 22976
rect 14556 22924 14608 22976
rect 16212 22924 16264 22976
rect 7896 22822 7948 22874
rect 7960 22822 8012 22874
rect 8024 22822 8076 22874
rect 8088 22822 8140 22874
rect 8152 22822 8204 22874
rect 14842 22822 14894 22874
rect 14906 22822 14958 22874
rect 14970 22822 15022 22874
rect 15034 22822 15086 22874
rect 15098 22822 15150 22874
rect 21788 22822 21840 22874
rect 21852 22822 21904 22874
rect 21916 22822 21968 22874
rect 21980 22822 22032 22874
rect 22044 22822 22096 22874
rect 28734 22822 28786 22874
rect 28798 22822 28850 22874
rect 28862 22822 28914 22874
rect 28926 22822 28978 22874
rect 28990 22822 29042 22874
rect 4160 22720 4212 22772
rect 6552 22720 6604 22772
rect 8300 22720 8352 22772
rect 3424 22652 3476 22704
rect 3700 22584 3752 22636
rect 4252 22584 4304 22636
rect 6368 22584 6420 22636
rect 7104 22627 7156 22636
rect 7104 22593 7113 22627
rect 7113 22593 7147 22627
rect 7147 22593 7156 22627
rect 11060 22652 11112 22704
rect 12440 22652 12492 22704
rect 7104 22584 7156 22593
rect 7656 22584 7708 22636
rect 9404 22627 9456 22636
rect 9404 22593 9413 22627
rect 9413 22593 9447 22627
rect 9447 22593 9456 22627
rect 9404 22584 9456 22593
rect 9680 22627 9732 22636
rect 9680 22593 9714 22627
rect 9714 22593 9732 22627
rect 9680 22584 9732 22593
rect 11152 22584 11204 22636
rect 12256 22627 12308 22636
rect 12256 22593 12264 22627
rect 12264 22593 12298 22627
rect 12298 22593 12308 22627
rect 12256 22584 12308 22593
rect 16948 22720 17000 22772
rect 19432 22763 19484 22772
rect 19432 22729 19441 22763
rect 19441 22729 19475 22763
rect 19475 22729 19484 22763
rect 19432 22720 19484 22729
rect 22560 22720 22612 22772
rect 23388 22720 23440 22772
rect 26424 22720 26476 22772
rect 15292 22652 15344 22704
rect 2044 22516 2096 22568
rect 11244 22516 11296 22568
rect 16212 22627 16264 22636
rect 16212 22593 16221 22627
rect 16221 22593 16255 22627
rect 16255 22593 16264 22627
rect 16212 22584 16264 22593
rect 17776 22584 17828 22636
rect 19800 22627 19852 22636
rect 19800 22593 19809 22627
rect 19809 22593 19843 22627
rect 19843 22593 19852 22627
rect 19800 22584 19852 22593
rect 19892 22584 19944 22636
rect 22652 22627 22704 22636
rect 22652 22593 22661 22627
rect 22661 22593 22695 22627
rect 22695 22593 22704 22627
rect 22652 22584 22704 22593
rect 26240 22584 26292 22636
rect 27528 22584 27580 22636
rect 13360 22559 13412 22568
rect 13360 22525 13369 22559
rect 13369 22525 13403 22559
rect 13403 22525 13412 22559
rect 13360 22516 13412 22525
rect 14188 22559 14240 22568
rect 14188 22525 14197 22559
rect 14197 22525 14231 22559
rect 14231 22525 14240 22559
rect 14188 22516 14240 22525
rect 15936 22559 15988 22568
rect 15936 22525 15945 22559
rect 15945 22525 15979 22559
rect 15979 22525 15988 22559
rect 15936 22516 15988 22525
rect 17960 22559 18012 22568
rect 17960 22525 17969 22559
rect 17969 22525 18003 22559
rect 18003 22525 18012 22559
rect 17960 22516 18012 22525
rect 4804 22448 4856 22500
rect 17684 22448 17736 22500
rect 17868 22448 17920 22500
rect 4160 22380 4212 22432
rect 10968 22380 11020 22432
rect 11980 22380 12032 22432
rect 17500 22423 17552 22432
rect 17500 22389 17509 22423
rect 17509 22389 17543 22423
rect 17543 22389 17552 22423
rect 17500 22380 17552 22389
rect 27252 22423 27304 22432
rect 27252 22389 27261 22423
rect 27261 22389 27295 22423
rect 27295 22389 27304 22423
rect 27252 22380 27304 22389
rect 4423 22278 4475 22330
rect 4487 22278 4539 22330
rect 4551 22278 4603 22330
rect 4615 22278 4667 22330
rect 4679 22278 4731 22330
rect 11369 22278 11421 22330
rect 11433 22278 11485 22330
rect 11497 22278 11549 22330
rect 11561 22278 11613 22330
rect 11625 22278 11677 22330
rect 18315 22278 18367 22330
rect 18379 22278 18431 22330
rect 18443 22278 18495 22330
rect 18507 22278 18559 22330
rect 18571 22278 18623 22330
rect 25261 22278 25313 22330
rect 25325 22278 25377 22330
rect 25389 22278 25441 22330
rect 25453 22278 25505 22330
rect 25517 22278 25569 22330
rect 3424 22219 3476 22228
rect 3424 22185 3433 22219
rect 3433 22185 3467 22219
rect 3467 22185 3476 22219
rect 3424 22176 3476 22185
rect 7656 22219 7708 22228
rect 7656 22185 7665 22219
rect 7665 22185 7699 22219
rect 7699 22185 7708 22219
rect 7656 22176 7708 22185
rect 17960 22176 18012 22228
rect 24032 22219 24084 22228
rect 7748 22108 7800 22160
rect 6460 22040 6512 22092
rect 8208 22040 8260 22092
rect 10416 22108 10468 22160
rect 12440 22083 12492 22092
rect 12440 22049 12449 22083
rect 12449 22049 12483 22083
rect 12483 22049 12492 22083
rect 15292 22083 15344 22092
rect 12440 22040 12492 22049
rect 15292 22049 15301 22083
rect 15301 22049 15335 22083
rect 15335 22049 15344 22083
rect 15292 22040 15344 22049
rect 24032 22185 24041 22219
rect 24041 22185 24075 22219
rect 24075 22185 24084 22219
rect 24032 22176 24084 22185
rect 27252 22176 27304 22228
rect 19984 22083 20036 22092
rect 19984 22049 19993 22083
rect 19993 22049 20027 22083
rect 20027 22049 20036 22083
rect 19984 22040 20036 22049
rect 27528 22040 27580 22092
rect 2044 22015 2096 22024
rect 2044 21981 2053 22015
rect 2053 21981 2087 22015
rect 2087 21981 2096 22015
rect 2044 21972 2096 21981
rect 2780 21972 2832 22024
rect 3056 21972 3108 22024
rect 4068 21972 4120 22024
rect 4252 21972 4304 22024
rect 5540 21972 5592 22024
rect 5816 21972 5868 22024
rect 10416 21972 10468 22024
rect 12256 21972 12308 22024
rect 12624 22015 12676 22024
rect 12624 21981 12633 22015
rect 12633 21981 12667 22015
rect 12667 21981 12676 22015
rect 12624 21972 12676 21981
rect 12808 22015 12860 22024
rect 12808 21981 12817 22015
rect 12817 21981 12851 22015
rect 12851 21981 12860 22015
rect 12808 21972 12860 21981
rect 13268 22015 13320 22024
rect 13268 21981 13277 22015
rect 13277 21981 13311 22015
rect 13311 21981 13320 22015
rect 13268 21972 13320 21981
rect 6368 21947 6420 21956
rect 6368 21913 6377 21947
rect 6377 21913 6411 21947
rect 6411 21913 6420 21947
rect 6368 21904 6420 21913
rect 9588 21904 9640 21956
rect 12532 21904 12584 21956
rect 13544 21947 13596 21956
rect 13544 21913 13553 21947
rect 13553 21913 13587 21947
rect 13587 21913 13596 21947
rect 13544 21904 13596 21913
rect 9404 21836 9456 21888
rect 9864 21836 9916 21888
rect 14464 21972 14516 22024
rect 16856 21972 16908 22024
rect 17316 21972 17368 22024
rect 17500 22015 17552 22024
rect 17500 21981 17534 22015
rect 17534 21981 17552 22015
rect 19616 22015 19668 22024
rect 17500 21972 17552 21981
rect 19616 21981 19625 22015
rect 19625 21981 19659 22015
rect 19659 21981 19668 22015
rect 19616 21972 19668 21981
rect 22744 21972 22796 22024
rect 26240 22015 26292 22024
rect 26240 21981 26249 22015
rect 26249 21981 26283 22015
rect 26283 21981 26292 22015
rect 26240 21972 26292 21981
rect 23204 21904 23256 21956
rect 28264 21904 28316 21956
rect 7896 21734 7948 21786
rect 7960 21734 8012 21786
rect 8024 21734 8076 21786
rect 8088 21734 8140 21786
rect 8152 21734 8204 21786
rect 14842 21734 14894 21786
rect 14906 21734 14958 21786
rect 14970 21734 15022 21786
rect 15034 21734 15086 21786
rect 15098 21734 15150 21786
rect 21788 21734 21840 21786
rect 21852 21734 21904 21786
rect 21916 21734 21968 21786
rect 21980 21734 22032 21786
rect 22044 21734 22096 21786
rect 28734 21734 28786 21786
rect 28798 21734 28850 21786
rect 28862 21734 28914 21786
rect 28926 21734 28978 21786
rect 28990 21734 29042 21786
rect 3700 21675 3752 21684
rect 2228 21564 2280 21616
rect 3148 21564 3200 21616
rect 3700 21641 3709 21675
rect 3709 21641 3743 21675
rect 3743 21641 3752 21675
rect 3700 21632 3752 21641
rect 9680 21632 9732 21684
rect 10140 21632 10192 21684
rect 11152 21675 11204 21684
rect 11152 21641 11161 21675
rect 11161 21641 11195 21675
rect 11195 21641 11204 21675
rect 11152 21632 11204 21641
rect 12808 21632 12860 21684
rect 13452 21632 13504 21684
rect 15936 21632 15988 21684
rect 4804 21564 4856 21616
rect 10876 21564 10928 21616
rect 3884 21539 3936 21548
rect 3884 21505 3893 21539
rect 3893 21505 3927 21539
rect 3927 21505 3936 21539
rect 3884 21496 3936 21505
rect 4160 21539 4212 21548
rect 4160 21505 4169 21539
rect 4169 21505 4203 21539
rect 4203 21505 4212 21539
rect 4160 21496 4212 21505
rect 6736 21539 6788 21548
rect 6736 21505 6745 21539
rect 6745 21505 6779 21539
rect 6779 21505 6788 21539
rect 6736 21496 6788 21505
rect 10140 21539 10192 21548
rect 10140 21505 10149 21539
rect 10149 21505 10183 21539
rect 10183 21505 10192 21539
rect 10140 21496 10192 21505
rect 10692 21496 10744 21548
rect 10968 21539 11020 21548
rect 10968 21505 10977 21539
rect 10977 21505 11011 21539
rect 11011 21505 11020 21539
rect 10968 21496 11020 21505
rect 13544 21564 13596 21616
rect 21548 21632 21600 21684
rect 22744 21632 22796 21684
rect 23204 21675 23256 21684
rect 23204 21641 23213 21675
rect 23213 21641 23247 21675
rect 23247 21641 23256 21675
rect 23204 21632 23256 21641
rect 24032 21632 24084 21684
rect 26240 21632 26292 21684
rect 28264 21675 28316 21684
rect 28264 21641 28273 21675
rect 28273 21641 28307 21675
rect 28307 21641 28316 21675
rect 28264 21632 28316 21641
rect 12992 21496 13044 21548
rect 14188 21496 14240 21548
rect 17316 21564 17368 21616
rect 17500 21564 17552 21616
rect 23480 21564 23532 21616
rect 23756 21564 23808 21616
rect 17224 21539 17276 21548
rect 17224 21505 17258 21539
rect 17258 21505 17276 21539
rect 17224 21496 17276 21505
rect 19708 21496 19760 21548
rect 21640 21496 21692 21548
rect 22836 21496 22888 21548
rect 26424 21539 26476 21548
rect 26424 21505 26433 21539
rect 26433 21505 26467 21539
rect 26467 21505 26476 21539
rect 26424 21496 26476 21505
rect 27436 21539 27488 21548
rect 27436 21505 27445 21539
rect 27445 21505 27479 21539
rect 27479 21505 27488 21539
rect 27436 21496 27488 21505
rect 3240 21471 3292 21480
rect 3240 21437 3249 21471
rect 3249 21437 3283 21471
rect 3283 21437 3292 21471
rect 3240 21428 3292 21437
rect 4068 21471 4120 21480
rect 4068 21437 4077 21471
rect 4077 21437 4111 21471
rect 4111 21437 4120 21471
rect 4068 21428 4120 21437
rect 10416 21471 10468 21480
rect 10416 21437 10425 21471
rect 10425 21437 10459 21471
rect 10459 21437 10468 21471
rect 10416 21428 10468 21437
rect 12348 21471 12400 21480
rect 12348 21437 12357 21471
rect 12357 21437 12391 21471
rect 12391 21437 12400 21471
rect 12348 21428 12400 21437
rect 14740 21471 14792 21480
rect 14740 21437 14749 21471
rect 14749 21437 14783 21471
rect 14783 21437 14792 21471
rect 14740 21428 14792 21437
rect 17960 21360 18012 21412
rect 2780 21335 2832 21344
rect 2780 21301 2789 21335
rect 2789 21301 2823 21335
rect 2823 21301 2832 21335
rect 2780 21292 2832 21301
rect 4896 21292 4948 21344
rect 5632 21292 5684 21344
rect 12256 21292 12308 21344
rect 12716 21292 12768 21344
rect 13820 21292 13872 21344
rect 21824 21292 21876 21344
rect 22284 21292 22336 21344
rect 23572 21292 23624 21344
rect 26240 21428 26292 21480
rect 27344 21471 27396 21480
rect 27344 21437 27353 21471
rect 27353 21437 27387 21471
rect 27387 21437 27396 21471
rect 27344 21428 27396 21437
rect 24768 21360 24820 21412
rect 25136 21292 25188 21344
rect 4423 21190 4475 21242
rect 4487 21190 4539 21242
rect 4551 21190 4603 21242
rect 4615 21190 4667 21242
rect 4679 21190 4731 21242
rect 11369 21190 11421 21242
rect 11433 21190 11485 21242
rect 11497 21190 11549 21242
rect 11561 21190 11613 21242
rect 11625 21190 11677 21242
rect 18315 21190 18367 21242
rect 18379 21190 18431 21242
rect 18443 21190 18495 21242
rect 18507 21190 18559 21242
rect 18571 21190 18623 21242
rect 25261 21190 25313 21242
rect 25325 21190 25377 21242
rect 25389 21190 25441 21242
rect 25453 21190 25505 21242
rect 25517 21190 25569 21242
rect 6736 21088 6788 21140
rect 9404 21088 9456 21140
rect 12992 21131 13044 21140
rect 12992 21097 13001 21131
rect 13001 21097 13035 21131
rect 13035 21097 13044 21131
rect 12992 21088 13044 21097
rect 13360 21088 13412 21140
rect 15936 21088 15988 21140
rect 17224 21088 17276 21140
rect 19984 21088 20036 21140
rect 16764 21020 16816 21072
rect 17132 21020 17184 21072
rect 5724 20952 5776 21004
rect 7748 20952 7800 21004
rect 9680 20952 9732 21004
rect 13452 20995 13504 21004
rect 4344 20884 4396 20936
rect 7656 20884 7708 20936
rect 10140 20884 10192 20936
rect 13452 20961 13461 20995
rect 13461 20961 13495 20995
rect 13495 20961 13504 20995
rect 13452 20952 13504 20961
rect 14648 20952 14700 21004
rect 17868 20995 17920 21004
rect 17868 20961 17877 20995
rect 17877 20961 17911 20995
rect 17911 20961 17920 20995
rect 17868 20952 17920 20961
rect 23664 20995 23716 21004
rect 23664 20961 23673 20995
rect 23673 20961 23707 20995
rect 23707 20961 23716 20995
rect 23664 20952 23716 20961
rect 5632 20859 5684 20868
rect 5632 20825 5641 20859
rect 5641 20825 5675 20859
rect 5675 20825 5684 20859
rect 5632 20816 5684 20825
rect 6368 20816 6420 20868
rect 9588 20816 9640 20868
rect 14464 20884 14516 20936
rect 17132 20884 17184 20936
rect 17960 20884 18012 20936
rect 20076 20884 20128 20936
rect 20536 20884 20588 20936
rect 21824 20927 21876 20936
rect 21824 20893 21833 20927
rect 21833 20893 21867 20927
rect 21867 20893 21876 20927
rect 21824 20884 21876 20893
rect 14556 20816 14608 20868
rect 20444 20816 20496 20868
rect 21272 20816 21324 20868
rect 22100 20927 22152 20936
rect 22100 20893 22109 20927
rect 22109 20893 22143 20927
rect 22143 20893 22152 20927
rect 22100 20884 22152 20893
rect 22284 20927 22336 20936
rect 22284 20893 22298 20927
rect 22298 20893 22332 20927
rect 22332 20893 22336 20927
rect 23572 20927 23624 20936
rect 22284 20884 22336 20893
rect 23572 20893 23581 20927
rect 23581 20893 23615 20927
rect 23615 20893 23624 20927
rect 23572 20884 23624 20893
rect 23848 20927 23900 20936
rect 23848 20893 23857 20927
rect 23857 20893 23891 20927
rect 23891 20893 23900 20927
rect 23848 20884 23900 20893
rect 24676 20952 24728 21004
rect 27896 20927 27948 20936
rect 22376 20816 22428 20868
rect 27896 20893 27905 20927
rect 27905 20893 27939 20927
rect 27939 20893 27948 20927
rect 27896 20884 27948 20893
rect 28172 20859 28224 20868
rect 2044 20791 2096 20800
rect 2044 20757 2053 20791
rect 2053 20757 2087 20791
rect 2087 20757 2096 20791
rect 2044 20748 2096 20757
rect 13360 20791 13412 20800
rect 13360 20757 13369 20791
rect 13369 20757 13403 20791
rect 13403 20757 13412 20791
rect 13360 20748 13412 20757
rect 14280 20791 14332 20800
rect 14280 20757 14289 20791
rect 14289 20757 14323 20791
rect 14323 20757 14332 20791
rect 14280 20748 14332 20757
rect 14740 20791 14792 20800
rect 14740 20757 14749 20791
rect 14749 20757 14783 20791
rect 14783 20757 14792 20791
rect 14740 20748 14792 20757
rect 21640 20748 21692 20800
rect 28172 20825 28181 20859
rect 28181 20825 28215 20859
rect 28215 20825 28224 20859
rect 28172 20816 28224 20825
rect 24860 20791 24912 20800
rect 24860 20757 24869 20791
rect 24869 20757 24903 20791
rect 24903 20757 24912 20791
rect 24860 20748 24912 20757
rect 7896 20646 7948 20698
rect 7960 20646 8012 20698
rect 8024 20646 8076 20698
rect 8088 20646 8140 20698
rect 8152 20646 8204 20698
rect 14842 20646 14894 20698
rect 14906 20646 14958 20698
rect 14970 20646 15022 20698
rect 15034 20646 15086 20698
rect 15098 20646 15150 20698
rect 21788 20646 21840 20698
rect 21852 20646 21904 20698
rect 21916 20646 21968 20698
rect 21980 20646 22032 20698
rect 22044 20646 22096 20698
rect 28734 20646 28786 20698
rect 28798 20646 28850 20698
rect 28862 20646 28914 20698
rect 28926 20646 28978 20698
rect 28990 20646 29042 20698
rect 3240 20544 3292 20596
rect 2780 20476 2832 20528
rect 5724 20544 5776 20596
rect 10140 20544 10192 20596
rect 11060 20587 11112 20596
rect 11060 20553 11069 20587
rect 11069 20553 11103 20587
rect 11103 20553 11112 20587
rect 11060 20544 11112 20553
rect 14740 20544 14792 20596
rect 20444 20587 20496 20596
rect 20444 20553 20453 20587
rect 20453 20553 20487 20587
rect 20487 20553 20496 20587
rect 20444 20544 20496 20553
rect 22376 20587 22428 20596
rect 22376 20553 22385 20587
rect 22385 20553 22419 20587
rect 22419 20553 22428 20587
rect 22376 20544 22428 20553
rect 4252 20408 4304 20460
rect 13820 20476 13872 20528
rect 14280 20476 14332 20528
rect 17132 20519 17184 20528
rect 17132 20485 17166 20519
rect 17166 20485 17184 20519
rect 17132 20476 17184 20485
rect 17776 20476 17828 20528
rect 4896 20408 4948 20460
rect 6000 20408 6052 20460
rect 7656 20408 7708 20460
rect 9864 20451 9916 20460
rect 9864 20417 9873 20451
rect 9873 20417 9907 20451
rect 9907 20417 9916 20451
rect 9864 20408 9916 20417
rect 10692 20451 10744 20460
rect 10692 20417 10701 20451
rect 10701 20417 10735 20451
rect 10735 20417 10744 20451
rect 10692 20408 10744 20417
rect 10876 20451 10928 20460
rect 10876 20417 10885 20451
rect 10885 20417 10919 20451
rect 10919 20417 10928 20451
rect 10876 20408 10928 20417
rect 11980 20451 12032 20460
rect 2044 20383 2096 20392
rect 2044 20349 2053 20383
rect 2053 20349 2087 20383
rect 2087 20349 2096 20383
rect 2044 20340 2096 20349
rect 3240 20340 3292 20392
rect 7104 20340 7156 20392
rect 7748 20340 7800 20392
rect 9404 20340 9456 20392
rect 9772 20383 9824 20392
rect 9772 20349 9781 20383
rect 9781 20349 9815 20383
rect 9815 20349 9824 20383
rect 9772 20340 9824 20349
rect 11980 20417 11989 20451
rect 11989 20417 12023 20451
rect 12023 20417 12032 20451
rect 11980 20408 12032 20417
rect 12164 20451 12216 20460
rect 12164 20417 12173 20451
rect 12173 20417 12207 20451
rect 12207 20417 12216 20451
rect 12164 20408 12216 20417
rect 13544 20408 13596 20460
rect 21640 20476 21692 20528
rect 22836 20476 22888 20528
rect 23388 20519 23440 20528
rect 23388 20485 23397 20519
rect 23397 20485 23431 20519
rect 23431 20485 23440 20519
rect 23388 20476 23440 20485
rect 24952 20408 25004 20460
rect 26424 20408 26476 20460
rect 27344 20451 27396 20460
rect 27344 20417 27353 20451
rect 27353 20417 27387 20451
rect 27387 20417 27396 20451
rect 27344 20408 27396 20417
rect 13636 20340 13688 20392
rect 16856 20383 16908 20392
rect 16856 20349 16865 20383
rect 16865 20349 16899 20383
rect 16899 20349 16908 20383
rect 16856 20340 16908 20349
rect 13176 20272 13228 20324
rect 3148 20204 3200 20256
rect 7564 20204 7616 20256
rect 9680 20247 9732 20256
rect 9680 20213 9689 20247
rect 9689 20213 9723 20247
rect 9723 20213 9732 20247
rect 9680 20204 9732 20213
rect 16764 20204 16816 20256
rect 22468 20340 22520 20392
rect 26240 20340 26292 20392
rect 27620 20272 27672 20324
rect 26792 20204 26844 20256
rect 4423 20102 4475 20154
rect 4487 20102 4539 20154
rect 4551 20102 4603 20154
rect 4615 20102 4667 20154
rect 4679 20102 4731 20154
rect 11369 20102 11421 20154
rect 11433 20102 11485 20154
rect 11497 20102 11549 20154
rect 11561 20102 11613 20154
rect 11625 20102 11677 20154
rect 18315 20102 18367 20154
rect 18379 20102 18431 20154
rect 18443 20102 18495 20154
rect 18507 20102 18559 20154
rect 18571 20102 18623 20154
rect 25261 20102 25313 20154
rect 25325 20102 25377 20154
rect 25389 20102 25441 20154
rect 25453 20102 25505 20154
rect 25517 20102 25569 20154
rect 7656 20000 7708 20052
rect 9864 20000 9916 20052
rect 10508 20043 10560 20052
rect 10508 20009 10517 20043
rect 10517 20009 10551 20043
rect 10551 20009 10560 20043
rect 10508 20000 10560 20009
rect 12164 20000 12216 20052
rect 17868 20000 17920 20052
rect 20076 20043 20128 20052
rect 20076 20009 20085 20043
rect 20085 20009 20119 20043
rect 20119 20009 20128 20043
rect 20076 20000 20128 20009
rect 21272 20043 21324 20052
rect 21272 20009 21281 20043
rect 21281 20009 21315 20043
rect 21315 20009 21324 20043
rect 21272 20000 21324 20009
rect 27344 20000 27396 20052
rect 9772 19864 9824 19916
rect 2044 19839 2096 19848
rect 2044 19805 2053 19839
rect 2053 19805 2087 19839
rect 2087 19805 2096 19839
rect 2044 19796 2096 19805
rect 2780 19728 2832 19780
rect 6644 19796 6696 19848
rect 9312 19839 9364 19848
rect 9312 19805 9321 19839
rect 9321 19805 9355 19839
rect 9355 19805 9364 19839
rect 9312 19796 9364 19805
rect 10600 19796 10652 19848
rect 12348 19864 12400 19916
rect 12716 19864 12768 19916
rect 14556 19907 14608 19916
rect 14556 19873 14565 19907
rect 14565 19873 14599 19907
rect 14599 19873 14608 19907
rect 14556 19864 14608 19873
rect 16764 19907 16816 19916
rect 16764 19873 16773 19907
rect 16773 19873 16807 19907
rect 16807 19873 16816 19907
rect 16764 19864 16816 19873
rect 12992 19839 13044 19848
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 12992 19796 13044 19805
rect 16028 19796 16080 19848
rect 16948 19839 17000 19848
rect 5908 19728 5960 19780
rect 7472 19728 7524 19780
rect 11612 19771 11664 19780
rect 11612 19737 11630 19771
rect 11630 19737 11664 19771
rect 11612 19728 11664 19737
rect 16488 19728 16540 19780
rect 4344 19660 4396 19712
rect 13360 19660 13412 19712
rect 16948 19805 16957 19839
rect 16957 19805 16991 19839
rect 16991 19805 17000 19839
rect 16948 19796 17000 19805
rect 22652 19907 22704 19916
rect 22652 19873 22661 19907
rect 22661 19873 22695 19907
rect 22695 19873 22704 19907
rect 22652 19864 22704 19873
rect 24768 19864 24820 19916
rect 25136 19907 25188 19916
rect 25136 19873 25145 19907
rect 25145 19873 25179 19907
rect 25179 19873 25188 19907
rect 26792 19907 26844 19916
rect 25136 19864 25188 19873
rect 26792 19873 26801 19907
rect 26801 19873 26835 19907
rect 26835 19873 26844 19907
rect 26792 19864 26844 19873
rect 24952 19839 25004 19848
rect 24952 19805 24961 19839
rect 24961 19805 24995 19839
rect 24995 19805 25004 19839
rect 24952 19796 25004 19805
rect 19616 19728 19668 19780
rect 20904 19771 20956 19780
rect 20904 19737 20913 19771
rect 20913 19737 20947 19771
rect 20947 19737 20956 19771
rect 20904 19728 20956 19737
rect 22284 19728 22336 19780
rect 17040 19660 17092 19712
rect 26332 19728 26384 19780
rect 28080 19728 28132 19780
rect 7896 19558 7948 19610
rect 7960 19558 8012 19610
rect 8024 19558 8076 19610
rect 8088 19558 8140 19610
rect 8152 19558 8204 19610
rect 14842 19558 14894 19610
rect 14906 19558 14958 19610
rect 14970 19558 15022 19610
rect 15034 19558 15086 19610
rect 15098 19558 15150 19610
rect 21788 19558 21840 19610
rect 21852 19558 21904 19610
rect 21916 19558 21968 19610
rect 21980 19558 22032 19610
rect 22044 19558 22096 19610
rect 28734 19558 28786 19610
rect 28798 19558 28850 19610
rect 28862 19558 28914 19610
rect 28926 19558 28978 19610
rect 28990 19558 29042 19610
rect 3148 19456 3200 19508
rect 5908 19499 5960 19508
rect 4344 19431 4396 19440
rect 4344 19397 4353 19431
rect 4353 19397 4387 19431
rect 4387 19397 4396 19431
rect 4344 19388 4396 19397
rect 2780 19295 2832 19304
rect 2780 19261 2789 19295
rect 2789 19261 2823 19295
rect 2823 19261 2832 19295
rect 3148 19295 3200 19304
rect 2780 19252 2832 19261
rect 3148 19261 3157 19295
rect 3157 19261 3191 19295
rect 3191 19261 3200 19295
rect 3148 19252 3200 19261
rect 3240 19295 3292 19304
rect 3240 19261 3249 19295
rect 3249 19261 3283 19295
rect 3283 19261 3292 19295
rect 4896 19363 4948 19372
rect 4896 19329 4905 19363
rect 4905 19329 4939 19363
rect 4939 19329 4948 19363
rect 5908 19465 5917 19499
rect 5917 19465 5951 19499
rect 5951 19465 5960 19499
rect 5908 19456 5960 19465
rect 6644 19499 6696 19508
rect 6644 19465 6653 19499
rect 6653 19465 6687 19499
rect 6687 19465 6696 19499
rect 6644 19456 6696 19465
rect 7748 19456 7800 19508
rect 9496 19499 9548 19508
rect 9496 19465 9505 19499
rect 9505 19465 9539 19499
rect 9539 19465 9548 19499
rect 9496 19456 9548 19465
rect 11612 19456 11664 19508
rect 4896 19320 4948 19329
rect 7104 19388 7156 19440
rect 7564 19388 7616 19440
rect 7656 19388 7708 19440
rect 13268 19456 13320 19508
rect 16304 19456 16356 19508
rect 16856 19499 16908 19508
rect 16856 19465 16865 19499
rect 16865 19465 16899 19499
rect 16899 19465 16908 19499
rect 16856 19456 16908 19465
rect 20904 19456 20956 19508
rect 22192 19499 22244 19508
rect 12164 19431 12216 19440
rect 6000 19363 6052 19372
rect 6000 19329 6009 19363
rect 6009 19329 6043 19363
rect 6043 19329 6052 19363
rect 6000 19320 6052 19329
rect 8300 19320 8352 19372
rect 9312 19320 9364 19372
rect 9772 19320 9824 19372
rect 12164 19397 12173 19431
rect 12173 19397 12207 19431
rect 12207 19397 12216 19431
rect 12164 19388 12216 19397
rect 16580 19388 16632 19440
rect 17776 19388 17828 19440
rect 17960 19388 18012 19440
rect 12072 19363 12124 19372
rect 12072 19329 12081 19363
rect 12081 19329 12115 19363
rect 12115 19329 12124 19363
rect 12072 19320 12124 19329
rect 12992 19320 13044 19372
rect 13268 19363 13320 19372
rect 3240 19252 3292 19261
rect 7104 19252 7156 19304
rect 9496 19252 9548 19304
rect 13268 19329 13277 19363
rect 13277 19329 13311 19363
rect 13311 19329 13320 19363
rect 13268 19320 13320 19329
rect 14188 19363 14240 19372
rect 14188 19329 14197 19363
rect 14197 19329 14231 19363
rect 14231 19329 14240 19363
rect 14188 19320 14240 19329
rect 16028 19363 16080 19372
rect 16028 19329 16037 19363
rect 16037 19329 16071 19363
rect 16071 19329 16080 19363
rect 16028 19320 16080 19329
rect 17040 19363 17092 19372
rect 17040 19329 17049 19363
rect 17049 19329 17083 19363
rect 17083 19329 17092 19363
rect 17040 19320 17092 19329
rect 20076 19388 20128 19440
rect 22192 19465 22201 19499
rect 22201 19465 22235 19499
rect 22235 19465 22244 19499
rect 22192 19456 22244 19465
rect 28080 19456 28132 19508
rect 21732 19388 21784 19440
rect 21272 19320 21324 19372
rect 22192 19363 22244 19372
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 22652 19363 22704 19372
rect 22652 19329 22661 19363
rect 22661 19329 22695 19363
rect 22695 19329 22704 19363
rect 22652 19320 22704 19329
rect 22928 19363 22980 19372
rect 22928 19329 22962 19363
rect 22962 19329 22980 19363
rect 22928 19320 22980 19329
rect 26332 19320 26384 19372
rect 27436 19363 27488 19372
rect 27436 19329 27445 19363
rect 27445 19329 27479 19363
rect 27479 19329 27488 19363
rect 27436 19320 27488 19329
rect 13544 19252 13596 19304
rect 14648 19252 14700 19304
rect 15200 19252 15252 19304
rect 17500 19252 17552 19304
rect 19616 19252 19668 19304
rect 23848 19252 23900 19304
rect 10600 19184 10652 19236
rect 13636 19184 13688 19236
rect 4252 19116 4304 19168
rect 5080 19116 5132 19168
rect 7564 19116 7616 19168
rect 9220 19116 9272 19168
rect 18236 19116 18288 19168
rect 19892 19116 19944 19168
rect 21180 19116 21232 19168
rect 22560 19184 22612 19236
rect 24032 19227 24084 19236
rect 24032 19193 24041 19227
rect 24041 19193 24075 19227
rect 24075 19193 24084 19227
rect 26240 19252 26292 19304
rect 24032 19184 24084 19193
rect 25964 19116 26016 19168
rect 4423 19014 4475 19066
rect 4487 19014 4539 19066
rect 4551 19014 4603 19066
rect 4615 19014 4667 19066
rect 4679 19014 4731 19066
rect 11369 19014 11421 19066
rect 11433 19014 11485 19066
rect 11497 19014 11549 19066
rect 11561 19014 11613 19066
rect 11625 19014 11677 19066
rect 18315 19014 18367 19066
rect 18379 19014 18431 19066
rect 18443 19014 18495 19066
rect 18507 19014 18559 19066
rect 18571 19014 18623 19066
rect 25261 19014 25313 19066
rect 25325 19014 25377 19066
rect 25389 19014 25441 19066
rect 25453 19014 25505 19066
rect 25517 19014 25569 19066
rect 9772 18912 9824 18964
rect 12532 18912 12584 18964
rect 21272 18955 21324 18964
rect 21272 18921 21281 18955
rect 21281 18921 21315 18955
rect 21315 18921 21324 18955
rect 21272 18912 21324 18921
rect 22928 18955 22980 18964
rect 22928 18921 22937 18955
rect 22937 18921 22971 18955
rect 22971 18921 22980 18955
rect 22928 18912 22980 18921
rect 26332 18912 26384 18964
rect 5540 18844 5592 18896
rect 2044 18776 2096 18828
rect 2872 18708 2924 18760
rect 5908 18819 5960 18828
rect 5908 18785 5917 18819
rect 5917 18785 5951 18819
rect 5951 18785 5960 18819
rect 5908 18776 5960 18785
rect 7472 18776 7524 18828
rect 13452 18819 13504 18828
rect 13452 18785 13478 18819
rect 13478 18785 13504 18819
rect 21180 18844 21232 18896
rect 21732 18819 21784 18828
rect 13452 18776 13504 18785
rect 5816 18708 5868 18760
rect 4344 18683 4396 18692
rect 4344 18649 4353 18683
rect 4353 18649 4387 18683
rect 4387 18649 4396 18683
rect 4344 18640 4396 18649
rect 9220 18708 9272 18760
rect 13544 18708 13596 18760
rect 14740 18708 14792 18760
rect 15292 18708 15344 18760
rect 21732 18785 21741 18819
rect 21741 18785 21775 18819
rect 21775 18785 21784 18819
rect 21732 18776 21784 18785
rect 22192 18844 22244 18896
rect 10600 18640 10652 18692
rect 13176 18683 13228 18692
rect 13176 18649 13185 18683
rect 13185 18649 13219 18683
rect 13219 18649 13228 18683
rect 13176 18640 13228 18649
rect 14280 18640 14332 18692
rect 13636 18572 13688 18624
rect 17408 18708 17460 18760
rect 18236 18751 18288 18760
rect 18236 18717 18245 18751
rect 18245 18717 18279 18751
rect 18279 18717 18288 18751
rect 18236 18708 18288 18717
rect 19800 18708 19852 18760
rect 19892 18751 19944 18760
rect 19892 18717 19901 18751
rect 19901 18717 19935 18751
rect 19935 18717 19944 18751
rect 20812 18751 20864 18760
rect 19892 18708 19944 18717
rect 20812 18717 20821 18751
rect 20821 18717 20855 18751
rect 20855 18717 20864 18751
rect 20812 18708 20864 18717
rect 24032 18708 24084 18760
rect 25964 18819 26016 18828
rect 25964 18785 25973 18819
rect 25973 18785 26007 18819
rect 26007 18785 26016 18819
rect 25964 18776 26016 18785
rect 18880 18615 18932 18624
rect 18880 18581 18889 18615
rect 18889 18581 18923 18615
rect 18923 18581 18932 18615
rect 18880 18572 18932 18581
rect 25136 18640 25188 18692
rect 26608 18640 26660 18692
rect 20260 18572 20312 18624
rect 21640 18615 21692 18624
rect 21640 18581 21649 18615
rect 21649 18581 21683 18615
rect 21683 18581 21692 18615
rect 21640 18572 21692 18581
rect 23020 18572 23072 18624
rect 7896 18470 7948 18522
rect 7960 18470 8012 18522
rect 8024 18470 8076 18522
rect 8088 18470 8140 18522
rect 8152 18470 8204 18522
rect 14842 18470 14894 18522
rect 14906 18470 14958 18522
rect 14970 18470 15022 18522
rect 15034 18470 15086 18522
rect 15098 18470 15150 18522
rect 21788 18470 21840 18522
rect 21852 18470 21904 18522
rect 21916 18470 21968 18522
rect 21980 18470 22032 18522
rect 22044 18470 22096 18522
rect 28734 18470 28786 18522
rect 28798 18470 28850 18522
rect 28862 18470 28914 18522
rect 28926 18470 28978 18522
rect 28990 18470 29042 18522
rect 14740 18368 14792 18420
rect 17408 18411 17460 18420
rect 17408 18377 17417 18411
rect 17417 18377 17451 18411
rect 17451 18377 17460 18411
rect 17408 18368 17460 18377
rect 19984 18368 20036 18420
rect 22192 18368 22244 18420
rect 26608 18411 26660 18420
rect 26608 18377 26617 18411
rect 26617 18377 26651 18411
rect 26651 18377 26660 18411
rect 26608 18368 26660 18377
rect 2872 18343 2924 18352
rect 2872 18309 2881 18343
rect 2881 18309 2915 18343
rect 2915 18309 2924 18343
rect 2872 18300 2924 18309
rect 5816 18300 5868 18352
rect 9588 18343 9640 18352
rect 9588 18309 9597 18343
rect 9597 18309 9631 18343
rect 9631 18309 9640 18343
rect 9588 18300 9640 18309
rect 17500 18300 17552 18352
rect 18880 18300 18932 18352
rect 20260 18300 20312 18352
rect 24676 18300 24728 18352
rect 3976 18232 4028 18284
rect 6736 18275 6788 18284
rect 6736 18241 6745 18275
rect 6745 18241 6779 18275
rect 6779 18241 6788 18275
rect 6736 18232 6788 18241
rect 12808 18232 12860 18284
rect 13084 18275 13136 18284
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 13728 18232 13780 18284
rect 14648 18232 14700 18284
rect 13820 18164 13872 18216
rect 14280 18164 14332 18216
rect 25136 18232 25188 18284
rect 25780 18275 25832 18284
rect 25780 18241 25789 18275
rect 25789 18241 25823 18275
rect 25823 18241 25832 18275
rect 25780 18232 25832 18241
rect 26240 18275 26292 18284
rect 26240 18241 26249 18275
rect 26249 18241 26283 18275
rect 26283 18241 26292 18275
rect 26240 18232 26292 18241
rect 18696 18207 18748 18216
rect 18696 18173 18705 18207
rect 18705 18173 18739 18207
rect 18739 18173 18748 18207
rect 18696 18164 18748 18173
rect 19708 18164 19760 18216
rect 13544 18139 13596 18148
rect 13544 18105 13553 18139
rect 13553 18105 13587 18139
rect 13587 18105 13596 18139
rect 13544 18096 13596 18105
rect 16580 18096 16632 18148
rect 2872 18028 2924 18080
rect 6552 18028 6604 18080
rect 13084 18028 13136 18080
rect 14372 18028 14424 18080
rect 15292 18028 15344 18080
rect 16948 18028 17000 18080
rect 24860 18071 24912 18080
rect 24860 18037 24869 18071
rect 24869 18037 24903 18071
rect 24903 18037 24912 18071
rect 24860 18028 24912 18037
rect 4423 17926 4475 17978
rect 4487 17926 4539 17978
rect 4551 17926 4603 17978
rect 4615 17926 4667 17978
rect 4679 17926 4731 17978
rect 11369 17926 11421 17978
rect 11433 17926 11485 17978
rect 11497 17926 11549 17978
rect 11561 17926 11613 17978
rect 11625 17926 11677 17978
rect 18315 17926 18367 17978
rect 18379 17926 18431 17978
rect 18443 17926 18495 17978
rect 18507 17926 18559 17978
rect 18571 17926 18623 17978
rect 25261 17926 25313 17978
rect 25325 17926 25377 17978
rect 25389 17926 25441 17978
rect 25453 17926 25505 17978
rect 25517 17926 25569 17978
rect 2872 17867 2924 17876
rect 2872 17833 2881 17867
rect 2881 17833 2915 17867
rect 2915 17833 2924 17867
rect 2872 17824 2924 17833
rect 3976 17824 4028 17876
rect 11244 17824 11296 17876
rect 19708 17824 19760 17876
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 3240 17620 3292 17672
rect 8300 17688 8352 17740
rect 9404 17731 9456 17740
rect 9404 17697 9413 17731
rect 9413 17697 9447 17731
rect 9447 17697 9456 17731
rect 9404 17688 9456 17697
rect 10600 17688 10652 17740
rect 13176 17688 13228 17740
rect 23112 17688 23164 17740
rect 6736 17620 6788 17672
rect 7288 17620 7340 17672
rect 13820 17620 13872 17672
rect 19984 17663 20036 17672
rect 19984 17629 19993 17663
rect 19993 17629 20027 17663
rect 20027 17629 20036 17663
rect 19984 17620 20036 17629
rect 24676 17620 24728 17672
rect 24860 17663 24912 17672
rect 24860 17629 24894 17663
rect 24894 17629 24912 17663
rect 24860 17620 24912 17629
rect 27620 17620 27672 17672
rect 6368 17552 6420 17604
rect 6828 17484 6880 17536
rect 7380 17552 7432 17604
rect 12348 17552 12400 17604
rect 13728 17552 13780 17604
rect 14648 17595 14700 17604
rect 14648 17561 14657 17595
rect 14657 17561 14691 17595
rect 14691 17561 14700 17595
rect 14648 17552 14700 17561
rect 15200 17552 15252 17604
rect 16856 17552 16908 17604
rect 21640 17552 21692 17604
rect 28172 17595 28224 17604
rect 28172 17561 28181 17595
rect 28181 17561 28215 17595
rect 28215 17561 28224 17595
rect 28172 17552 28224 17561
rect 9956 17484 10008 17536
rect 12992 17484 13044 17536
rect 14372 17484 14424 17536
rect 17224 17484 17276 17536
rect 22284 17484 22336 17536
rect 24032 17484 24084 17536
rect 25136 17484 25188 17536
rect 25320 17484 25372 17536
rect 7896 17382 7948 17434
rect 7960 17382 8012 17434
rect 8024 17382 8076 17434
rect 8088 17382 8140 17434
rect 8152 17382 8204 17434
rect 14842 17382 14894 17434
rect 14906 17382 14958 17434
rect 14970 17382 15022 17434
rect 15034 17382 15086 17434
rect 15098 17382 15150 17434
rect 21788 17382 21840 17434
rect 21852 17382 21904 17434
rect 21916 17382 21968 17434
rect 21980 17382 22032 17434
rect 22044 17382 22096 17434
rect 28734 17382 28786 17434
rect 28798 17382 28850 17434
rect 28862 17382 28914 17434
rect 28926 17382 28978 17434
rect 28990 17382 29042 17434
rect 2964 17144 3016 17196
rect 4068 17144 4120 17196
rect 6736 17280 6788 17332
rect 14372 17280 14424 17332
rect 16856 17280 16908 17332
rect 5816 17144 5868 17196
rect 5908 17187 5960 17196
rect 5908 17153 5917 17187
rect 5917 17153 5951 17187
rect 5951 17153 5960 17187
rect 5908 17144 5960 17153
rect 7656 17144 7708 17196
rect 10600 17144 10652 17196
rect 11796 17144 11848 17196
rect 13084 17144 13136 17196
rect 13820 17187 13872 17196
rect 13820 17153 13829 17187
rect 13829 17153 13863 17187
rect 13863 17153 13872 17187
rect 13820 17144 13872 17153
rect 7380 17076 7432 17128
rect 13728 17076 13780 17128
rect 5540 17008 5592 17060
rect 12992 17008 13044 17060
rect 14648 17212 14700 17264
rect 15016 17187 15068 17196
rect 15016 17153 15025 17187
rect 15025 17153 15059 17187
rect 15059 17153 15068 17187
rect 15016 17144 15068 17153
rect 15200 17187 15252 17196
rect 15200 17153 15209 17187
rect 15209 17153 15243 17187
rect 15243 17153 15252 17187
rect 15200 17144 15252 17153
rect 17224 17212 17276 17264
rect 22284 17255 22336 17264
rect 22284 17221 22293 17255
rect 22293 17221 22327 17255
rect 22327 17221 22336 17255
rect 22284 17212 22336 17221
rect 22744 17212 22796 17264
rect 24032 17255 24084 17264
rect 24032 17221 24041 17255
rect 24041 17221 24075 17255
rect 24075 17221 24084 17255
rect 27896 17280 27948 17332
rect 24032 17212 24084 17221
rect 24492 17187 24544 17196
rect 24492 17153 24501 17187
rect 24501 17153 24535 17187
rect 24535 17153 24544 17187
rect 24492 17144 24544 17153
rect 25044 17212 25096 17264
rect 27252 17255 27304 17264
rect 27252 17221 27261 17255
rect 27261 17221 27295 17255
rect 27295 17221 27304 17255
rect 27252 17212 27304 17221
rect 24768 17144 24820 17196
rect 25320 17187 25372 17196
rect 25320 17153 25329 17187
rect 25329 17153 25363 17187
rect 25363 17153 25372 17187
rect 25320 17144 25372 17153
rect 26332 17187 26384 17196
rect 14740 17076 14792 17128
rect 15292 17076 15344 17128
rect 14280 17008 14332 17060
rect 15016 17008 15068 17060
rect 22284 17076 22336 17128
rect 22652 17076 22704 17128
rect 26332 17153 26341 17187
rect 26341 17153 26375 17187
rect 26375 17153 26384 17187
rect 26332 17144 26384 17153
rect 26884 17144 26936 17196
rect 2320 16940 2372 16992
rect 5724 16940 5776 16992
rect 9680 16940 9732 16992
rect 13084 16983 13136 16992
rect 13084 16949 13093 16983
rect 13093 16949 13127 16983
rect 13127 16949 13136 16983
rect 13084 16940 13136 16949
rect 14556 16940 14608 16992
rect 15200 16940 15252 16992
rect 15752 16940 15804 16992
rect 18236 16940 18288 16992
rect 4423 16838 4475 16890
rect 4487 16838 4539 16890
rect 4551 16838 4603 16890
rect 4615 16838 4667 16890
rect 4679 16838 4731 16890
rect 11369 16838 11421 16890
rect 11433 16838 11485 16890
rect 11497 16838 11549 16890
rect 11561 16838 11613 16890
rect 11625 16838 11677 16890
rect 18315 16838 18367 16890
rect 18379 16838 18431 16890
rect 18443 16838 18495 16890
rect 18507 16838 18559 16890
rect 18571 16838 18623 16890
rect 25261 16838 25313 16890
rect 25325 16838 25377 16890
rect 25389 16838 25441 16890
rect 25453 16838 25505 16890
rect 25517 16838 25569 16890
rect 8300 16779 8352 16788
rect 8300 16745 8309 16779
rect 8309 16745 8343 16779
rect 8343 16745 8352 16779
rect 8300 16736 8352 16745
rect 6552 16643 6604 16652
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 6552 16600 6604 16609
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 10600 16736 10652 16788
rect 12348 16779 12400 16788
rect 12348 16745 12357 16779
rect 12357 16745 12391 16779
rect 12391 16745 12400 16779
rect 12348 16736 12400 16745
rect 23112 16736 23164 16788
rect 26332 16736 26384 16788
rect 27620 16779 27672 16788
rect 27620 16745 27629 16779
rect 27629 16745 27663 16779
rect 27663 16745 27672 16779
rect 27620 16736 27672 16745
rect 11704 16643 11756 16652
rect 11704 16609 11713 16643
rect 11713 16609 11747 16643
rect 11747 16609 11756 16643
rect 11704 16600 11756 16609
rect 2596 16532 2648 16584
rect 3240 16532 3292 16584
rect 2044 16396 2096 16448
rect 3332 16396 3384 16448
rect 5540 16396 5592 16448
rect 7012 16396 7064 16448
rect 12256 16532 12308 16584
rect 13084 16600 13136 16652
rect 14188 16600 14240 16652
rect 16580 16668 16632 16720
rect 24032 16711 24084 16720
rect 24032 16677 24041 16711
rect 24041 16677 24075 16711
rect 24075 16677 24084 16711
rect 24032 16668 24084 16677
rect 24768 16668 24820 16720
rect 14648 16643 14700 16652
rect 12992 16575 13044 16584
rect 12992 16541 13001 16575
rect 13001 16541 13035 16575
rect 13035 16541 13044 16575
rect 12992 16532 13044 16541
rect 13176 16575 13228 16584
rect 13176 16541 13185 16575
rect 13185 16541 13219 16575
rect 13219 16541 13228 16575
rect 13176 16532 13228 16541
rect 9220 16464 9272 16516
rect 12900 16464 12952 16516
rect 13728 16532 13780 16584
rect 14648 16609 14657 16643
rect 14657 16609 14691 16643
rect 14691 16609 14700 16643
rect 14648 16600 14700 16609
rect 14740 16575 14792 16584
rect 14740 16541 14749 16575
rect 14749 16541 14783 16575
rect 14783 16541 14792 16575
rect 14740 16532 14792 16541
rect 15200 16532 15252 16584
rect 18236 16643 18288 16652
rect 18236 16609 18245 16643
rect 18245 16609 18279 16643
rect 18279 16609 18288 16643
rect 18236 16600 18288 16609
rect 20628 16600 20680 16652
rect 22284 16643 22336 16652
rect 22284 16609 22293 16643
rect 22293 16609 22327 16643
rect 22327 16609 22336 16643
rect 22284 16600 22336 16609
rect 26884 16600 26936 16652
rect 24492 16532 24544 16584
rect 25044 16575 25096 16584
rect 25044 16541 25053 16575
rect 25053 16541 25087 16575
rect 25087 16541 25096 16575
rect 25044 16532 25096 16541
rect 27252 16575 27304 16584
rect 27252 16541 27261 16575
rect 27261 16541 27295 16575
rect 27295 16541 27304 16575
rect 27252 16532 27304 16541
rect 13820 16464 13872 16516
rect 14096 16464 14148 16516
rect 22468 16464 22520 16516
rect 9496 16396 9548 16448
rect 12072 16396 12124 16448
rect 18880 16439 18932 16448
rect 18880 16405 18889 16439
rect 18889 16405 18923 16439
rect 18923 16405 18932 16439
rect 18880 16396 18932 16405
rect 22836 16464 22888 16516
rect 25136 16464 25188 16516
rect 22928 16396 22980 16448
rect 7896 16294 7948 16346
rect 7960 16294 8012 16346
rect 8024 16294 8076 16346
rect 8088 16294 8140 16346
rect 8152 16294 8204 16346
rect 14842 16294 14894 16346
rect 14906 16294 14958 16346
rect 14970 16294 15022 16346
rect 15034 16294 15086 16346
rect 15098 16294 15150 16346
rect 21788 16294 21840 16346
rect 21852 16294 21904 16346
rect 21916 16294 21968 16346
rect 21980 16294 22032 16346
rect 22044 16294 22096 16346
rect 28734 16294 28786 16346
rect 28798 16294 28850 16346
rect 28862 16294 28914 16346
rect 28926 16294 28978 16346
rect 28990 16294 29042 16346
rect 9220 16192 9272 16244
rect 9404 16192 9456 16244
rect 11796 16192 11848 16244
rect 13084 16192 13136 16244
rect 13452 16235 13504 16244
rect 13452 16201 13461 16235
rect 13461 16201 13495 16235
rect 13495 16201 13504 16235
rect 13452 16192 13504 16201
rect 2320 16167 2372 16176
rect 2320 16133 2329 16167
rect 2329 16133 2363 16167
rect 2363 16133 2372 16167
rect 2320 16124 2372 16133
rect 3332 16124 3384 16176
rect 4068 16167 4120 16176
rect 4068 16133 4077 16167
rect 4077 16133 4111 16167
rect 4111 16133 4120 16167
rect 4068 16124 4120 16133
rect 9312 16124 9364 16176
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 5816 16056 5868 16108
rect 11980 16056 12032 16108
rect 12256 16124 12308 16176
rect 15936 16167 15988 16176
rect 15936 16133 15945 16167
rect 15945 16133 15979 16167
rect 15979 16133 15988 16167
rect 15936 16124 15988 16133
rect 16488 16124 16540 16176
rect 12624 16056 12676 16108
rect 13176 16056 13228 16108
rect 13728 16056 13780 16108
rect 14740 16099 14792 16108
rect 14740 16065 14749 16099
rect 14749 16065 14783 16099
rect 14783 16065 14792 16099
rect 14740 16056 14792 16065
rect 17776 16099 17828 16108
rect 17776 16065 17810 16099
rect 17810 16065 17828 16099
rect 17776 16056 17828 16065
rect 6552 16031 6604 16040
rect 6552 15997 6561 16031
rect 6561 15997 6595 16031
rect 6595 15997 6604 16031
rect 6552 15988 6604 15997
rect 7380 16031 7432 16040
rect 7380 15997 7389 16031
rect 7389 15997 7423 16031
rect 7423 15997 7432 16031
rect 7380 15988 7432 15997
rect 9588 15988 9640 16040
rect 11060 15988 11112 16040
rect 11704 15988 11756 16040
rect 15752 16031 15804 16040
rect 15752 15997 15761 16031
rect 15761 15997 15795 16031
rect 15795 15997 15804 16031
rect 15752 15988 15804 15997
rect 17408 15988 17460 16040
rect 17500 16031 17552 16040
rect 17500 15997 17509 16031
rect 17509 15997 17543 16031
rect 17543 15997 17552 16031
rect 17500 15988 17552 15997
rect 12440 15920 12492 15972
rect 12900 15920 12952 15972
rect 10968 15852 11020 15904
rect 11980 15852 12032 15904
rect 14464 15852 14516 15904
rect 16672 15920 16724 15972
rect 18880 16124 18932 16176
rect 22744 16192 22796 16244
rect 22928 16192 22980 16244
rect 24032 16192 24084 16244
rect 22468 16124 22520 16176
rect 22376 16099 22428 16108
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 22284 15988 22336 16040
rect 22928 16056 22980 16108
rect 23020 16056 23072 16108
rect 23112 15988 23164 16040
rect 23848 15988 23900 16040
rect 16580 15852 16632 15904
rect 18880 15895 18932 15904
rect 18880 15861 18889 15895
rect 18889 15861 18923 15895
rect 18923 15861 18932 15895
rect 18880 15852 18932 15861
rect 20628 15920 20680 15972
rect 21640 15852 21692 15904
rect 4423 15750 4475 15802
rect 4487 15750 4539 15802
rect 4551 15750 4603 15802
rect 4615 15750 4667 15802
rect 4679 15750 4731 15802
rect 11369 15750 11421 15802
rect 11433 15750 11485 15802
rect 11497 15750 11549 15802
rect 11561 15750 11613 15802
rect 11625 15750 11677 15802
rect 18315 15750 18367 15802
rect 18379 15750 18431 15802
rect 18443 15750 18495 15802
rect 18507 15750 18559 15802
rect 18571 15750 18623 15802
rect 25261 15750 25313 15802
rect 25325 15750 25377 15802
rect 25389 15750 25441 15802
rect 25453 15750 25505 15802
rect 25517 15750 25569 15802
rect 7288 15691 7340 15700
rect 7288 15657 7297 15691
rect 7297 15657 7331 15691
rect 7331 15657 7340 15691
rect 7288 15648 7340 15657
rect 17408 15648 17460 15700
rect 22836 15691 22888 15700
rect 22836 15657 22845 15691
rect 22845 15657 22879 15691
rect 22879 15657 22888 15691
rect 22836 15648 22888 15657
rect 11060 15580 11112 15632
rect 14096 15580 14148 15632
rect 4344 15512 4396 15564
rect 2596 15487 2648 15496
rect 2596 15453 2605 15487
rect 2605 15453 2639 15487
rect 2639 15453 2648 15487
rect 2596 15444 2648 15453
rect 3240 15444 3292 15496
rect 5540 15487 5592 15496
rect 5540 15453 5549 15487
rect 5549 15453 5583 15487
rect 5583 15453 5592 15487
rect 5540 15444 5592 15453
rect 9680 15487 9732 15496
rect 9680 15453 9689 15487
rect 9689 15453 9723 15487
rect 9723 15453 9732 15487
rect 9680 15444 9732 15453
rect 10968 15512 11020 15564
rect 12440 15555 12492 15564
rect 12440 15521 12449 15555
rect 12449 15521 12483 15555
rect 12483 15521 12492 15555
rect 12440 15512 12492 15521
rect 20536 15512 20588 15564
rect 20904 15512 20956 15564
rect 2780 15376 2832 15428
rect 5724 15376 5776 15428
rect 6552 15376 6604 15428
rect 9956 15419 10008 15428
rect 9956 15385 9965 15419
rect 9965 15385 9999 15419
rect 9999 15385 10008 15419
rect 9956 15376 10008 15385
rect 12624 15419 12676 15428
rect 12624 15385 12633 15419
rect 12633 15385 12667 15419
rect 12667 15385 12676 15419
rect 12624 15376 12676 15385
rect 12808 15419 12860 15428
rect 12808 15385 12817 15419
rect 12817 15385 12851 15419
rect 12851 15385 12860 15419
rect 12808 15376 12860 15385
rect 12992 15376 13044 15428
rect 13268 15376 13320 15428
rect 16580 15444 16632 15496
rect 20720 15444 20772 15496
rect 22376 15444 22428 15496
rect 22928 15487 22980 15496
rect 22928 15453 22937 15487
rect 22937 15453 22971 15487
rect 22971 15453 22980 15487
rect 22928 15444 22980 15453
rect 26148 15487 26200 15496
rect 26148 15453 26157 15487
rect 26157 15453 26191 15487
rect 26191 15453 26200 15487
rect 26148 15444 26200 15453
rect 17500 15376 17552 15428
rect 1860 15351 1912 15360
rect 1860 15317 1869 15351
rect 1869 15317 1903 15351
rect 1903 15317 1912 15351
rect 1860 15308 1912 15317
rect 2504 15351 2556 15360
rect 2504 15317 2513 15351
rect 2513 15317 2547 15351
rect 2547 15317 2556 15351
rect 2504 15308 2556 15317
rect 3240 15351 3292 15360
rect 3240 15317 3249 15351
rect 3249 15317 3283 15351
rect 3283 15317 3292 15351
rect 3240 15308 3292 15317
rect 10508 15308 10560 15360
rect 11060 15308 11112 15360
rect 11244 15351 11296 15360
rect 11244 15317 11253 15351
rect 11253 15317 11287 15351
rect 11287 15317 11296 15351
rect 11244 15308 11296 15317
rect 13452 15308 13504 15360
rect 14740 15308 14792 15360
rect 25964 15308 26016 15360
rect 7896 15206 7948 15258
rect 7960 15206 8012 15258
rect 8024 15206 8076 15258
rect 8088 15206 8140 15258
rect 8152 15206 8204 15258
rect 14842 15206 14894 15258
rect 14906 15206 14958 15258
rect 14970 15206 15022 15258
rect 15034 15206 15086 15258
rect 15098 15206 15150 15258
rect 21788 15206 21840 15258
rect 21852 15206 21904 15258
rect 21916 15206 21968 15258
rect 21980 15206 22032 15258
rect 22044 15206 22096 15258
rect 28734 15206 28786 15258
rect 28798 15206 28850 15258
rect 28862 15206 28914 15258
rect 28926 15206 28978 15258
rect 28990 15206 29042 15258
rect 17776 15104 17828 15156
rect 17960 15104 18012 15156
rect 24952 15147 25004 15156
rect 24952 15113 24961 15147
rect 24961 15113 24995 15147
rect 24995 15113 25004 15147
rect 24952 15104 25004 15113
rect 2504 15036 2556 15088
rect 3240 15036 3292 15088
rect 1860 14968 1912 15020
rect 5080 15011 5132 15020
rect 5080 14977 5089 15011
rect 5089 14977 5123 15011
rect 5123 14977 5132 15011
rect 5080 14968 5132 14977
rect 6552 15011 6604 15020
rect 6552 14977 6561 15011
rect 6561 14977 6595 15011
rect 6595 14977 6604 15011
rect 6552 14968 6604 14977
rect 7472 15011 7524 15020
rect 7472 14977 7481 15011
rect 7481 14977 7515 15011
rect 7515 14977 7524 15011
rect 7472 14968 7524 14977
rect 10416 14968 10468 15020
rect 11244 14968 11296 15020
rect 12348 14968 12400 15020
rect 13452 15011 13504 15020
rect 13452 14977 13461 15011
rect 13461 14977 13495 15011
rect 13495 14977 13504 15011
rect 13452 14968 13504 14977
rect 13728 14968 13780 15020
rect 2596 14900 2648 14952
rect 6644 14807 6696 14816
rect 6644 14773 6653 14807
rect 6653 14773 6687 14807
rect 6687 14773 6696 14807
rect 6644 14764 6696 14773
rect 7564 14807 7616 14816
rect 7564 14773 7573 14807
rect 7573 14773 7607 14807
rect 7607 14773 7616 14807
rect 7564 14764 7616 14773
rect 12900 14900 12952 14952
rect 15568 15011 15620 15020
rect 15568 14977 15577 15011
rect 15577 14977 15611 15011
rect 15611 14977 15620 15011
rect 15568 14968 15620 14977
rect 24768 15036 24820 15088
rect 25044 15036 25096 15088
rect 20720 15011 20772 15020
rect 20720 14977 20729 15011
rect 20729 14977 20763 15011
rect 20763 14977 20772 15011
rect 21364 15011 21416 15020
rect 20720 14968 20772 14977
rect 21364 14977 21373 15011
rect 21373 14977 21407 15011
rect 21407 14977 21416 15011
rect 21364 14968 21416 14977
rect 26792 14968 26844 15020
rect 27988 14968 28040 15020
rect 14280 14875 14332 14884
rect 14280 14841 14289 14875
rect 14289 14841 14323 14875
rect 14323 14841 14332 14875
rect 14280 14832 14332 14841
rect 14832 14832 14884 14884
rect 9956 14764 10008 14816
rect 10876 14764 10928 14816
rect 13452 14764 13504 14816
rect 13728 14764 13780 14816
rect 15292 14900 15344 14952
rect 16028 14900 16080 14952
rect 18236 14900 18288 14952
rect 18880 14900 18932 14952
rect 19616 14807 19668 14816
rect 19616 14773 19625 14807
rect 19625 14773 19659 14807
rect 19659 14773 19668 14807
rect 19616 14764 19668 14773
rect 20352 14764 20404 14816
rect 21272 14807 21324 14816
rect 21272 14773 21281 14807
rect 21281 14773 21315 14807
rect 21315 14773 21324 14807
rect 21272 14764 21324 14773
rect 26516 14943 26568 14952
rect 26148 14832 26200 14884
rect 26516 14909 26525 14943
rect 26525 14909 26559 14943
rect 26559 14909 26568 14943
rect 26516 14900 26568 14909
rect 27436 14832 27488 14884
rect 27252 14807 27304 14816
rect 27252 14773 27261 14807
rect 27261 14773 27295 14807
rect 27295 14773 27304 14807
rect 27252 14764 27304 14773
rect 4423 14662 4475 14714
rect 4487 14662 4539 14714
rect 4551 14662 4603 14714
rect 4615 14662 4667 14714
rect 4679 14662 4731 14714
rect 11369 14662 11421 14714
rect 11433 14662 11485 14714
rect 11497 14662 11549 14714
rect 11561 14662 11613 14714
rect 11625 14662 11677 14714
rect 18315 14662 18367 14714
rect 18379 14662 18431 14714
rect 18443 14662 18495 14714
rect 18507 14662 18559 14714
rect 18571 14662 18623 14714
rect 25261 14662 25313 14714
rect 25325 14662 25377 14714
rect 25389 14662 25441 14714
rect 25453 14662 25505 14714
rect 25517 14662 25569 14714
rect 5540 14492 5592 14544
rect 2780 14399 2832 14408
rect 2780 14365 2789 14399
rect 2789 14365 2823 14399
rect 2823 14365 2832 14399
rect 2780 14356 2832 14365
rect 3056 14356 3108 14408
rect 6552 14424 6604 14476
rect 5540 14356 5592 14408
rect 9588 14560 9640 14612
rect 11244 14560 11296 14612
rect 12808 14560 12860 14612
rect 13452 14560 13504 14612
rect 15568 14560 15620 14612
rect 26148 14560 26200 14612
rect 18696 14492 18748 14544
rect 10508 14467 10560 14476
rect 10508 14433 10517 14467
rect 10517 14433 10551 14467
rect 10551 14433 10560 14467
rect 10508 14424 10560 14433
rect 12900 14424 12952 14476
rect 14188 14424 14240 14476
rect 20352 14467 20404 14476
rect 9588 14356 9640 14408
rect 9956 14356 10008 14408
rect 12348 14399 12400 14408
rect 12348 14365 12357 14399
rect 12357 14365 12391 14399
rect 12391 14365 12400 14399
rect 12348 14356 12400 14365
rect 5908 14331 5960 14340
rect 5908 14297 5917 14331
rect 5917 14297 5951 14331
rect 5951 14297 5960 14331
rect 5908 14288 5960 14297
rect 6644 14288 6696 14340
rect 7472 14288 7524 14340
rect 12624 14288 12676 14340
rect 14556 14356 14608 14408
rect 14832 14399 14884 14408
rect 14832 14365 14841 14399
rect 14841 14365 14875 14399
rect 14875 14365 14884 14399
rect 20352 14433 20361 14467
rect 20361 14433 20395 14467
rect 20395 14433 20404 14467
rect 20352 14424 20404 14433
rect 21272 14424 21324 14476
rect 21364 14424 21416 14476
rect 24952 14424 25004 14476
rect 25964 14467 26016 14476
rect 25964 14433 25973 14467
rect 25973 14433 26007 14467
rect 26007 14433 26016 14467
rect 25964 14424 26016 14433
rect 14832 14356 14884 14365
rect 13820 14288 13872 14340
rect 14372 14288 14424 14340
rect 17500 14288 17552 14340
rect 21180 14288 21232 14340
rect 26516 14288 26568 14340
rect 1584 14220 1636 14272
rect 2320 14220 2372 14272
rect 3332 14263 3384 14272
rect 3332 14229 3341 14263
rect 3341 14229 3375 14263
rect 3375 14229 3384 14263
rect 3332 14220 3384 14229
rect 5080 14263 5132 14272
rect 5080 14229 5089 14263
rect 5089 14229 5123 14263
rect 5123 14229 5132 14263
rect 5080 14220 5132 14229
rect 8208 14263 8260 14272
rect 8208 14229 8217 14263
rect 8217 14229 8251 14263
rect 8251 14229 8260 14263
rect 8208 14220 8260 14229
rect 13452 14220 13504 14272
rect 15660 14220 15712 14272
rect 17224 14220 17276 14272
rect 20720 14220 20772 14272
rect 7896 14118 7948 14170
rect 7960 14118 8012 14170
rect 8024 14118 8076 14170
rect 8088 14118 8140 14170
rect 8152 14118 8204 14170
rect 14842 14118 14894 14170
rect 14906 14118 14958 14170
rect 14970 14118 15022 14170
rect 15034 14118 15086 14170
rect 15098 14118 15150 14170
rect 21788 14118 21840 14170
rect 21852 14118 21904 14170
rect 21916 14118 21968 14170
rect 21980 14118 22032 14170
rect 22044 14118 22096 14170
rect 28734 14118 28786 14170
rect 28798 14118 28850 14170
rect 28862 14118 28914 14170
rect 28926 14118 28978 14170
rect 28990 14118 29042 14170
rect 5540 14059 5592 14068
rect 5540 14025 5549 14059
rect 5549 14025 5583 14059
rect 5583 14025 5592 14059
rect 5540 14016 5592 14025
rect 5908 14016 5960 14068
rect 9588 14016 9640 14068
rect 10416 14059 10468 14068
rect 10416 14025 10425 14059
rect 10425 14025 10459 14059
rect 10459 14025 10468 14059
rect 10416 14016 10468 14025
rect 10876 14059 10928 14068
rect 10876 14025 10885 14059
rect 10885 14025 10919 14059
rect 10919 14025 10928 14059
rect 10876 14016 10928 14025
rect 2320 13991 2372 14000
rect 2320 13957 2329 13991
rect 2329 13957 2363 13991
rect 2363 13957 2372 13991
rect 2320 13948 2372 13957
rect 3332 13948 3384 14000
rect 8208 13991 8260 14000
rect 8208 13957 8217 13991
rect 8217 13957 8251 13991
rect 8251 13957 8260 13991
rect 8208 13948 8260 13957
rect 9864 13948 9916 14000
rect 4804 13923 4856 13932
rect 4804 13889 4813 13923
rect 4813 13889 4847 13923
rect 4847 13889 4856 13923
rect 4804 13880 4856 13889
rect 7472 13880 7524 13932
rect 7564 13880 7616 13932
rect 10784 13923 10836 13932
rect 10784 13889 10793 13923
rect 10793 13889 10827 13923
rect 10827 13889 10836 13923
rect 10784 13880 10836 13889
rect 12164 13923 12216 13932
rect 12164 13889 12173 13923
rect 12173 13889 12207 13923
rect 12207 13889 12216 13923
rect 12164 13880 12216 13889
rect 14280 14016 14332 14068
rect 15384 14016 15436 14068
rect 13452 13948 13504 14000
rect 17224 13948 17276 14000
rect 24768 14016 24820 14068
rect 14188 13880 14240 13932
rect 15476 13923 15528 13932
rect 2044 13855 2096 13864
rect 2044 13821 2053 13855
rect 2053 13821 2087 13855
rect 2087 13821 2096 13855
rect 2044 13812 2096 13821
rect 2780 13812 2832 13864
rect 5816 13812 5868 13864
rect 10968 13855 11020 13864
rect 10968 13821 10977 13855
rect 10977 13821 11011 13855
rect 11011 13821 11020 13855
rect 10968 13812 11020 13821
rect 12624 13812 12676 13864
rect 13360 13676 13412 13728
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 15660 13923 15712 13932
rect 15660 13889 15669 13923
rect 15669 13889 15703 13923
rect 15703 13889 15712 13923
rect 15660 13880 15712 13889
rect 17408 13880 17460 13932
rect 17776 13880 17828 13932
rect 21180 13991 21232 14000
rect 21180 13957 21189 13991
rect 21189 13957 21223 13991
rect 21223 13957 21232 13991
rect 21180 13948 21232 13957
rect 27804 13948 27856 14000
rect 21456 13880 21508 13932
rect 21548 13880 21600 13932
rect 23112 13923 23164 13932
rect 23112 13889 23146 13923
rect 23146 13889 23164 13923
rect 26424 13923 26476 13932
rect 23112 13880 23164 13889
rect 26424 13889 26433 13923
rect 26433 13889 26467 13923
rect 26467 13889 26476 13923
rect 26424 13880 26476 13889
rect 26792 13880 26844 13932
rect 27344 13880 27396 13932
rect 17592 13812 17644 13864
rect 17960 13812 18012 13864
rect 19432 13812 19484 13864
rect 20628 13855 20680 13864
rect 20628 13821 20637 13855
rect 20637 13821 20671 13855
rect 20671 13821 20680 13855
rect 20628 13812 20680 13821
rect 20812 13812 20864 13864
rect 21088 13744 21140 13796
rect 27436 13855 27488 13864
rect 27436 13821 27445 13855
rect 27445 13821 27479 13855
rect 27479 13821 27488 13855
rect 27436 13812 27488 13821
rect 18236 13719 18288 13728
rect 18236 13685 18245 13719
rect 18245 13685 18279 13719
rect 18279 13685 18288 13719
rect 18236 13676 18288 13685
rect 23572 13676 23624 13728
rect 26240 13676 26292 13728
rect 4423 13574 4475 13626
rect 4487 13574 4539 13626
rect 4551 13574 4603 13626
rect 4615 13574 4667 13626
rect 4679 13574 4731 13626
rect 11369 13574 11421 13626
rect 11433 13574 11485 13626
rect 11497 13574 11549 13626
rect 11561 13574 11613 13626
rect 11625 13574 11677 13626
rect 18315 13574 18367 13626
rect 18379 13574 18431 13626
rect 18443 13574 18495 13626
rect 18507 13574 18559 13626
rect 18571 13574 18623 13626
rect 25261 13574 25313 13626
rect 25325 13574 25377 13626
rect 25389 13574 25441 13626
rect 25453 13574 25505 13626
rect 25517 13574 25569 13626
rect 2044 13472 2096 13524
rect 4804 13336 4856 13388
rect 5816 13379 5868 13388
rect 5816 13345 5825 13379
rect 5825 13345 5859 13379
rect 5859 13345 5868 13379
rect 5816 13336 5868 13345
rect 23112 13515 23164 13524
rect 23112 13481 23121 13515
rect 23121 13481 23155 13515
rect 23155 13481 23164 13515
rect 23112 13472 23164 13481
rect 27988 13515 28040 13524
rect 27988 13481 27997 13515
rect 27997 13481 28031 13515
rect 28031 13481 28040 13515
rect 27988 13472 28040 13481
rect 9864 13447 9916 13456
rect 9864 13413 9873 13447
rect 9873 13413 9907 13447
rect 9907 13413 9916 13447
rect 9864 13404 9916 13413
rect 14648 13404 14700 13456
rect 3056 13311 3108 13320
rect 3056 13277 3065 13311
rect 3065 13277 3099 13311
rect 3099 13277 3108 13311
rect 3056 13268 3108 13277
rect 6552 13311 6604 13320
rect 6552 13277 6561 13311
rect 6561 13277 6595 13311
rect 6595 13277 6604 13311
rect 6552 13268 6604 13277
rect 9956 13268 10008 13320
rect 10968 13311 11020 13320
rect 10968 13277 10977 13311
rect 10977 13277 11011 13311
rect 11011 13277 11020 13311
rect 10968 13268 11020 13277
rect 11704 13311 11756 13320
rect 11704 13277 11713 13311
rect 11713 13277 11747 13311
rect 11747 13277 11756 13311
rect 11704 13268 11756 13277
rect 3608 13200 3660 13252
rect 5080 13200 5132 13252
rect 6644 13200 6696 13252
rect 7196 13200 7248 13252
rect 9312 13200 9364 13252
rect 23572 13379 23624 13388
rect 12164 13311 12216 13320
rect 12164 13277 12173 13311
rect 12173 13277 12207 13311
rect 12207 13277 12216 13311
rect 12164 13268 12216 13277
rect 12992 13311 13044 13320
rect 12992 13277 13001 13311
rect 13001 13277 13035 13311
rect 13035 13277 13044 13311
rect 12992 13268 13044 13277
rect 14372 13268 14424 13320
rect 15292 13268 15344 13320
rect 15476 13268 15528 13320
rect 16488 13268 16540 13320
rect 17592 13311 17644 13320
rect 17592 13277 17601 13311
rect 17601 13277 17635 13311
rect 17635 13277 17644 13311
rect 17592 13268 17644 13277
rect 17684 13311 17736 13320
rect 17684 13277 17694 13311
rect 17694 13277 17728 13311
rect 17728 13277 17736 13311
rect 17960 13311 18012 13320
rect 17684 13268 17736 13277
rect 17960 13277 17969 13311
rect 17969 13277 18003 13311
rect 18003 13277 18012 13311
rect 17960 13268 18012 13277
rect 18236 13268 18288 13320
rect 19524 13311 19576 13320
rect 19524 13277 19533 13311
rect 19533 13277 19567 13311
rect 19567 13277 19576 13311
rect 19524 13268 19576 13277
rect 12808 13200 12860 13252
rect 16856 13200 16908 13252
rect 17040 13200 17092 13252
rect 23572 13345 23581 13379
rect 23581 13345 23615 13379
rect 23615 13345 23624 13379
rect 23572 13336 23624 13345
rect 23756 13379 23808 13388
rect 23756 13345 23765 13379
rect 23765 13345 23799 13379
rect 23799 13345 23808 13379
rect 23756 13336 23808 13345
rect 24584 13379 24636 13388
rect 24584 13345 24593 13379
rect 24593 13345 24627 13379
rect 24627 13345 24636 13379
rect 24584 13336 24636 13345
rect 26240 13379 26292 13388
rect 26240 13345 26249 13379
rect 26249 13345 26283 13379
rect 26283 13345 26292 13379
rect 26240 13336 26292 13345
rect 27252 13336 27304 13388
rect 20996 13268 21048 13320
rect 23480 13311 23532 13320
rect 23480 13277 23489 13311
rect 23489 13277 23523 13311
rect 23523 13277 23532 13311
rect 23480 13268 23532 13277
rect 1860 13132 1912 13184
rect 2964 13175 3016 13184
rect 2964 13141 2973 13175
rect 2973 13141 3007 13175
rect 3007 13141 3016 13175
rect 2964 13132 3016 13141
rect 7012 13132 7064 13184
rect 11152 13132 11204 13184
rect 14648 13132 14700 13184
rect 16948 13132 17000 13184
rect 26424 13200 26476 13252
rect 27804 13200 27856 13252
rect 19432 13132 19484 13184
rect 19984 13132 20036 13184
rect 22376 13175 22428 13184
rect 22376 13141 22385 13175
rect 22385 13141 22419 13175
rect 22419 13141 22428 13175
rect 22376 13132 22428 13141
rect 7896 13030 7948 13082
rect 7960 13030 8012 13082
rect 8024 13030 8076 13082
rect 8088 13030 8140 13082
rect 8152 13030 8204 13082
rect 14842 13030 14894 13082
rect 14906 13030 14958 13082
rect 14970 13030 15022 13082
rect 15034 13030 15086 13082
rect 15098 13030 15150 13082
rect 21788 13030 21840 13082
rect 21852 13030 21904 13082
rect 21916 13030 21968 13082
rect 21980 13030 22032 13082
rect 22044 13030 22096 13082
rect 28734 13030 28786 13082
rect 28798 13030 28850 13082
rect 28862 13030 28914 13082
rect 28926 13030 28978 13082
rect 28990 13030 29042 13082
rect 6644 12928 6696 12980
rect 7012 12971 7064 12980
rect 7012 12937 7021 12971
rect 7021 12937 7055 12971
rect 7055 12937 7064 12971
rect 7012 12928 7064 12937
rect 13452 12971 13504 12980
rect 1860 12903 1912 12912
rect 1860 12869 1869 12903
rect 1869 12869 1903 12903
rect 1903 12869 1912 12903
rect 1860 12860 1912 12869
rect 3608 12903 3660 12912
rect 3608 12869 3617 12903
rect 3617 12869 3651 12903
rect 3651 12869 3660 12903
rect 3608 12860 3660 12869
rect 6092 12860 6144 12912
rect 1584 12835 1636 12844
rect 1584 12801 1593 12835
rect 1593 12801 1627 12835
rect 1627 12801 1636 12835
rect 1584 12792 1636 12801
rect 2964 12792 3016 12844
rect 4804 12792 4856 12844
rect 5724 12792 5776 12844
rect 6552 12792 6604 12844
rect 10784 12860 10836 12912
rect 9772 12792 9824 12844
rect 13452 12937 13461 12971
rect 13461 12937 13495 12971
rect 13495 12937 13504 12971
rect 13452 12928 13504 12937
rect 16856 12971 16908 12980
rect 16856 12937 16865 12971
rect 16865 12937 16899 12971
rect 16899 12937 16908 12971
rect 16856 12928 16908 12937
rect 16948 12928 17000 12980
rect 20996 12971 21048 12980
rect 20996 12937 21005 12971
rect 21005 12937 21039 12971
rect 21039 12937 21048 12971
rect 20996 12928 21048 12937
rect 14740 12903 14792 12912
rect 14740 12869 14749 12903
rect 14749 12869 14783 12903
rect 14783 12869 14792 12903
rect 14740 12860 14792 12869
rect 15384 12903 15436 12912
rect 15384 12869 15393 12903
rect 15393 12869 15427 12903
rect 15427 12869 15436 12903
rect 15384 12860 15436 12869
rect 17684 12860 17736 12912
rect 7196 12767 7248 12776
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 13360 12724 13412 12776
rect 9956 12656 10008 12708
rect 10876 12656 10928 12708
rect 15660 12792 15712 12844
rect 16672 12792 16724 12844
rect 17224 12835 17276 12844
rect 17224 12801 17233 12835
rect 17233 12801 17267 12835
rect 17267 12801 17276 12835
rect 17224 12792 17276 12801
rect 21088 12860 21140 12912
rect 19432 12792 19484 12844
rect 24584 12928 24636 12980
rect 22468 12860 22520 12912
rect 28172 12903 28224 12912
rect 28172 12869 28181 12903
rect 28181 12869 28215 12903
rect 28215 12869 28224 12903
rect 28172 12860 28224 12869
rect 22376 12792 22428 12844
rect 22560 12835 22612 12844
rect 22560 12801 22594 12835
rect 22594 12801 22612 12835
rect 26332 12835 26384 12844
rect 22560 12792 22612 12801
rect 26332 12801 26341 12835
rect 26341 12801 26375 12835
rect 26375 12801 26384 12835
rect 26332 12792 26384 12801
rect 26424 12792 26476 12844
rect 27436 12792 27488 12844
rect 27620 12792 27672 12844
rect 17500 12767 17552 12776
rect 17500 12733 17509 12767
rect 17509 12733 17543 12767
rect 17543 12733 17552 12767
rect 17500 12724 17552 12733
rect 21272 12767 21324 12776
rect 21272 12733 21281 12767
rect 21281 12733 21315 12767
rect 21315 12733 21324 12767
rect 21272 12724 21324 12733
rect 5448 12588 5500 12640
rect 8484 12631 8536 12640
rect 8484 12597 8493 12631
rect 8493 12597 8527 12631
rect 8527 12597 8536 12631
rect 8484 12588 8536 12597
rect 10692 12588 10744 12640
rect 19800 12588 19852 12640
rect 19892 12588 19944 12640
rect 20904 12588 20956 12640
rect 23664 12631 23716 12640
rect 23664 12597 23673 12631
rect 23673 12597 23707 12631
rect 23707 12597 23716 12631
rect 23664 12588 23716 12597
rect 26424 12631 26476 12640
rect 26424 12597 26433 12631
rect 26433 12597 26467 12631
rect 26467 12597 26476 12631
rect 26424 12588 26476 12597
rect 26700 12588 26752 12640
rect 4423 12486 4475 12538
rect 4487 12486 4539 12538
rect 4551 12486 4603 12538
rect 4615 12486 4667 12538
rect 4679 12486 4731 12538
rect 11369 12486 11421 12538
rect 11433 12486 11485 12538
rect 11497 12486 11549 12538
rect 11561 12486 11613 12538
rect 11625 12486 11677 12538
rect 18315 12486 18367 12538
rect 18379 12486 18431 12538
rect 18443 12486 18495 12538
rect 18507 12486 18559 12538
rect 18571 12486 18623 12538
rect 25261 12486 25313 12538
rect 25325 12486 25377 12538
rect 25389 12486 25441 12538
rect 25453 12486 25505 12538
rect 25517 12486 25569 12538
rect 9772 12384 9824 12436
rect 14188 12384 14240 12436
rect 17040 12384 17092 12436
rect 17592 12384 17644 12436
rect 19432 12427 19484 12436
rect 19432 12393 19441 12427
rect 19441 12393 19475 12427
rect 19475 12393 19484 12427
rect 19432 12384 19484 12393
rect 21272 12384 21324 12436
rect 22560 12384 22612 12436
rect 27436 12384 27488 12436
rect 10784 12316 10836 12368
rect 5724 12291 5776 12300
rect 5724 12257 5733 12291
rect 5733 12257 5767 12291
rect 5767 12257 5776 12291
rect 5724 12248 5776 12257
rect 9312 12291 9364 12300
rect 9312 12257 9321 12291
rect 9321 12257 9355 12291
rect 9355 12257 9364 12291
rect 9312 12248 9364 12257
rect 10968 12291 11020 12300
rect 10968 12257 10977 12291
rect 10977 12257 11011 12291
rect 11011 12257 11020 12291
rect 10968 12248 11020 12257
rect 13912 12248 13964 12300
rect 19800 12316 19852 12368
rect 14832 12291 14884 12300
rect 14832 12257 14841 12291
rect 14841 12257 14875 12291
rect 14875 12257 14884 12291
rect 14832 12248 14884 12257
rect 16948 12291 17000 12300
rect 16948 12257 16957 12291
rect 16957 12257 16991 12291
rect 16991 12257 17000 12291
rect 16948 12248 17000 12257
rect 19892 12291 19944 12300
rect 19892 12257 19901 12291
rect 19901 12257 19935 12291
rect 19935 12257 19944 12291
rect 19892 12248 19944 12257
rect 20076 12248 20128 12300
rect 23756 12248 23808 12300
rect 26424 12291 26476 12300
rect 26424 12257 26433 12291
rect 26433 12257 26467 12291
rect 26467 12257 26476 12291
rect 26424 12248 26476 12257
rect 26700 12291 26752 12300
rect 26700 12257 26709 12291
rect 26709 12257 26743 12291
rect 26743 12257 26752 12291
rect 26700 12248 26752 12257
rect 4896 12180 4948 12232
rect 8484 12180 8536 12232
rect 9220 12180 9272 12232
rect 11244 12223 11296 12232
rect 11244 12189 11253 12223
rect 11253 12189 11287 12223
rect 11287 12189 11296 12223
rect 11244 12180 11296 12189
rect 4804 12112 4856 12164
rect 6552 12112 6604 12164
rect 10876 12112 10928 12164
rect 13452 12180 13504 12232
rect 14004 12180 14056 12232
rect 15200 12180 15252 12232
rect 15660 12223 15712 12232
rect 15660 12189 15669 12223
rect 15669 12189 15703 12223
rect 15703 12189 15712 12223
rect 15660 12180 15712 12189
rect 20812 12223 20864 12232
rect 16672 12112 16724 12164
rect 20812 12189 20821 12223
rect 20821 12189 20855 12223
rect 20855 12189 20864 12223
rect 20812 12180 20864 12189
rect 23020 12223 23072 12232
rect 23020 12189 23029 12223
rect 23029 12189 23063 12223
rect 23063 12189 23072 12223
rect 23020 12180 23072 12189
rect 23664 12180 23716 12232
rect 26332 12180 26384 12232
rect 27988 12112 28040 12164
rect 7012 12044 7064 12096
rect 9496 12087 9548 12096
rect 9496 12053 9505 12087
rect 9505 12053 9539 12087
rect 9539 12053 9548 12087
rect 9496 12044 9548 12053
rect 11888 12044 11940 12096
rect 12072 12087 12124 12096
rect 12072 12053 12081 12087
rect 12081 12053 12115 12087
rect 12115 12053 12124 12087
rect 12072 12044 12124 12053
rect 12256 12044 12308 12096
rect 25044 12044 25096 12096
rect 7896 11942 7948 11994
rect 7960 11942 8012 11994
rect 8024 11942 8076 11994
rect 8088 11942 8140 11994
rect 8152 11942 8204 11994
rect 14842 11942 14894 11994
rect 14906 11942 14958 11994
rect 14970 11942 15022 11994
rect 15034 11942 15086 11994
rect 15098 11942 15150 11994
rect 21788 11942 21840 11994
rect 21852 11942 21904 11994
rect 21916 11942 21968 11994
rect 21980 11942 22032 11994
rect 22044 11942 22096 11994
rect 28734 11942 28786 11994
rect 28798 11942 28850 11994
rect 28862 11942 28914 11994
rect 28926 11942 28978 11994
rect 28990 11942 29042 11994
rect 6552 11883 6604 11892
rect 6552 11849 6561 11883
rect 6561 11849 6595 11883
rect 6595 11849 6604 11883
rect 6552 11840 6604 11849
rect 7012 11883 7064 11892
rect 7012 11849 7021 11883
rect 7021 11849 7055 11883
rect 7055 11849 7064 11883
rect 7012 11840 7064 11849
rect 11060 11840 11112 11892
rect 12072 11840 12124 11892
rect 9864 11772 9916 11824
rect 2320 11679 2372 11688
rect 2320 11645 2329 11679
rect 2329 11645 2363 11679
rect 2363 11645 2372 11679
rect 2320 11636 2372 11645
rect 4160 11704 4212 11756
rect 6368 11704 6420 11756
rect 9680 11704 9732 11756
rect 10692 11747 10744 11756
rect 10692 11713 10701 11747
rect 10701 11713 10735 11747
rect 10735 11713 10744 11747
rect 10692 11704 10744 11713
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 12256 11772 12308 11824
rect 16764 11840 16816 11892
rect 20076 11840 20128 11892
rect 26332 11840 26384 11892
rect 13728 11815 13780 11824
rect 13728 11781 13737 11815
rect 13737 11781 13771 11815
rect 13771 11781 13780 11815
rect 13728 11772 13780 11781
rect 16580 11772 16632 11824
rect 25044 11815 25096 11824
rect 25044 11781 25053 11815
rect 25053 11781 25087 11815
rect 25087 11781 25096 11815
rect 25044 11772 25096 11781
rect 25688 11772 25740 11824
rect 27988 11815 28040 11824
rect 27988 11781 27997 11815
rect 27997 11781 28031 11815
rect 28031 11781 28040 11815
rect 27988 11772 28040 11781
rect 14648 11704 14700 11756
rect 16672 11704 16724 11756
rect 17132 11747 17184 11756
rect 17132 11713 17166 11747
rect 17166 11713 17184 11747
rect 17132 11704 17184 11713
rect 4252 11679 4304 11688
rect 4252 11645 4261 11679
rect 4261 11645 4295 11679
rect 4295 11645 4304 11679
rect 4252 11636 4304 11645
rect 7196 11679 7248 11688
rect 7196 11645 7205 11679
rect 7205 11645 7239 11679
rect 7239 11645 7248 11679
rect 7196 11636 7248 11645
rect 10784 11679 10836 11688
rect 10784 11645 10793 11679
rect 10793 11645 10827 11679
rect 10827 11645 10836 11679
rect 10784 11636 10836 11645
rect 11980 11679 12032 11688
rect 11980 11645 11989 11679
rect 11989 11645 12023 11679
rect 12023 11645 12032 11679
rect 11980 11636 12032 11645
rect 14740 11636 14792 11688
rect 20168 11704 20220 11756
rect 24676 11704 24728 11756
rect 27344 11704 27396 11756
rect 19892 11636 19944 11688
rect 20628 11679 20680 11688
rect 20628 11645 20637 11679
rect 20637 11645 20671 11679
rect 20671 11645 20680 11679
rect 20628 11636 20680 11645
rect 21272 11636 21324 11688
rect 22468 11636 22520 11688
rect 23664 11636 23716 11688
rect 24768 11679 24820 11688
rect 24768 11645 24777 11679
rect 24777 11645 24811 11679
rect 24811 11645 24820 11679
rect 24768 11636 24820 11645
rect 27528 11636 27580 11688
rect 20904 11568 20956 11620
rect 8484 11500 8536 11552
rect 11796 11500 11848 11552
rect 18144 11500 18196 11552
rect 19340 11543 19392 11552
rect 19340 11509 19349 11543
rect 19349 11509 19383 11543
rect 19383 11509 19392 11543
rect 19340 11500 19392 11509
rect 19524 11500 19576 11552
rect 19892 11500 19944 11552
rect 23940 11543 23992 11552
rect 23940 11509 23949 11543
rect 23949 11509 23983 11543
rect 23983 11509 23992 11543
rect 23940 11500 23992 11509
rect 4423 11398 4475 11450
rect 4487 11398 4539 11450
rect 4551 11398 4603 11450
rect 4615 11398 4667 11450
rect 4679 11398 4731 11450
rect 11369 11398 11421 11450
rect 11433 11398 11485 11450
rect 11497 11398 11549 11450
rect 11561 11398 11613 11450
rect 11625 11398 11677 11450
rect 18315 11398 18367 11450
rect 18379 11398 18431 11450
rect 18443 11398 18495 11450
rect 18507 11398 18559 11450
rect 18571 11398 18623 11450
rect 25261 11398 25313 11450
rect 25325 11398 25377 11450
rect 25389 11398 25441 11450
rect 25453 11398 25505 11450
rect 25517 11398 25569 11450
rect 6368 11296 6420 11348
rect 2964 11228 3016 11280
rect 7012 11228 7064 11280
rect 11980 11296 12032 11348
rect 17132 11339 17184 11348
rect 17132 11305 17141 11339
rect 17141 11305 17175 11339
rect 17175 11305 17184 11339
rect 17132 11296 17184 11305
rect 19616 11339 19668 11348
rect 19616 11305 19625 11339
rect 19625 11305 19659 11339
rect 19659 11305 19668 11339
rect 19616 11296 19668 11305
rect 19892 11339 19944 11348
rect 19892 11305 19901 11339
rect 19901 11305 19935 11339
rect 19935 11305 19944 11339
rect 19892 11296 19944 11305
rect 24768 11339 24820 11348
rect 24768 11305 24777 11339
rect 24777 11305 24811 11339
rect 24811 11305 24820 11339
rect 24768 11296 24820 11305
rect 14188 11228 14240 11280
rect 19708 11228 19760 11280
rect 9036 11160 9088 11212
rect 9220 11203 9272 11212
rect 9220 11169 9229 11203
rect 9229 11169 9263 11203
rect 9263 11169 9272 11203
rect 9220 11160 9272 11169
rect 10232 11160 10284 11212
rect 11060 11160 11112 11212
rect 14740 11203 14792 11212
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 1584 11092 1636 11101
rect 5448 11135 5500 11144
rect 5448 11101 5457 11135
rect 5457 11101 5491 11135
rect 5491 11101 5500 11135
rect 5448 11092 5500 11101
rect 5632 11092 5684 11144
rect 9128 11092 9180 11144
rect 11244 11092 11296 11144
rect 1860 11067 1912 11076
rect 1860 11033 1869 11067
rect 1869 11033 1903 11067
rect 1903 11033 1912 11067
rect 1860 11024 1912 11033
rect 2320 11024 2372 11076
rect 13728 11092 13780 11144
rect 14740 11169 14749 11203
rect 14749 11169 14783 11203
rect 14783 11169 14792 11203
rect 14740 11160 14792 11169
rect 14832 11160 14884 11212
rect 17408 11160 17460 11212
rect 19340 11160 19392 11212
rect 16764 11092 16816 11144
rect 18144 11092 18196 11144
rect 20904 11160 20956 11212
rect 25688 11203 25740 11212
rect 20720 11092 20772 11144
rect 25688 11169 25697 11203
rect 25697 11169 25731 11203
rect 25731 11169 25740 11203
rect 25688 11160 25740 11169
rect 26056 11160 26108 11212
rect 24676 11135 24728 11144
rect 24676 11101 24685 11135
rect 24685 11101 24719 11135
rect 24719 11101 24728 11135
rect 24676 11092 24728 11101
rect 27344 11160 27396 11212
rect 26608 11135 26660 11144
rect 26608 11101 26617 11135
rect 26617 11101 26651 11135
rect 26651 11101 26660 11135
rect 26608 11092 26660 11101
rect 27528 11092 27580 11144
rect 13084 11024 13136 11076
rect 19432 11067 19484 11076
rect 7104 10956 7156 11008
rect 7656 10956 7708 11008
rect 12164 10956 12216 11008
rect 14280 10999 14332 11008
rect 14280 10965 14289 10999
rect 14289 10965 14323 10999
rect 14323 10965 14332 10999
rect 14280 10956 14332 10965
rect 19432 11033 19441 11067
rect 19441 11033 19475 11067
rect 19475 11033 19484 11067
rect 19432 11024 19484 11033
rect 23480 11024 23532 11076
rect 23664 11024 23716 11076
rect 20536 10999 20588 11008
rect 20536 10965 20545 10999
rect 20545 10965 20579 10999
rect 20579 10965 20588 10999
rect 20536 10956 20588 10965
rect 22836 10956 22888 11008
rect 7896 10854 7948 10906
rect 7960 10854 8012 10906
rect 8024 10854 8076 10906
rect 8088 10854 8140 10906
rect 8152 10854 8204 10906
rect 14842 10854 14894 10906
rect 14906 10854 14958 10906
rect 14970 10854 15022 10906
rect 15034 10854 15086 10906
rect 15098 10854 15150 10906
rect 21788 10854 21840 10906
rect 21852 10854 21904 10906
rect 21916 10854 21968 10906
rect 21980 10854 22032 10906
rect 22044 10854 22096 10906
rect 28734 10854 28786 10906
rect 28798 10854 28850 10906
rect 28862 10854 28914 10906
rect 28926 10854 28978 10906
rect 28990 10854 29042 10906
rect 1860 10752 1912 10804
rect 14740 10752 14792 10804
rect 7656 10684 7708 10736
rect 8116 10684 8168 10736
rect 9128 10727 9180 10736
rect 9128 10693 9137 10727
rect 9137 10693 9171 10727
rect 9171 10693 9180 10727
rect 9128 10684 9180 10693
rect 14280 10684 14332 10736
rect 19708 10727 19760 10736
rect 19708 10693 19717 10727
rect 19717 10693 19751 10727
rect 19751 10693 19760 10727
rect 19708 10684 19760 10693
rect 23940 10752 23992 10804
rect 24676 10752 24728 10804
rect 24124 10684 24176 10736
rect 2964 10659 3016 10668
rect 2964 10625 2973 10659
rect 2973 10625 3007 10659
rect 3007 10625 3016 10659
rect 2964 10616 3016 10625
rect 4988 10616 5040 10668
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 14556 10616 14608 10668
rect 17224 10659 17276 10668
rect 17224 10625 17233 10659
rect 17233 10625 17267 10659
rect 17267 10625 17276 10659
rect 17224 10616 17276 10625
rect 4344 10548 4396 10600
rect 17408 10591 17460 10600
rect 17408 10557 17417 10591
rect 17417 10557 17451 10591
rect 17451 10557 17460 10591
rect 20812 10616 20864 10668
rect 22836 10659 22888 10668
rect 22836 10625 22845 10659
rect 22845 10625 22879 10659
rect 22879 10625 22888 10659
rect 22836 10616 22888 10625
rect 27896 10659 27948 10668
rect 27896 10625 27905 10659
rect 27905 10625 27939 10659
rect 27939 10625 27948 10659
rect 27896 10616 27948 10625
rect 21456 10591 21508 10600
rect 17408 10548 17460 10557
rect 17868 10480 17920 10532
rect 5632 10412 5684 10464
rect 16764 10412 16816 10464
rect 20260 10412 20312 10464
rect 21456 10557 21465 10591
rect 21465 10557 21499 10591
rect 21499 10557 21508 10591
rect 21456 10548 21508 10557
rect 21824 10548 21876 10600
rect 28172 10591 28224 10600
rect 28172 10557 28181 10591
rect 28181 10557 28215 10591
rect 28215 10557 28224 10591
rect 28172 10548 28224 10557
rect 23572 10412 23624 10464
rect 4423 10310 4475 10362
rect 4487 10310 4539 10362
rect 4551 10310 4603 10362
rect 4615 10310 4667 10362
rect 4679 10310 4731 10362
rect 11369 10310 11421 10362
rect 11433 10310 11485 10362
rect 11497 10310 11549 10362
rect 11561 10310 11613 10362
rect 11625 10310 11677 10362
rect 18315 10310 18367 10362
rect 18379 10310 18431 10362
rect 18443 10310 18495 10362
rect 18507 10310 18559 10362
rect 18571 10310 18623 10362
rect 25261 10310 25313 10362
rect 25325 10310 25377 10362
rect 25389 10310 25441 10362
rect 25453 10310 25505 10362
rect 25517 10310 25569 10362
rect 1584 10208 1636 10260
rect 9772 10208 9824 10260
rect 2964 10140 3016 10192
rect 4160 10115 4212 10124
rect 4160 10081 4169 10115
rect 4169 10081 4203 10115
rect 4203 10081 4212 10115
rect 4160 10072 4212 10081
rect 2780 10004 2832 10056
rect 4252 10047 4304 10056
rect 4252 10013 4261 10047
rect 4261 10013 4295 10047
rect 4295 10013 4304 10047
rect 4252 10004 4304 10013
rect 9312 10140 9364 10192
rect 4988 10115 5040 10124
rect 4988 10081 4997 10115
rect 4997 10081 5031 10115
rect 5031 10081 5040 10115
rect 4988 10072 5040 10081
rect 6092 10115 6144 10124
rect 6092 10081 6101 10115
rect 6101 10081 6135 10115
rect 6135 10081 6144 10115
rect 6092 10072 6144 10081
rect 8116 10072 8168 10124
rect 5540 9936 5592 9988
rect 12348 10115 12400 10124
rect 12348 10081 12357 10115
rect 12357 10081 12391 10115
rect 12391 10081 12400 10115
rect 12348 10072 12400 10081
rect 12624 10072 12676 10124
rect 10876 9936 10928 9988
rect 14556 10004 14608 10056
rect 16672 10208 16724 10260
rect 17868 10251 17920 10260
rect 17868 10217 17877 10251
rect 17877 10217 17911 10251
rect 17911 10217 17920 10251
rect 17868 10208 17920 10217
rect 19432 10208 19484 10260
rect 20904 10208 20956 10260
rect 20260 10115 20312 10124
rect 20260 10081 20269 10115
rect 20269 10081 20303 10115
rect 20303 10081 20312 10115
rect 20260 10072 20312 10081
rect 20536 10115 20588 10124
rect 20536 10081 20545 10115
rect 20545 10081 20579 10115
rect 20579 10081 20588 10115
rect 20536 10072 20588 10081
rect 26608 10140 26660 10192
rect 27620 10183 27672 10192
rect 27620 10149 27629 10183
rect 27629 10149 27663 10183
rect 27663 10149 27672 10183
rect 27620 10140 27672 10149
rect 24124 10072 24176 10124
rect 26516 10072 26568 10124
rect 16764 10047 16816 10056
rect 16764 10013 16798 10047
rect 16798 10013 16816 10047
rect 16764 10004 16816 10013
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 23020 10047 23072 10056
rect 23020 10013 23029 10047
rect 23029 10013 23063 10047
rect 23063 10013 23072 10047
rect 23020 10004 23072 10013
rect 20812 9936 20864 9988
rect 21272 9936 21324 9988
rect 21824 9936 21876 9988
rect 27620 10004 27672 10056
rect 25964 9936 26016 9988
rect 12164 9911 12216 9920
rect 12164 9877 12173 9911
rect 12173 9877 12207 9911
rect 12207 9877 12216 9911
rect 12164 9868 12216 9877
rect 19340 9868 19392 9920
rect 7896 9766 7948 9818
rect 7960 9766 8012 9818
rect 8024 9766 8076 9818
rect 8088 9766 8140 9818
rect 8152 9766 8204 9818
rect 14842 9766 14894 9818
rect 14906 9766 14958 9818
rect 14970 9766 15022 9818
rect 15034 9766 15086 9818
rect 15098 9766 15150 9818
rect 21788 9766 21840 9818
rect 21852 9766 21904 9818
rect 21916 9766 21968 9818
rect 21980 9766 22032 9818
rect 22044 9766 22096 9818
rect 28734 9766 28786 9818
rect 28798 9766 28850 9818
rect 28862 9766 28914 9818
rect 28926 9766 28978 9818
rect 28990 9766 29042 9818
rect 26516 9707 26568 9716
rect 26516 9673 26525 9707
rect 26525 9673 26559 9707
rect 26559 9673 26568 9707
rect 26516 9664 26568 9673
rect 27620 9707 27672 9716
rect 27620 9673 27629 9707
rect 27629 9673 27663 9707
rect 27663 9673 27672 9707
rect 27620 9664 27672 9673
rect 4344 9596 4396 9648
rect 10600 9639 10652 9648
rect 2780 9571 2832 9580
rect 2780 9537 2789 9571
rect 2789 9537 2823 9571
rect 2823 9537 2832 9571
rect 2780 9528 2832 9537
rect 4068 9528 4120 9580
rect 5632 9528 5684 9580
rect 9588 9571 9640 9580
rect 9588 9537 9597 9571
rect 9597 9537 9631 9571
rect 9631 9537 9640 9571
rect 9588 9528 9640 9537
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 10232 9571 10284 9580
rect 10232 9537 10241 9571
rect 10241 9537 10275 9571
rect 10275 9537 10284 9571
rect 10232 9528 10284 9537
rect 10600 9605 10609 9639
rect 10609 9605 10643 9639
rect 10643 9605 10652 9639
rect 10600 9596 10652 9605
rect 19340 9596 19392 9648
rect 20628 9596 20680 9648
rect 23020 9596 23072 9648
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 10876 9528 10928 9580
rect 14648 9528 14700 9580
rect 15108 9528 15160 9580
rect 18512 9528 18564 9580
rect 20352 9528 20404 9580
rect 4896 9460 4948 9512
rect 10784 9392 10836 9444
rect 18788 9460 18840 9512
rect 19800 9460 19852 9512
rect 26424 9571 26476 9580
rect 26424 9537 26433 9571
rect 26433 9537 26467 9571
rect 26467 9537 26476 9571
rect 26424 9528 26476 9537
rect 26608 9571 26660 9580
rect 26608 9537 26617 9571
rect 26617 9537 26651 9571
rect 26651 9537 26660 9571
rect 26608 9528 26660 9537
rect 20812 9460 20864 9512
rect 27252 9460 27304 9512
rect 2596 9324 2648 9376
rect 14372 9324 14424 9376
rect 17132 9324 17184 9376
rect 27804 9392 27856 9444
rect 20260 9324 20312 9376
rect 4423 9222 4475 9274
rect 4487 9222 4539 9274
rect 4551 9222 4603 9274
rect 4615 9222 4667 9274
rect 4679 9222 4731 9274
rect 11369 9222 11421 9274
rect 11433 9222 11485 9274
rect 11497 9222 11549 9274
rect 11561 9222 11613 9274
rect 11625 9222 11677 9274
rect 18315 9222 18367 9274
rect 18379 9222 18431 9274
rect 18443 9222 18495 9274
rect 18507 9222 18559 9274
rect 18571 9222 18623 9274
rect 25261 9222 25313 9274
rect 25325 9222 25377 9274
rect 25389 9222 25441 9274
rect 25453 9222 25505 9274
rect 25517 9222 25569 9274
rect 10508 9163 10560 9172
rect 10508 9129 10517 9163
rect 10517 9129 10551 9163
rect 10551 9129 10560 9163
rect 10508 9120 10560 9129
rect 18788 9163 18840 9172
rect 18788 9129 18797 9163
rect 18797 9129 18831 9163
rect 18831 9129 18840 9163
rect 18788 9120 18840 9129
rect 26884 9163 26936 9172
rect 26884 9129 26893 9163
rect 26893 9129 26927 9163
rect 26927 9129 26936 9163
rect 26884 9120 26936 9129
rect 10600 9052 10652 9104
rect 2688 9027 2740 9036
rect 2688 8993 2697 9027
rect 2697 8993 2731 9027
rect 2731 8993 2740 9027
rect 2688 8984 2740 8993
rect 4160 8984 4212 9036
rect 5540 8984 5592 9036
rect 7012 9027 7064 9036
rect 7012 8993 7021 9027
rect 7021 8993 7055 9027
rect 7055 8993 7064 9027
rect 7012 8984 7064 8993
rect 7288 9027 7340 9036
rect 7288 8993 7297 9027
rect 7297 8993 7331 9027
rect 7331 8993 7340 9027
rect 7288 8984 7340 8993
rect 2504 8916 2556 8968
rect 4252 8916 4304 8968
rect 6920 8959 6972 8968
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 9404 8916 9456 8968
rect 11520 8984 11572 9036
rect 11704 9027 11756 9036
rect 11704 8993 11713 9027
rect 11713 8993 11747 9027
rect 11747 8993 11756 9027
rect 11704 8984 11756 8993
rect 9772 8916 9824 8968
rect 12164 8916 12216 8968
rect 4068 8848 4120 8900
rect 9588 8848 9640 8900
rect 14188 8916 14240 8968
rect 14648 8916 14700 8968
rect 15108 8916 15160 8968
rect 15844 8916 15896 8968
rect 15384 8891 15436 8900
rect 3332 8780 3384 8832
rect 5448 8780 5500 8832
rect 15384 8857 15393 8891
rect 15393 8857 15427 8891
rect 15427 8857 15436 8891
rect 15384 8848 15436 8857
rect 16672 8848 16724 8900
rect 25780 9052 25832 9104
rect 27436 9052 27488 9104
rect 18696 8959 18748 8968
rect 18696 8925 18705 8959
rect 18705 8925 18739 8959
rect 18739 8925 18748 8959
rect 18696 8916 18748 8925
rect 19800 8984 19852 9036
rect 20352 8984 20404 9036
rect 22284 8984 22336 9036
rect 22744 8984 22796 9036
rect 23848 9027 23900 9036
rect 20168 8916 20220 8968
rect 20260 8916 20312 8968
rect 23848 8993 23857 9027
rect 23857 8993 23891 9027
rect 23891 8993 23900 9027
rect 23848 8984 23900 8993
rect 26608 8984 26660 9036
rect 23664 8959 23716 8968
rect 23664 8925 23673 8959
rect 23673 8925 23707 8959
rect 23707 8925 23716 8959
rect 23664 8916 23716 8925
rect 26424 8916 26476 8968
rect 27252 8959 27304 8968
rect 27252 8925 27261 8959
rect 27261 8925 27295 8959
rect 27295 8925 27304 8959
rect 27252 8916 27304 8925
rect 27804 8916 27856 8968
rect 28356 8891 28408 8900
rect 28356 8857 28365 8891
rect 28365 8857 28399 8891
rect 28399 8857 28408 8891
rect 28356 8848 28408 8857
rect 11060 8823 11112 8832
rect 11060 8789 11069 8823
rect 11069 8789 11103 8823
rect 11103 8789 11112 8823
rect 11060 8780 11112 8789
rect 11520 8823 11572 8832
rect 11520 8789 11529 8823
rect 11529 8789 11563 8823
rect 11563 8789 11572 8823
rect 11520 8780 11572 8789
rect 12164 8780 12216 8832
rect 16856 8780 16908 8832
rect 22836 8823 22888 8832
rect 22836 8789 22845 8823
rect 22845 8789 22879 8823
rect 22879 8789 22888 8823
rect 22836 8780 22888 8789
rect 23112 8780 23164 8832
rect 25136 8780 25188 8832
rect 7896 8678 7948 8730
rect 7960 8678 8012 8730
rect 8024 8678 8076 8730
rect 8088 8678 8140 8730
rect 8152 8678 8204 8730
rect 14842 8678 14894 8730
rect 14906 8678 14958 8730
rect 14970 8678 15022 8730
rect 15034 8678 15086 8730
rect 15098 8678 15150 8730
rect 21788 8678 21840 8730
rect 21852 8678 21904 8730
rect 21916 8678 21968 8730
rect 21980 8678 22032 8730
rect 22044 8678 22096 8730
rect 28734 8678 28786 8730
rect 28798 8678 28850 8730
rect 28862 8678 28914 8730
rect 28926 8678 28978 8730
rect 28990 8678 29042 8730
rect 4068 8619 4120 8628
rect 4068 8585 4077 8619
rect 4077 8585 4111 8619
rect 4111 8585 4120 8619
rect 4068 8576 4120 8585
rect 7012 8576 7064 8628
rect 7748 8576 7800 8628
rect 10876 8619 10928 8628
rect 10876 8585 10885 8619
rect 10885 8585 10919 8619
rect 10919 8585 10928 8619
rect 10876 8576 10928 8585
rect 15844 8619 15896 8628
rect 15844 8585 15853 8619
rect 15853 8585 15887 8619
rect 15887 8585 15896 8619
rect 15844 8576 15896 8585
rect 18696 8576 18748 8628
rect 22836 8576 22888 8628
rect 2596 8551 2648 8560
rect 2596 8517 2605 8551
rect 2605 8517 2639 8551
rect 2639 8517 2648 8551
rect 2596 8508 2648 8517
rect 3332 8508 3384 8560
rect 11520 8508 11572 8560
rect 14372 8551 14424 8560
rect 14372 8517 14381 8551
rect 14381 8517 14415 8551
rect 14415 8517 14424 8551
rect 14372 8508 14424 8517
rect 15384 8508 15436 8560
rect 17132 8551 17184 8560
rect 17132 8517 17141 8551
rect 17141 8517 17175 8551
rect 17175 8517 17184 8551
rect 17132 8508 17184 8517
rect 18144 8508 18196 8560
rect 23112 8551 23164 8560
rect 23112 8517 23121 8551
rect 23121 8517 23155 8551
rect 23155 8517 23164 8551
rect 23112 8508 23164 8517
rect 25136 8576 25188 8628
rect 27896 8576 27948 8628
rect 4988 8440 5040 8492
rect 5724 8440 5776 8492
rect 7380 8440 7432 8492
rect 9404 8440 9456 8492
rect 10784 8440 10836 8492
rect 11796 8440 11848 8492
rect 13636 8483 13688 8492
rect 13636 8449 13645 8483
rect 13645 8449 13679 8483
rect 13679 8449 13688 8483
rect 13636 8440 13688 8449
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 22744 8440 22796 8492
rect 27528 8440 27580 8492
rect 28356 8440 28408 8492
rect 2320 8415 2372 8424
rect 2320 8381 2329 8415
rect 2329 8381 2363 8415
rect 2363 8381 2372 8415
rect 2320 8372 2372 8381
rect 27436 8415 27488 8424
rect 27436 8381 27445 8415
rect 27445 8381 27479 8415
rect 27479 8381 27488 8415
rect 27436 8372 27488 8381
rect 11888 8347 11940 8356
rect 11888 8313 11897 8347
rect 11897 8313 11931 8347
rect 11931 8313 11940 8347
rect 11888 8304 11940 8313
rect 4423 8134 4475 8186
rect 4487 8134 4539 8186
rect 4551 8134 4603 8186
rect 4615 8134 4667 8186
rect 4679 8134 4731 8186
rect 11369 8134 11421 8186
rect 11433 8134 11485 8186
rect 11497 8134 11549 8186
rect 11561 8134 11613 8186
rect 11625 8134 11677 8186
rect 18315 8134 18367 8186
rect 18379 8134 18431 8186
rect 18443 8134 18495 8186
rect 18507 8134 18559 8186
rect 18571 8134 18623 8186
rect 25261 8134 25313 8186
rect 25325 8134 25377 8186
rect 25389 8134 25441 8186
rect 25453 8134 25505 8186
rect 25517 8134 25569 8186
rect 2320 8032 2372 8084
rect 5540 8032 5592 8084
rect 9312 8075 9364 8084
rect 9312 8041 9321 8075
rect 9321 8041 9355 8075
rect 9355 8041 9364 8075
rect 9312 8032 9364 8041
rect 12164 8075 12216 8084
rect 12164 8041 12173 8075
rect 12173 8041 12207 8075
rect 12207 8041 12216 8075
rect 12164 8032 12216 8041
rect 13636 8032 13688 8084
rect 10692 7896 10744 7948
rect 3332 7871 3384 7880
rect 3332 7837 3341 7871
rect 3341 7837 3375 7871
rect 3375 7837 3384 7871
rect 3332 7828 3384 7837
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 9036 7828 9088 7880
rect 10876 7828 10928 7880
rect 11060 7871 11112 7880
rect 11060 7837 11094 7871
rect 11094 7837 11112 7871
rect 11060 7828 11112 7837
rect 15660 8032 15712 8084
rect 27252 8032 27304 8084
rect 27804 8075 27856 8084
rect 27804 8041 27813 8075
rect 27813 8041 27847 8075
rect 27847 8041 27856 8075
rect 27804 8032 27856 8041
rect 14648 7896 14700 7948
rect 13912 7828 13964 7880
rect 16672 7871 16724 7880
rect 16672 7837 16681 7871
rect 16681 7837 16715 7871
rect 16715 7837 16724 7871
rect 16672 7828 16724 7837
rect 18144 7896 18196 7948
rect 19984 7896 20036 7948
rect 21640 7896 21692 7948
rect 22192 7939 22244 7948
rect 22192 7905 22201 7939
rect 22201 7905 22235 7939
rect 22235 7905 22244 7939
rect 22192 7896 22244 7905
rect 19340 7828 19392 7880
rect 24768 7871 24820 7880
rect 24768 7837 24777 7871
rect 24777 7837 24811 7871
rect 24811 7837 24820 7871
rect 24768 7828 24820 7837
rect 6920 7803 6972 7812
rect 6920 7769 6929 7803
rect 6929 7769 6963 7803
rect 6963 7769 6972 7803
rect 6920 7760 6972 7769
rect 9588 7803 9640 7812
rect 9588 7769 9597 7803
rect 9597 7769 9631 7803
rect 9631 7769 9640 7803
rect 9588 7760 9640 7769
rect 15200 7760 15252 7812
rect 21180 7760 21232 7812
rect 22468 7803 22520 7812
rect 22468 7769 22477 7803
rect 22477 7769 22511 7803
rect 22511 7769 22520 7803
rect 22468 7760 22520 7769
rect 25964 7760 26016 7812
rect 27988 7828 28040 7880
rect 2412 7692 2464 7744
rect 9128 7735 9180 7744
rect 9128 7701 9137 7735
rect 9137 7701 9171 7735
rect 9171 7701 9180 7735
rect 9128 7692 9180 7701
rect 22192 7692 22244 7744
rect 25412 7692 25464 7744
rect 25688 7692 25740 7744
rect 26424 7735 26476 7744
rect 26424 7701 26433 7735
rect 26433 7701 26467 7735
rect 26467 7701 26476 7735
rect 26424 7692 26476 7701
rect 26608 7735 26660 7744
rect 26608 7701 26617 7735
rect 26617 7701 26651 7735
rect 26651 7701 26660 7735
rect 26608 7692 26660 7701
rect 27620 7692 27672 7744
rect 7896 7590 7948 7642
rect 7960 7590 8012 7642
rect 8024 7590 8076 7642
rect 8088 7590 8140 7642
rect 8152 7590 8204 7642
rect 14842 7590 14894 7642
rect 14906 7590 14958 7642
rect 14970 7590 15022 7642
rect 15034 7590 15086 7642
rect 15098 7590 15150 7642
rect 21788 7590 21840 7642
rect 21852 7590 21904 7642
rect 21916 7590 21968 7642
rect 21980 7590 22032 7642
rect 22044 7590 22096 7642
rect 28734 7590 28786 7642
rect 28798 7590 28850 7642
rect 28862 7590 28914 7642
rect 28926 7590 28978 7642
rect 28990 7590 29042 7642
rect 3332 7488 3384 7540
rect 7012 7488 7064 7540
rect 7380 7531 7432 7540
rect 7380 7497 7389 7531
rect 7389 7497 7423 7531
rect 7423 7497 7432 7531
rect 7380 7488 7432 7497
rect 7748 7488 7800 7540
rect 9496 7488 9548 7540
rect 19340 7488 19392 7540
rect 20168 7488 20220 7540
rect 21180 7531 21232 7540
rect 21180 7497 21189 7531
rect 21189 7497 21223 7531
rect 21223 7497 21232 7531
rect 21180 7488 21232 7497
rect 22468 7488 22520 7540
rect 23572 7531 23624 7540
rect 23572 7497 23581 7531
rect 23581 7497 23615 7531
rect 23615 7497 23624 7531
rect 23572 7488 23624 7497
rect 25412 7488 25464 7540
rect 2412 7463 2464 7472
rect 2412 7429 2421 7463
rect 2421 7429 2455 7463
rect 2455 7429 2464 7463
rect 2412 7420 2464 7429
rect 3424 7420 3476 7472
rect 4896 7420 4948 7472
rect 4988 7352 5040 7404
rect 15200 7420 15252 7472
rect 19708 7420 19760 7472
rect 25044 7420 25096 7472
rect 26424 7488 26476 7540
rect 26516 7488 26568 7540
rect 27528 7531 27580 7540
rect 27528 7497 27537 7531
rect 27537 7497 27571 7531
rect 27571 7497 27580 7531
rect 27528 7488 27580 7497
rect 14648 7352 14700 7404
rect 22192 7352 22244 7404
rect 22652 7352 22704 7404
rect 25136 7395 25188 7404
rect 25136 7361 25145 7395
rect 25145 7361 25179 7395
rect 25179 7361 25188 7395
rect 25136 7352 25188 7361
rect 25412 7395 25464 7404
rect 25412 7361 25421 7395
rect 25421 7361 25455 7395
rect 25455 7361 25464 7395
rect 25412 7352 25464 7361
rect 26332 7352 26384 7404
rect 26516 7352 26568 7404
rect 27988 7395 28040 7404
rect 2136 7327 2188 7336
rect 2136 7293 2145 7327
rect 2145 7293 2179 7327
rect 2179 7293 2188 7327
rect 2136 7284 2188 7293
rect 7012 7216 7064 7268
rect 9496 7284 9548 7336
rect 10508 7284 10560 7336
rect 11704 7284 11756 7336
rect 13820 7284 13872 7336
rect 14188 7327 14240 7336
rect 14188 7293 14197 7327
rect 14197 7293 14231 7327
rect 14231 7293 14240 7327
rect 14188 7284 14240 7293
rect 23848 7327 23900 7336
rect 23848 7293 23857 7327
rect 23857 7293 23891 7327
rect 23891 7293 23900 7327
rect 23848 7284 23900 7293
rect 12348 7216 12400 7268
rect 27988 7361 27997 7395
rect 27997 7361 28031 7395
rect 28031 7361 28040 7395
rect 27988 7352 28040 7361
rect 25964 7216 26016 7268
rect 5816 7191 5868 7200
rect 5816 7157 5825 7191
rect 5825 7157 5859 7191
rect 5859 7157 5868 7191
rect 5816 7148 5868 7157
rect 10600 7148 10652 7200
rect 25044 7148 25096 7200
rect 26516 7148 26568 7200
rect 28080 7191 28132 7200
rect 28080 7157 28089 7191
rect 28089 7157 28123 7191
rect 28123 7157 28132 7191
rect 28080 7148 28132 7157
rect 4423 7046 4475 7098
rect 4487 7046 4539 7098
rect 4551 7046 4603 7098
rect 4615 7046 4667 7098
rect 4679 7046 4731 7098
rect 11369 7046 11421 7098
rect 11433 7046 11485 7098
rect 11497 7046 11549 7098
rect 11561 7046 11613 7098
rect 11625 7046 11677 7098
rect 18315 7046 18367 7098
rect 18379 7046 18431 7098
rect 18443 7046 18495 7098
rect 18507 7046 18559 7098
rect 18571 7046 18623 7098
rect 25261 7046 25313 7098
rect 25325 7046 25377 7098
rect 25389 7046 25441 7098
rect 25453 7046 25505 7098
rect 25517 7046 25569 7098
rect 4896 6987 4948 6996
rect 4896 6953 4905 6987
rect 4905 6953 4939 6987
rect 4939 6953 4948 6987
rect 4896 6944 4948 6953
rect 7288 6944 7340 6996
rect 27988 6944 28040 6996
rect 2688 6851 2740 6860
rect 2688 6817 2697 6851
rect 2697 6817 2731 6851
rect 2731 6817 2740 6851
rect 2688 6808 2740 6817
rect 3424 6851 3476 6860
rect 3424 6817 3433 6851
rect 3433 6817 3467 6851
rect 3467 6817 3476 6851
rect 3424 6808 3476 6817
rect 2504 6740 2556 6792
rect 5816 6740 5868 6792
rect 6736 6808 6788 6860
rect 7012 6740 7064 6792
rect 9128 6808 9180 6860
rect 10876 6851 10928 6860
rect 10876 6817 10885 6851
rect 10885 6817 10919 6851
rect 10919 6817 10928 6851
rect 10876 6808 10928 6817
rect 12716 6808 12768 6860
rect 6092 6647 6144 6656
rect 6092 6613 6101 6647
rect 6101 6613 6135 6647
rect 6135 6613 6144 6647
rect 6092 6604 6144 6613
rect 6460 6647 6512 6656
rect 6460 6613 6469 6647
rect 6469 6613 6503 6647
rect 6503 6613 6512 6647
rect 6460 6604 6512 6613
rect 6552 6647 6604 6656
rect 6552 6613 6561 6647
rect 6561 6613 6595 6647
rect 6595 6613 6604 6647
rect 7748 6672 7800 6724
rect 9680 6740 9732 6792
rect 10232 6740 10284 6792
rect 10600 6783 10652 6792
rect 10600 6749 10618 6783
rect 10618 6749 10652 6783
rect 10600 6740 10652 6749
rect 11704 6740 11756 6792
rect 14004 6808 14056 6860
rect 17132 6851 17184 6860
rect 17132 6817 17141 6851
rect 17141 6817 17175 6851
rect 17175 6817 17184 6851
rect 17132 6808 17184 6817
rect 13084 6740 13136 6792
rect 19432 6783 19484 6792
rect 11796 6672 11848 6724
rect 6552 6604 6604 6613
rect 9496 6647 9548 6656
rect 9496 6613 9505 6647
rect 9505 6613 9539 6647
rect 9539 6613 9548 6647
rect 9496 6604 9548 6613
rect 12256 6647 12308 6656
rect 12256 6613 12265 6647
rect 12265 6613 12299 6647
rect 12299 6613 12308 6647
rect 12256 6604 12308 6613
rect 12624 6647 12676 6656
rect 12624 6613 12633 6647
rect 12633 6613 12667 6647
rect 12667 6613 12676 6647
rect 12624 6604 12676 6613
rect 12716 6647 12768 6656
rect 12716 6613 12725 6647
rect 12725 6613 12759 6647
rect 12759 6613 12768 6647
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 20720 6740 20772 6792
rect 21640 6740 21692 6792
rect 22652 6783 22704 6792
rect 22652 6749 22661 6783
rect 22661 6749 22695 6783
rect 22695 6749 22704 6783
rect 22652 6740 22704 6749
rect 17592 6672 17644 6724
rect 28080 6740 28132 6792
rect 26424 6672 26476 6724
rect 12716 6604 12768 6613
rect 18144 6604 18196 6656
rect 18512 6604 18564 6656
rect 19524 6647 19576 6656
rect 19524 6613 19533 6647
rect 19533 6613 19567 6647
rect 19567 6613 19576 6647
rect 19524 6604 19576 6613
rect 26608 6604 26660 6656
rect 7896 6502 7948 6554
rect 7960 6502 8012 6554
rect 8024 6502 8076 6554
rect 8088 6502 8140 6554
rect 8152 6502 8204 6554
rect 14842 6502 14894 6554
rect 14906 6502 14958 6554
rect 14970 6502 15022 6554
rect 15034 6502 15086 6554
rect 15098 6502 15150 6554
rect 21788 6502 21840 6554
rect 21852 6502 21904 6554
rect 21916 6502 21968 6554
rect 21980 6502 22032 6554
rect 22044 6502 22096 6554
rect 28734 6502 28786 6554
rect 28798 6502 28850 6554
rect 28862 6502 28914 6554
rect 28926 6502 28978 6554
rect 28990 6502 29042 6554
rect 2136 6400 2188 6452
rect 6460 6400 6512 6452
rect 12624 6400 12676 6452
rect 12716 6400 12768 6452
rect 17592 6443 17644 6452
rect 17592 6409 17601 6443
rect 17601 6409 17635 6443
rect 17635 6409 17644 6443
rect 17592 6400 17644 6409
rect 6552 6332 6604 6384
rect 12256 6332 12308 6384
rect 19432 6400 19484 6452
rect 25044 6400 25096 6452
rect 2596 6264 2648 6316
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 7104 6264 7156 6316
rect 5816 6196 5868 6248
rect 9496 6264 9548 6316
rect 9956 6264 10008 6316
rect 10876 6264 10928 6316
rect 17040 6264 17092 6316
rect 19524 6332 19576 6384
rect 18512 6307 18564 6316
rect 9588 6196 9640 6248
rect 16856 6196 16908 6248
rect 18512 6273 18521 6307
rect 18521 6273 18555 6307
rect 18555 6273 18564 6307
rect 18512 6264 18564 6273
rect 19432 6264 19484 6316
rect 18144 6239 18196 6248
rect 18144 6205 18153 6239
rect 18153 6205 18187 6239
rect 18187 6205 18196 6239
rect 18144 6196 18196 6205
rect 19524 6196 19576 6248
rect 20720 6264 20772 6316
rect 21272 6264 21324 6316
rect 27896 6307 27948 6316
rect 27896 6273 27905 6307
rect 27905 6273 27939 6307
rect 27939 6273 27948 6307
rect 27896 6264 27948 6273
rect 6736 6128 6788 6180
rect 22652 6196 22704 6248
rect 28172 6239 28224 6248
rect 28172 6205 28181 6239
rect 28181 6205 28215 6239
rect 28215 6205 28224 6239
rect 28172 6196 28224 6205
rect 4068 6060 4120 6112
rect 7656 6060 7708 6112
rect 8484 6060 8536 6112
rect 19800 6060 19852 6112
rect 20536 6103 20588 6112
rect 20536 6069 20545 6103
rect 20545 6069 20579 6103
rect 20579 6069 20588 6103
rect 20536 6060 20588 6069
rect 22100 6060 22152 6112
rect 24768 6060 24820 6112
rect 4423 5958 4475 6010
rect 4487 5958 4539 6010
rect 4551 5958 4603 6010
rect 4615 5958 4667 6010
rect 4679 5958 4731 6010
rect 11369 5958 11421 6010
rect 11433 5958 11485 6010
rect 11497 5958 11549 6010
rect 11561 5958 11613 6010
rect 11625 5958 11677 6010
rect 18315 5958 18367 6010
rect 18379 5958 18431 6010
rect 18443 5958 18495 6010
rect 18507 5958 18559 6010
rect 18571 5958 18623 6010
rect 25261 5958 25313 6010
rect 25325 5958 25377 6010
rect 25389 5958 25441 6010
rect 25453 5958 25505 6010
rect 25517 5958 25569 6010
rect 4804 5856 4856 5908
rect 6552 5856 6604 5908
rect 7748 5856 7800 5908
rect 9956 5856 10008 5908
rect 10692 5856 10744 5908
rect 13912 5856 13964 5908
rect 15108 5856 15160 5908
rect 17132 5856 17184 5908
rect 21272 5899 21324 5908
rect 21272 5865 21281 5899
rect 21281 5865 21315 5899
rect 21315 5865 21324 5899
rect 21272 5856 21324 5865
rect 4988 5720 5040 5772
rect 10508 5763 10560 5772
rect 10508 5729 10517 5763
rect 10517 5729 10551 5763
rect 10551 5729 10560 5763
rect 10508 5720 10560 5729
rect 12716 5720 12768 5772
rect 2504 5652 2556 5704
rect 3332 5652 3384 5704
rect 6092 5652 6144 5704
rect 7288 5695 7340 5704
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 8300 5695 8352 5704
rect 8300 5661 8309 5695
rect 8309 5661 8343 5695
rect 8343 5661 8352 5695
rect 8300 5652 8352 5661
rect 8484 5695 8536 5704
rect 8484 5661 8493 5695
rect 8493 5661 8527 5695
rect 8527 5661 8536 5695
rect 8484 5652 8536 5661
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 14556 5720 14608 5772
rect 17040 5720 17092 5772
rect 19800 5763 19852 5772
rect 19800 5729 19809 5763
rect 19809 5729 19843 5763
rect 19843 5729 19852 5763
rect 19800 5720 19852 5729
rect 4160 5584 4212 5636
rect 3424 5559 3476 5568
rect 3424 5525 3433 5559
rect 3433 5525 3467 5559
rect 3467 5525 3476 5559
rect 3424 5516 3476 5525
rect 4344 5516 4396 5568
rect 7564 5627 7616 5636
rect 7564 5593 7573 5627
rect 7573 5593 7607 5627
rect 7607 5593 7616 5627
rect 10232 5627 10284 5636
rect 7564 5584 7616 5593
rect 10232 5593 10241 5627
rect 10241 5593 10275 5627
rect 10275 5593 10284 5627
rect 10232 5584 10284 5593
rect 15108 5652 15160 5704
rect 15752 5695 15804 5704
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 19524 5695 19576 5704
rect 19524 5661 19533 5695
rect 19533 5661 19567 5695
rect 19567 5661 19576 5695
rect 19524 5652 19576 5661
rect 21640 5652 21692 5704
rect 22100 5652 22152 5704
rect 27804 5695 27856 5704
rect 27804 5661 27813 5695
rect 27813 5661 27847 5695
rect 27847 5661 27856 5695
rect 27804 5652 27856 5661
rect 15292 5516 15344 5568
rect 16764 5584 16816 5636
rect 20536 5584 20588 5636
rect 27252 5584 27304 5636
rect 16948 5516 17000 5568
rect 21640 5516 21692 5568
rect 26424 5559 26476 5568
rect 26424 5525 26433 5559
rect 26433 5525 26467 5559
rect 26467 5525 26476 5559
rect 26424 5516 26476 5525
rect 7896 5414 7948 5466
rect 7960 5414 8012 5466
rect 8024 5414 8076 5466
rect 8088 5414 8140 5466
rect 8152 5414 8204 5466
rect 14842 5414 14894 5466
rect 14906 5414 14958 5466
rect 14970 5414 15022 5466
rect 15034 5414 15086 5466
rect 15098 5414 15150 5466
rect 21788 5414 21840 5466
rect 21852 5414 21904 5466
rect 21916 5414 21968 5466
rect 21980 5414 22032 5466
rect 22044 5414 22096 5466
rect 28734 5414 28786 5466
rect 28798 5414 28850 5466
rect 28862 5414 28914 5466
rect 28926 5414 28978 5466
rect 28990 5414 29042 5466
rect 2596 5355 2648 5364
rect 2596 5321 2605 5355
rect 2605 5321 2639 5355
rect 2639 5321 2648 5355
rect 2596 5312 2648 5321
rect 7288 5312 7340 5364
rect 7564 5312 7616 5364
rect 15752 5355 15804 5364
rect 15752 5321 15761 5355
rect 15761 5321 15795 5355
rect 15795 5321 15804 5355
rect 15752 5312 15804 5321
rect 16764 5312 16816 5364
rect 25688 5312 25740 5364
rect 27252 5355 27304 5364
rect 27252 5321 27261 5355
rect 27261 5321 27295 5355
rect 27295 5321 27304 5355
rect 27252 5312 27304 5321
rect 27804 5312 27856 5364
rect 3424 5244 3476 5296
rect 4068 5287 4120 5296
rect 4068 5253 4077 5287
rect 4077 5253 4111 5287
rect 4111 5253 4120 5287
rect 4068 5244 4120 5253
rect 8484 5244 8536 5296
rect 15292 5244 15344 5296
rect 4344 5219 4396 5228
rect 4344 5185 4353 5219
rect 4353 5185 4387 5219
rect 4387 5185 4396 5219
rect 4344 5176 4396 5185
rect 6552 5176 6604 5228
rect 5540 5108 5592 5160
rect 6828 5108 6880 5160
rect 8300 5176 8352 5228
rect 16856 5219 16908 5228
rect 16856 5185 16865 5219
rect 16865 5185 16899 5219
rect 16899 5185 16908 5219
rect 16856 5176 16908 5185
rect 17040 5219 17092 5228
rect 17040 5185 17049 5219
rect 17049 5185 17083 5219
rect 17083 5185 17092 5219
rect 17040 5176 17092 5185
rect 21548 5176 21600 5228
rect 22192 5219 22244 5228
rect 22192 5185 22201 5219
rect 22201 5185 22235 5219
rect 22235 5185 22244 5219
rect 26424 5244 26476 5296
rect 22192 5176 22244 5185
rect 26148 5176 26200 5228
rect 26332 5219 26384 5228
rect 26332 5185 26341 5219
rect 26341 5185 26375 5219
rect 26375 5185 26384 5219
rect 26332 5176 26384 5185
rect 27528 5176 27580 5228
rect 13912 5108 13964 5160
rect 14280 5151 14332 5160
rect 14280 5117 14289 5151
rect 14289 5117 14323 5151
rect 14323 5117 14332 5151
rect 14280 5108 14332 5117
rect 25964 5151 26016 5160
rect 25964 5117 25973 5151
rect 25973 5117 26007 5151
rect 26007 5117 26016 5151
rect 25964 5108 26016 5117
rect 22284 4972 22336 5024
rect 22744 5015 22796 5024
rect 22744 4981 22753 5015
rect 22753 4981 22787 5015
rect 22787 4981 22796 5015
rect 22744 4972 22796 4981
rect 26700 4972 26752 5024
rect 4423 4870 4475 4922
rect 4487 4870 4539 4922
rect 4551 4870 4603 4922
rect 4615 4870 4667 4922
rect 4679 4870 4731 4922
rect 11369 4870 11421 4922
rect 11433 4870 11485 4922
rect 11497 4870 11549 4922
rect 11561 4870 11613 4922
rect 11625 4870 11677 4922
rect 18315 4870 18367 4922
rect 18379 4870 18431 4922
rect 18443 4870 18495 4922
rect 18507 4870 18559 4922
rect 18571 4870 18623 4922
rect 25261 4870 25313 4922
rect 25325 4870 25377 4922
rect 25389 4870 25441 4922
rect 25453 4870 25505 4922
rect 25517 4870 25569 4922
rect 26332 4768 26384 4820
rect 27252 4768 27304 4820
rect 27436 4768 27488 4820
rect 27896 4811 27948 4820
rect 27896 4777 27905 4811
rect 27905 4777 27939 4811
rect 27939 4777 27948 4811
rect 27896 4768 27948 4777
rect 4160 4632 4212 4684
rect 6828 4632 6880 4684
rect 6736 4607 6788 4616
rect 6736 4573 6745 4607
rect 6745 4573 6779 4607
rect 6779 4573 6788 4607
rect 6736 4564 6788 4573
rect 8300 4564 8352 4616
rect 11060 4632 11112 4684
rect 21272 4632 21324 4684
rect 28264 4675 28316 4684
rect 28264 4641 28273 4675
rect 28273 4641 28307 4675
rect 28307 4641 28316 4675
rect 28264 4632 28316 4641
rect 10692 4607 10744 4616
rect 6644 4496 6696 4548
rect 9772 4496 9824 4548
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 13820 4564 13872 4616
rect 19524 4564 19576 4616
rect 20628 4564 20680 4616
rect 22652 4607 22704 4616
rect 22652 4573 22661 4607
rect 22661 4573 22695 4607
rect 22695 4573 22704 4607
rect 22652 4564 22704 4573
rect 23296 4564 23348 4616
rect 25964 4564 26016 4616
rect 26240 4564 26292 4616
rect 10600 4496 10652 4548
rect 13636 4496 13688 4548
rect 21640 4496 21692 4548
rect 22928 4539 22980 4548
rect 22928 4505 22962 4539
rect 22962 4505 22980 4539
rect 22928 4496 22980 4505
rect 25596 4496 25648 4548
rect 27712 4564 27764 4616
rect 27436 4496 27488 4548
rect 4344 4428 4396 4480
rect 7380 4471 7432 4480
rect 7380 4437 7389 4471
rect 7389 4437 7423 4471
rect 7423 4437 7432 4471
rect 7380 4428 7432 4437
rect 8392 4428 8444 4480
rect 9680 4428 9732 4480
rect 11704 4428 11756 4480
rect 22192 4428 22244 4480
rect 25688 4471 25740 4480
rect 25688 4437 25697 4471
rect 25697 4437 25731 4471
rect 25731 4437 25740 4471
rect 25688 4428 25740 4437
rect 25964 4428 26016 4480
rect 26700 4471 26752 4480
rect 26700 4437 26709 4471
rect 26709 4437 26743 4471
rect 26743 4437 26752 4471
rect 26700 4428 26752 4437
rect 28356 4428 28408 4480
rect 7896 4326 7948 4378
rect 7960 4326 8012 4378
rect 8024 4326 8076 4378
rect 8088 4326 8140 4378
rect 8152 4326 8204 4378
rect 14842 4326 14894 4378
rect 14906 4326 14958 4378
rect 14970 4326 15022 4378
rect 15034 4326 15086 4378
rect 15098 4326 15150 4378
rect 21788 4326 21840 4378
rect 21852 4326 21904 4378
rect 21916 4326 21968 4378
rect 21980 4326 22032 4378
rect 22044 4326 22096 4378
rect 28734 4326 28786 4378
rect 28798 4326 28850 4378
rect 28862 4326 28914 4378
rect 28926 4326 28978 4378
rect 28990 4326 29042 4378
rect 6736 4224 6788 4276
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 4344 4156 4396 4208
rect 5080 4156 5132 4208
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6644 4088 6696 4097
rect 6828 4088 6880 4140
rect 10600 4224 10652 4276
rect 11060 4267 11112 4276
rect 11060 4233 11069 4267
rect 11069 4233 11103 4267
rect 11103 4233 11112 4267
rect 11060 4224 11112 4233
rect 27712 4267 27764 4276
rect 10876 4156 10928 4208
rect 13636 4156 13688 4208
rect 25688 4156 25740 4208
rect 27712 4233 27721 4267
rect 27721 4233 27755 4267
rect 27755 4233 27764 4267
rect 27712 4224 27764 4233
rect 28264 4267 28316 4276
rect 28264 4233 28273 4267
rect 28273 4233 28307 4267
rect 28307 4233 28316 4267
rect 28264 4224 28316 4233
rect 11060 4088 11112 4140
rect 12164 4088 12216 4140
rect 17224 4131 17276 4140
rect 17224 4097 17233 4131
rect 17233 4097 17267 4131
rect 17267 4097 17276 4131
rect 17224 4088 17276 4097
rect 19984 4088 20036 4140
rect 24676 4088 24728 4140
rect 25596 4131 25648 4140
rect 25596 4097 25605 4131
rect 25605 4097 25639 4131
rect 25639 4097 25648 4131
rect 25596 4088 25648 4097
rect 25964 4131 26016 4140
rect 25964 4097 25973 4131
rect 25973 4097 26007 4131
rect 26007 4097 26016 4131
rect 26240 4131 26292 4140
rect 25964 4088 26016 4097
rect 26240 4097 26249 4131
rect 26249 4097 26283 4131
rect 26283 4097 26292 4131
rect 26240 4088 26292 4097
rect 27252 4088 27304 4140
rect 27528 4131 27580 4140
rect 27528 4097 27537 4131
rect 27537 4097 27571 4131
rect 27571 4097 27580 4131
rect 27528 4088 27580 4097
rect 28356 4131 28408 4140
rect 28356 4097 28365 4131
rect 28365 4097 28399 4131
rect 28399 4097 28408 4131
rect 28356 4088 28408 4097
rect 8300 4063 8352 4072
rect 8300 4029 8309 4063
rect 8309 4029 8343 4063
rect 8343 4029 8352 4063
rect 8300 4020 8352 4029
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 9680 4020 9732 4072
rect 12624 4020 12676 4072
rect 14004 4020 14056 4072
rect 14280 4020 14332 4072
rect 16120 4020 16172 4072
rect 20628 4020 20680 4072
rect 3332 3884 3384 3936
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 7012 3884 7064 3936
rect 9772 3884 9824 3936
rect 12256 3884 12308 3936
rect 14648 3884 14700 3936
rect 19708 3884 19760 3936
rect 19800 3884 19852 3936
rect 26148 4020 26200 4072
rect 25596 3884 25648 3936
rect 27160 3884 27212 3936
rect 4423 3782 4475 3834
rect 4487 3782 4539 3834
rect 4551 3782 4603 3834
rect 4615 3782 4667 3834
rect 4679 3782 4731 3834
rect 11369 3782 11421 3834
rect 11433 3782 11485 3834
rect 11497 3782 11549 3834
rect 11561 3782 11613 3834
rect 11625 3782 11677 3834
rect 18315 3782 18367 3834
rect 18379 3782 18431 3834
rect 18443 3782 18495 3834
rect 18507 3782 18559 3834
rect 18571 3782 18623 3834
rect 25261 3782 25313 3834
rect 25325 3782 25377 3834
rect 25389 3782 25441 3834
rect 25453 3782 25505 3834
rect 25517 3782 25569 3834
rect 6644 3680 6696 3732
rect 4160 3587 4212 3596
rect 4160 3553 4169 3587
rect 4169 3553 4203 3587
rect 4203 3553 4212 3587
rect 4160 3544 4212 3553
rect 2504 3476 2556 3528
rect 6736 3612 6788 3664
rect 9312 3680 9364 3732
rect 9404 3612 9456 3664
rect 5080 3587 5132 3596
rect 5080 3553 5089 3587
rect 5089 3553 5123 3587
rect 5123 3553 5132 3587
rect 5080 3544 5132 3553
rect 7012 3587 7064 3596
rect 7012 3553 7021 3587
rect 7021 3553 7055 3587
rect 7055 3553 7064 3587
rect 7012 3544 7064 3553
rect 6184 3383 6236 3392
rect 6184 3349 6193 3383
rect 6193 3349 6227 3383
rect 6227 3349 6236 3383
rect 6184 3340 6236 3349
rect 8300 3476 8352 3528
rect 11060 3680 11112 3732
rect 11888 3680 11940 3732
rect 16120 3723 16172 3732
rect 16120 3689 16129 3723
rect 16129 3689 16163 3723
rect 16163 3689 16172 3723
rect 16120 3680 16172 3689
rect 19800 3680 19852 3732
rect 19984 3723 20036 3732
rect 19984 3689 19993 3723
rect 19993 3689 20027 3723
rect 20027 3689 20036 3723
rect 19984 3680 20036 3689
rect 22928 3680 22980 3732
rect 24676 3723 24728 3732
rect 24676 3689 24685 3723
rect 24685 3689 24719 3723
rect 24719 3689 24728 3723
rect 24676 3680 24728 3689
rect 26148 3680 26200 3732
rect 12256 3587 12308 3596
rect 12256 3553 12265 3587
rect 12265 3553 12299 3587
rect 12299 3553 12308 3587
rect 12256 3544 12308 3553
rect 16580 3587 16632 3596
rect 16580 3553 16589 3587
rect 16589 3553 16623 3587
rect 16623 3553 16632 3587
rect 19524 3587 19576 3596
rect 16580 3544 16632 3553
rect 19524 3553 19533 3587
rect 19533 3553 19567 3587
rect 19567 3553 19576 3587
rect 19524 3544 19576 3553
rect 22192 3544 22244 3596
rect 12624 3476 12676 3528
rect 13728 3476 13780 3528
rect 13912 3476 13964 3528
rect 16304 3476 16356 3528
rect 17224 3476 17276 3528
rect 19616 3519 19668 3528
rect 19616 3485 19625 3519
rect 19625 3485 19659 3519
rect 19659 3485 19668 3519
rect 19616 3476 19668 3485
rect 20628 3476 20680 3528
rect 25596 3476 25648 3528
rect 27252 3519 27304 3528
rect 27252 3485 27261 3519
rect 27261 3485 27295 3519
rect 27295 3485 27304 3519
rect 27252 3476 27304 3485
rect 27528 3476 27580 3528
rect 7288 3408 7340 3460
rect 11704 3408 11756 3460
rect 22284 3408 22336 3460
rect 7104 3340 7156 3392
rect 14740 3340 14792 3392
rect 17960 3383 18012 3392
rect 17960 3349 17969 3383
rect 17969 3349 18003 3383
rect 18003 3349 18012 3383
rect 17960 3340 18012 3349
rect 7896 3238 7948 3290
rect 7960 3238 8012 3290
rect 8024 3238 8076 3290
rect 8088 3238 8140 3290
rect 8152 3238 8204 3290
rect 14842 3238 14894 3290
rect 14906 3238 14958 3290
rect 14970 3238 15022 3290
rect 15034 3238 15086 3290
rect 15098 3238 15150 3290
rect 21788 3238 21840 3290
rect 21852 3238 21904 3290
rect 21916 3238 21968 3290
rect 21980 3238 22032 3290
rect 22044 3238 22096 3290
rect 28734 3238 28786 3290
rect 28798 3238 28850 3290
rect 28862 3238 28914 3290
rect 28926 3238 28978 3290
rect 28990 3238 29042 3290
rect 6184 3136 6236 3188
rect 10876 3179 10928 3188
rect 4160 3068 4212 3120
rect 7380 3068 7432 3120
rect 10876 3145 10885 3179
rect 10885 3145 10919 3179
rect 10919 3145 10928 3179
rect 10876 3136 10928 3145
rect 14004 3179 14056 3188
rect 14004 3145 14013 3179
rect 14013 3145 14047 3179
rect 14047 3145 14056 3179
rect 14004 3136 14056 3145
rect 14740 3136 14792 3188
rect 19524 3136 19576 3188
rect 19616 3136 19668 3188
rect 17960 3068 18012 3120
rect 8392 3043 8444 3052
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 9772 3000 9824 3052
rect 10692 3000 10744 3052
rect 12440 3000 12492 3052
rect 22744 3068 22796 3120
rect 25964 3136 26016 3188
rect 27252 3136 27304 3188
rect 6920 2932 6972 2984
rect 12624 2975 12676 2984
rect 12624 2941 12633 2975
rect 12633 2941 12667 2975
rect 12667 2941 12676 2975
rect 12624 2932 12676 2941
rect 16304 2975 16356 2984
rect 16304 2941 16313 2975
rect 16313 2941 16347 2975
rect 16347 2941 16356 2975
rect 16304 2932 16356 2941
rect 20628 3000 20680 3052
rect 25596 3000 25648 3052
rect 27160 3043 27212 3052
rect 27160 3009 27169 3043
rect 27169 3009 27203 3043
rect 27203 3009 27212 3043
rect 27160 3000 27212 3009
rect 27436 3000 27488 3052
rect 19708 2975 19760 2984
rect 7104 2864 7156 2916
rect 19708 2941 19717 2975
rect 19717 2941 19751 2975
rect 19751 2941 19760 2975
rect 19708 2932 19760 2941
rect 22928 2932 22980 2984
rect 23296 2932 23348 2984
rect 20628 2796 20680 2848
rect 27896 2796 27948 2848
rect 4423 2694 4475 2746
rect 4487 2694 4539 2746
rect 4551 2694 4603 2746
rect 4615 2694 4667 2746
rect 4679 2694 4731 2746
rect 11369 2694 11421 2746
rect 11433 2694 11485 2746
rect 11497 2694 11549 2746
rect 11561 2694 11613 2746
rect 11625 2694 11677 2746
rect 18315 2694 18367 2746
rect 18379 2694 18431 2746
rect 18443 2694 18495 2746
rect 18507 2694 18559 2746
rect 18571 2694 18623 2746
rect 25261 2694 25313 2746
rect 25325 2694 25377 2746
rect 25389 2694 25441 2746
rect 25453 2694 25505 2746
rect 25517 2694 25569 2746
rect 7288 2635 7340 2644
rect 7288 2601 7297 2635
rect 7297 2601 7331 2635
rect 7331 2601 7340 2635
rect 7288 2592 7340 2601
rect 12440 2592 12492 2644
rect 13728 2499 13780 2508
rect 13728 2465 13737 2499
rect 13737 2465 13771 2499
rect 13771 2465 13780 2499
rect 13728 2456 13780 2465
rect 7104 2388 7156 2440
rect 27896 2431 27948 2440
rect 27896 2397 27905 2431
rect 27905 2397 27939 2431
rect 27939 2397 27948 2431
rect 27896 2388 27948 2397
rect 14648 2320 14700 2372
rect 28172 2363 28224 2372
rect 28172 2329 28181 2363
rect 28181 2329 28215 2363
rect 28215 2329 28224 2363
rect 28172 2320 28224 2329
rect 7896 2150 7948 2202
rect 7960 2150 8012 2202
rect 8024 2150 8076 2202
rect 8088 2150 8140 2202
rect 8152 2150 8204 2202
rect 14842 2150 14894 2202
rect 14906 2150 14958 2202
rect 14970 2150 15022 2202
rect 15034 2150 15086 2202
rect 15098 2150 15150 2202
rect 21788 2150 21840 2202
rect 21852 2150 21904 2202
rect 21916 2150 21968 2202
rect 21980 2150 22032 2202
rect 22044 2150 22096 2202
rect 28734 2150 28786 2202
rect 28798 2150 28850 2202
rect 28862 2150 28914 2202
rect 28926 2150 28978 2202
rect 28990 2150 29042 2202
<< metal2 >>
rect 2042 29200 2098 30000
rect 5722 29200 5778 30000
rect 9402 29322 9458 30000
rect 9402 29294 9628 29322
rect 9402 29200 9458 29294
rect 2056 24886 2084 29200
rect 4423 27772 4731 27781
rect 4423 27770 4429 27772
rect 4485 27770 4509 27772
rect 4565 27770 4589 27772
rect 4645 27770 4669 27772
rect 4725 27770 4731 27772
rect 4485 27718 4487 27770
rect 4667 27718 4669 27770
rect 4423 27716 4429 27718
rect 4485 27716 4509 27718
rect 4565 27716 4589 27718
rect 4645 27716 4669 27718
rect 4725 27716 4731 27718
rect 4423 27707 4731 27716
rect 5736 27470 5764 29200
rect 9600 27470 9628 29294
rect 13082 29200 13138 30000
rect 16762 29322 16818 30000
rect 20442 29322 20498 30000
rect 16762 29294 17080 29322
rect 16762 29200 16818 29294
rect 11369 27772 11677 27781
rect 11369 27770 11375 27772
rect 11431 27770 11455 27772
rect 11511 27770 11535 27772
rect 11591 27770 11615 27772
rect 11671 27770 11677 27772
rect 11431 27718 11433 27770
rect 11613 27718 11615 27770
rect 11369 27716 11375 27718
rect 11431 27716 11455 27718
rect 11511 27716 11535 27718
rect 11591 27716 11615 27718
rect 11671 27716 11677 27718
rect 11369 27707 11677 27716
rect 13096 27470 13124 29200
rect 17052 27470 17080 29294
rect 20442 29294 20668 29322
rect 20442 29200 20498 29294
rect 18315 27772 18623 27781
rect 18315 27770 18321 27772
rect 18377 27770 18401 27772
rect 18457 27770 18481 27772
rect 18537 27770 18561 27772
rect 18617 27770 18623 27772
rect 18377 27718 18379 27770
rect 18559 27718 18561 27770
rect 18315 27716 18321 27718
rect 18377 27716 18401 27718
rect 18457 27716 18481 27718
rect 18537 27716 18561 27718
rect 18617 27716 18623 27718
rect 18315 27707 18623 27716
rect 17684 27532 17736 27538
rect 17684 27474 17736 27480
rect 3332 27464 3384 27470
rect 3332 27406 3384 27412
rect 5724 27464 5776 27470
rect 5724 27406 5776 27412
rect 9588 27464 9640 27470
rect 9588 27406 9640 27412
rect 13084 27464 13136 27470
rect 13084 27406 13136 27412
rect 17040 27464 17092 27470
rect 17040 27406 17092 27412
rect 3148 27328 3200 27334
rect 3148 27270 3200 27276
rect 2872 26988 2924 26994
rect 2872 26930 2924 26936
rect 2884 26602 2912 26930
rect 2792 26574 2912 26602
rect 2136 26240 2188 26246
rect 2136 26182 2188 26188
rect 2148 25906 2176 26182
rect 2792 26042 2820 26574
rect 2872 26376 2924 26382
rect 2872 26318 2924 26324
rect 2780 26036 2832 26042
rect 2780 25978 2832 25984
rect 2136 25900 2188 25906
rect 2136 25842 2188 25848
rect 2884 25838 2912 26318
rect 3160 26314 3188 27270
rect 3344 26314 3372 27406
rect 4528 27396 4580 27402
rect 4528 27338 4580 27344
rect 12624 27396 12676 27402
rect 12624 27338 12676 27344
rect 13728 27396 13780 27402
rect 13728 27338 13780 27344
rect 4540 27062 4568 27338
rect 6920 27328 6972 27334
rect 6920 27270 6972 27276
rect 3424 27056 3476 27062
rect 3424 26998 3476 27004
rect 4528 27056 4580 27062
rect 4528 26998 4580 27004
rect 5264 27056 5316 27062
rect 5264 26998 5316 27004
rect 3436 26450 3464 26998
rect 4160 26784 4212 26790
rect 4160 26726 4212 26732
rect 4172 26586 4200 26726
rect 4423 26684 4731 26693
rect 4423 26682 4429 26684
rect 4485 26682 4509 26684
rect 4565 26682 4589 26684
rect 4645 26682 4669 26684
rect 4725 26682 4731 26684
rect 4485 26630 4487 26682
rect 4667 26630 4669 26682
rect 4423 26628 4429 26630
rect 4485 26628 4509 26630
rect 4565 26628 4589 26630
rect 4645 26628 4669 26630
rect 4725 26628 4731 26630
rect 4423 26619 4731 26628
rect 4160 26580 4212 26586
rect 4160 26522 4212 26528
rect 3424 26444 3476 26450
rect 3424 26386 3476 26392
rect 3148 26308 3200 26314
rect 3148 26250 3200 26256
rect 3332 26308 3384 26314
rect 3332 26250 3384 26256
rect 2872 25832 2924 25838
rect 2872 25774 2924 25780
rect 2044 24880 2096 24886
rect 2044 24822 2096 24828
rect 2884 24750 2912 25774
rect 4172 25702 4200 26522
rect 4988 26512 5040 26518
rect 4988 26454 5040 26460
rect 4436 26308 4488 26314
rect 4436 26250 4488 26256
rect 4344 26240 4396 26246
rect 4344 26182 4396 26188
rect 4356 25922 4384 26182
rect 4448 26042 4476 26250
rect 4896 26240 4948 26246
rect 4896 26182 4948 26188
rect 4436 26036 4488 26042
rect 4436 25978 4488 25984
rect 4264 25906 4384 25922
rect 4264 25900 4396 25906
rect 4264 25894 4344 25900
rect 4160 25696 4212 25702
rect 4160 25638 4212 25644
rect 4172 25378 4200 25638
rect 4264 25498 4292 25894
rect 4344 25842 4396 25848
rect 4448 25786 4476 25978
rect 4356 25758 4476 25786
rect 4804 25832 4856 25838
rect 4804 25774 4856 25780
rect 4252 25492 4304 25498
rect 4252 25434 4304 25440
rect 4172 25350 4292 25378
rect 3148 25288 3200 25294
rect 3148 25230 3200 25236
rect 4160 25288 4212 25294
rect 4160 25230 4212 25236
rect 2964 25152 3016 25158
rect 2964 25094 3016 25100
rect 2976 24818 3004 25094
rect 2964 24812 3016 24818
rect 2964 24754 3016 24760
rect 2872 24744 2924 24750
rect 2872 24686 2924 24692
rect 2780 24200 2832 24206
rect 2780 24142 2832 24148
rect 2792 23254 2820 24142
rect 2884 23866 2912 24686
rect 3160 24410 3188 25230
rect 4068 25152 4120 25158
rect 4068 25094 4120 25100
rect 3976 24880 4028 24886
rect 3976 24822 4028 24828
rect 3148 24404 3200 24410
rect 3148 24346 3200 24352
rect 3884 24064 3936 24070
rect 3884 24006 3936 24012
rect 2872 23860 2924 23866
rect 2872 23802 2924 23808
rect 2780 23248 2832 23254
rect 2780 23190 2832 23196
rect 2228 23112 2280 23118
rect 2228 23054 2280 23060
rect 3056 23112 3108 23118
rect 3056 23054 3108 23060
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 2044 22568 2096 22574
rect 2044 22510 2096 22516
rect 2056 22030 2084 22510
rect 2044 22024 2096 22030
rect 2044 21966 2096 21972
rect 2056 20806 2084 21966
rect 2240 21622 2268 23054
rect 2780 22976 2832 22982
rect 2780 22918 2832 22924
rect 2792 22030 2820 22918
rect 3068 22030 3096 23054
rect 3436 22710 3464 23054
rect 3424 22704 3476 22710
rect 3424 22646 3476 22652
rect 3436 22234 3464 22646
rect 3700 22636 3752 22642
rect 3700 22578 3752 22584
rect 3424 22228 3476 22234
rect 3424 22170 3476 22176
rect 2780 22024 2832 22030
rect 2780 21966 2832 21972
rect 3056 22024 3108 22030
rect 3056 21966 3108 21972
rect 3712 21690 3740 22578
rect 3700 21684 3752 21690
rect 3700 21626 3752 21632
rect 2228 21616 2280 21622
rect 2228 21558 2280 21564
rect 3148 21616 3200 21622
rect 3148 21558 3200 21564
rect 2780 21344 2832 21350
rect 2780 21286 2832 21292
rect 2044 20800 2096 20806
rect 2044 20742 2096 20748
rect 2056 20398 2084 20742
rect 2792 20534 2820 21286
rect 2780 20528 2832 20534
rect 2780 20470 2832 20476
rect 2044 20392 2096 20398
rect 2044 20334 2096 20340
rect 2056 19854 2084 20334
rect 3160 20262 3188 21558
rect 3896 21554 3924 24006
rect 3988 23118 4016 24822
rect 4080 24206 4108 25094
rect 4172 24954 4200 25230
rect 4264 25158 4292 25350
rect 4356 25294 4384 25758
rect 4423 25596 4731 25605
rect 4423 25594 4429 25596
rect 4485 25594 4509 25596
rect 4565 25594 4589 25596
rect 4645 25594 4669 25596
rect 4725 25594 4731 25596
rect 4485 25542 4487 25594
rect 4667 25542 4669 25594
rect 4423 25540 4429 25542
rect 4485 25540 4509 25542
rect 4565 25540 4589 25542
rect 4645 25540 4669 25542
rect 4725 25540 4731 25542
rect 4423 25531 4731 25540
rect 4816 25498 4844 25774
rect 4804 25492 4856 25498
rect 4804 25434 4856 25440
rect 4344 25288 4396 25294
rect 4344 25230 4396 25236
rect 4908 25226 4936 26182
rect 5000 25906 5028 26454
rect 5080 26376 5132 26382
rect 5080 26318 5132 26324
rect 4988 25900 5040 25906
rect 4988 25842 5040 25848
rect 5092 25362 5120 26318
rect 5276 25838 5304 26998
rect 6932 26994 6960 27270
rect 7896 27228 8204 27237
rect 7896 27226 7902 27228
rect 7958 27226 7982 27228
rect 8038 27226 8062 27228
rect 8118 27226 8142 27228
rect 8198 27226 8204 27228
rect 7958 27174 7960 27226
rect 8140 27174 8142 27226
rect 7896 27172 7902 27174
rect 7958 27172 7982 27174
rect 8038 27172 8062 27174
rect 8118 27172 8142 27174
rect 8198 27172 8204 27174
rect 7896 27163 8204 27172
rect 6920 26988 6972 26994
rect 6920 26930 6972 26936
rect 8300 26988 8352 26994
rect 8300 26930 8352 26936
rect 9496 26988 9548 26994
rect 9496 26930 9548 26936
rect 10416 26988 10468 26994
rect 10416 26930 10468 26936
rect 12256 26988 12308 26994
rect 12256 26930 12308 26936
rect 6552 26784 6604 26790
rect 6552 26726 6604 26732
rect 6564 26450 6592 26726
rect 6552 26444 6604 26450
rect 6552 26386 6604 26392
rect 6276 26376 6328 26382
rect 6276 26318 6328 26324
rect 5264 25832 5316 25838
rect 5264 25774 5316 25780
rect 5080 25356 5132 25362
rect 5080 25298 5132 25304
rect 5276 25226 5304 25774
rect 6288 25498 6316 26318
rect 6644 25832 6696 25838
rect 6644 25774 6696 25780
rect 6276 25492 6328 25498
rect 6276 25434 6328 25440
rect 6368 25288 6420 25294
rect 6368 25230 6420 25236
rect 4896 25220 4948 25226
rect 4896 25162 4948 25168
rect 5264 25220 5316 25226
rect 5264 25162 5316 25168
rect 4252 25152 4304 25158
rect 4252 25094 4304 25100
rect 4160 24948 4212 24954
rect 4160 24890 4212 24896
rect 4423 24508 4731 24517
rect 4423 24506 4429 24508
rect 4485 24506 4509 24508
rect 4565 24506 4589 24508
rect 4645 24506 4669 24508
rect 4725 24506 4731 24508
rect 4485 24454 4487 24506
rect 4667 24454 4669 24506
rect 4423 24452 4429 24454
rect 4485 24452 4509 24454
rect 4565 24452 4589 24454
rect 4645 24452 4669 24454
rect 4725 24452 4731 24454
rect 4423 24443 4731 24452
rect 5276 24274 5304 25162
rect 5264 24268 5316 24274
rect 5264 24210 5316 24216
rect 6380 24206 6408 25230
rect 4068 24200 4120 24206
rect 4068 24142 4120 24148
rect 6368 24200 6420 24206
rect 6368 24142 6420 24148
rect 4080 23322 4108 24142
rect 4252 24132 4304 24138
rect 4252 24074 4304 24080
rect 4068 23316 4120 23322
rect 4068 23258 4120 23264
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 4080 22794 4108 23258
rect 4080 22778 4200 22794
rect 4080 22772 4212 22778
rect 4080 22766 4160 22772
rect 4160 22714 4212 22720
rect 4172 22522 4200 22714
rect 4264 22642 4292 24074
rect 6380 23866 6408 24142
rect 6368 23860 6420 23866
rect 6368 23802 6420 23808
rect 4344 23724 4396 23730
rect 4344 23666 4396 23672
rect 4356 22982 4384 23666
rect 6552 23656 6604 23662
rect 6552 23598 6604 23604
rect 4423 23420 4731 23429
rect 4423 23418 4429 23420
rect 4485 23418 4509 23420
rect 4565 23418 4589 23420
rect 4645 23418 4669 23420
rect 4725 23418 4731 23420
rect 4485 23366 4487 23418
rect 4667 23366 4669 23418
rect 4423 23364 4429 23366
rect 4485 23364 4509 23366
rect 4565 23364 4589 23366
rect 4645 23364 4669 23366
rect 4725 23364 4731 23366
rect 4423 23355 4731 23364
rect 5816 23112 5868 23118
rect 5816 23054 5868 23060
rect 6460 23112 6512 23118
rect 6460 23054 6512 23060
rect 4344 22976 4396 22982
rect 4344 22918 4396 22924
rect 4252 22636 4304 22642
rect 4252 22578 4304 22584
rect 4172 22494 4292 22522
rect 4160 22432 4212 22438
rect 4160 22374 4212 22380
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 3884 21548 3936 21554
rect 3884 21490 3936 21496
rect 4080 21486 4108 21966
rect 4172 21554 4200 22374
rect 4264 22030 4292 22494
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 3240 21480 3292 21486
rect 3240 21422 3292 21428
rect 4068 21480 4120 21486
rect 4068 21422 4120 21428
rect 3252 20602 3280 21422
rect 4356 20942 4384 22918
rect 4804 22500 4856 22506
rect 4804 22442 4856 22448
rect 4423 22332 4731 22341
rect 4423 22330 4429 22332
rect 4485 22330 4509 22332
rect 4565 22330 4589 22332
rect 4645 22330 4669 22332
rect 4725 22330 4731 22332
rect 4485 22278 4487 22330
rect 4667 22278 4669 22330
rect 4423 22276 4429 22278
rect 4485 22276 4509 22278
rect 4565 22276 4589 22278
rect 4645 22276 4669 22278
rect 4725 22276 4731 22278
rect 4423 22267 4731 22276
rect 4816 22094 4844 22442
rect 5828 22094 5856 23054
rect 6368 22976 6420 22982
rect 6368 22918 6420 22924
rect 6380 22642 6408 22918
rect 6368 22636 6420 22642
rect 6368 22578 6420 22584
rect 6472 22098 6500 23054
rect 6564 22778 6592 23598
rect 6656 23186 6684 25774
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 6840 23798 6868 24006
rect 6828 23792 6880 23798
rect 6828 23734 6880 23740
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 6736 22976 6788 22982
rect 6736 22918 6788 22924
rect 6552 22772 6604 22778
rect 6552 22714 6604 22720
rect 4816 22066 4936 22094
rect 4804 21616 4856 21622
rect 4804 21558 4856 21564
rect 4423 21244 4731 21253
rect 4423 21242 4429 21244
rect 4485 21242 4509 21244
rect 4565 21242 4589 21244
rect 4645 21242 4669 21244
rect 4725 21242 4731 21244
rect 4485 21190 4487 21242
rect 4667 21190 4669 21242
rect 4423 21188 4429 21190
rect 4485 21188 4509 21190
rect 4565 21188 4589 21190
rect 4645 21188 4669 21190
rect 4725 21188 4731 21190
rect 4423 21179 4731 21188
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 3240 20596 3292 20602
rect 3240 20538 3292 20544
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 3240 20392 3292 20398
rect 3240 20334 3292 20340
rect 3148 20256 3200 20262
rect 3148 20198 3200 20204
rect 2044 19848 2096 19854
rect 2044 19790 2096 19796
rect 2056 18834 2084 19790
rect 2780 19780 2832 19786
rect 2780 19722 2832 19728
rect 2792 19310 2820 19722
rect 3160 19514 3188 20198
rect 3148 19508 3200 19514
rect 3148 19450 3200 19456
rect 3160 19310 3188 19450
rect 3252 19310 3280 20334
rect 2780 19304 2832 19310
rect 2780 19246 2832 19252
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 3240 19304 3292 19310
rect 3240 19246 3292 19252
rect 2044 18828 2096 18834
rect 2044 18770 2096 18776
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2884 18358 2912 18702
rect 2872 18352 2924 18358
rect 2872 18294 2924 18300
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 2884 17882 2912 18022
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 3252 17678 3280 19246
rect 4264 19174 4292 20402
rect 4816 20346 4844 21558
rect 4908 21350 4936 22066
rect 5552 22066 5856 22094
rect 6460 22092 6512 22098
rect 5552 22030 5580 22066
rect 6460 22034 6512 22040
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5816 22024 5868 22030
rect 5816 21966 5868 21972
rect 4896 21344 4948 21350
rect 4896 21286 4948 21292
rect 4908 20466 4936 21286
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 4816 20318 4936 20346
rect 4423 20156 4731 20165
rect 4423 20154 4429 20156
rect 4485 20154 4509 20156
rect 4565 20154 4589 20156
rect 4645 20154 4669 20156
rect 4725 20154 4731 20156
rect 4485 20102 4487 20154
rect 4667 20102 4669 20154
rect 4423 20100 4429 20102
rect 4485 20100 4509 20102
rect 4565 20100 4589 20102
rect 4645 20100 4669 20102
rect 4725 20100 4731 20102
rect 4423 20091 4731 20100
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 4356 19446 4384 19654
rect 4344 19440 4396 19446
rect 4344 19382 4396 19388
rect 4908 19378 4936 20318
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4423 19068 4731 19077
rect 4423 19066 4429 19068
rect 4485 19066 4509 19068
rect 4565 19066 4589 19068
rect 4645 19066 4669 19068
rect 4725 19066 4731 19068
rect 4485 19014 4487 19066
rect 4667 19014 4669 19066
rect 4423 19012 4429 19014
rect 4485 19012 4509 19014
rect 4565 19012 4589 19014
rect 4645 19012 4669 19014
rect 4725 19012 4731 19014
rect 4423 19003 4731 19012
rect 4344 18692 4396 18698
rect 4344 18634 4396 18640
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 3988 17882 4016 18226
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 2976 17202 3004 17614
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2320 16992 2372 16998
rect 2320 16934 2372 16940
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 2056 16114 2084 16390
rect 2332 16182 2360 16934
rect 3252 16590 3280 17614
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 2596 16584 2648 16590
rect 2596 16526 2648 16532
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 2320 16176 2372 16182
rect 2320 16118 2372 16124
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 2608 15502 2636 16526
rect 3252 15502 3280 16526
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3344 16182 3372 16390
rect 4080 16182 4108 17138
rect 3332 16176 3384 16182
rect 3332 16118 3384 16124
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 4356 15570 4384 18634
rect 4423 17980 4731 17989
rect 4423 17978 4429 17980
rect 4485 17978 4509 17980
rect 4565 17978 4589 17980
rect 4645 17978 4669 17980
rect 4725 17978 4731 17980
rect 4485 17926 4487 17978
rect 4667 17926 4669 17978
rect 4423 17924 4429 17926
rect 4485 17924 4509 17926
rect 4565 17924 4589 17926
rect 4645 17924 4669 17926
rect 4725 17924 4731 17926
rect 4423 17915 4731 17924
rect 4423 16892 4731 16901
rect 4423 16890 4429 16892
rect 4485 16890 4509 16892
rect 4565 16890 4589 16892
rect 4645 16890 4669 16892
rect 4725 16890 4731 16892
rect 4485 16838 4487 16890
rect 4667 16838 4669 16890
rect 4423 16836 4429 16838
rect 4485 16836 4509 16838
rect 4565 16836 4589 16838
rect 4645 16836 4669 16838
rect 4725 16836 4731 16838
rect 4423 16827 4731 16836
rect 4423 15804 4731 15813
rect 4423 15802 4429 15804
rect 4485 15802 4509 15804
rect 4565 15802 4589 15804
rect 4645 15802 4669 15804
rect 4725 15802 4731 15804
rect 4485 15750 4487 15802
rect 4667 15750 4669 15802
rect 4423 15748 4429 15750
rect 4485 15748 4509 15750
rect 4565 15748 4589 15750
rect 4645 15748 4669 15750
rect 4725 15748 4731 15750
rect 4423 15739 4731 15748
rect 4344 15564 4396 15570
rect 4344 15506 4396 15512
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 2504 15360 2556 15366
rect 2504 15302 2556 15308
rect 1872 15026 1900 15302
rect 2516 15094 2544 15302
rect 2504 15088 2556 15094
rect 2504 15030 2556 15036
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 2608 14958 2636 15438
rect 2780 15428 2832 15434
rect 2780 15370 2832 15376
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2792 14414 2820 15370
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3252 15094 3280 15302
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 4423 14716 4731 14725
rect 4423 14714 4429 14716
rect 4485 14714 4509 14716
rect 4565 14714 4589 14716
rect 4645 14714 4669 14716
rect 4725 14714 4731 14716
rect 4485 14662 4487 14714
rect 4667 14662 4669 14714
rect 4423 14660 4429 14662
rect 4485 14660 4509 14662
rect 4565 14660 4589 14662
rect 4645 14660 4669 14662
rect 4725 14660 4731 14662
rect 4423 14651 4731 14660
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 1584 14272 1636 14278
rect 1584 14214 1636 14220
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 1596 12850 1624 14214
rect 2332 14006 2360 14214
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 2792 13870 2820 14350
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2056 13530 2084 13806
rect 2044 13524 2096 13530
rect 2044 13466 2096 13472
rect 3068 13326 3096 14350
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3344 14006 3372 14214
rect 3332 14000 3384 14006
rect 3332 13942 3384 13948
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 4423 13628 4731 13637
rect 4423 13626 4429 13628
rect 4485 13626 4509 13628
rect 4565 13626 4589 13628
rect 4645 13626 4669 13628
rect 4725 13626 4731 13628
rect 4485 13574 4487 13626
rect 4667 13574 4669 13626
rect 4423 13572 4429 13574
rect 4485 13572 4509 13574
rect 4565 13572 4589 13574
rect 4645 13572 4669 13574
rect 4725 13572 4731 13574
rect 4423 13563 4731 13572
rect 4816 13394 4844 13874
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 3608 13252 3660 13258
rect 3608 13194 3660 13200
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 1872 12918 1900 13126
rect 1860 12912 1912 12918
rect 1860 12854 1912 12860
rect 2976 12850 3004 13126
rect 3620 12918 3648 13194
rect 3608 12912 3660 12918
rect 3608 12854 3660 12860
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4423 12540 4731 12549
rect 4423 12538 4429 12540
rect 4485 12538 4509 12540
rect 4565 12538 4589 12540
rect 4645 12538 4669 12540
rect 4725 12538 4731 12540
rect 4485 12486 4487 12538
rect 4667 12486 4669 12538
rect 4423 12484 4429 12486
rect 4485 12484 4509 12486
rect 4565 12484 4589 12486
rect 4645 12484 4669 12486
rect 4725 12484 4731 12486
rect 4423 12475 4731 12484
rect 4816 12170 4844 12786
rect 4908 12238 4936 19314
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 5092 15026 5120 19110
rect 5552 18902 5580 21966
rect 5632 21344 5684 21350
rect 5632 21286 5684 21292
rect 5644 20874 5672 21286
rect 5724 21004 5776 21010
rect 5724 20946 5776 20952
rect 5632 20868 5684 20874
rect 5632 20810 5684 20816
rect 5736 20602 5764 20946
rect 5724 20596 5776 20602
rect 5724 20538 5776 20544
rect 5540 18896 5592 18902
rect 5540 18838 5592 18844
rect 5828 18766 5856 21966
rect 6368 21956 6420 21962
rect 6368 21898 6420 21904
rect 6380 20874 6408 21898
rect 6748 21554 6776 22918
rect 6932 22094 6960 26930
rect 8312 26450 8340 26930
rect 8760 26920 8812 26926
rect 8760 26862 8812 26868
rect 8392 26784 8444 26790
rect 8392 26726 8444 26732
rect 8300 26444 8352 26450
rect 8300 26386 8352 26392
rect 7656 26376 7708 26382
rect 7656 26318 7708 26324
rect 7668 25974 7696 26318
rect 7896 26140 8204 26149
rect 7896 26138 7902 26140
rect 7958 26138 7982 26140
rect 8038 26138 8062 26140
rect 8118 26138 8142 26140
rect 8198 26138 8204 26140
rect 7958 26086 7960 26138
rect 8140 26086 8142 26138
rect 7896 26084 7902 26086
rect 7958 26084 7982 26086
rect 8038 26084 8062 26086
rect 8118 26084 8142 26086
rect 8198 26084 8204 26086
rect 7896 26075 8204 26084
rect 7656 25968 7708 25974
rect 7656 25910 7708 25916
rect 8404 25906 8432 26726
rect 8772 26586 8800 26862
rect 8760 26580 8812 26586
rect 8760 26522 8812 26528
rect 8668 26240 8720 26246
rect 8668 26182 8720 26188
rect 8680 25974 8708 26182
rect 8668 25968 8720 25974
rect 8668 25910 8720 25916
rect 8392 25900 8444 25906
rect 8392 25842 8444 25848
rect 8772 25838 8800 26522
rect 9312 26444 9364 26450
rect 9312 26386 9364 26392
rect 8760 25832 8812 25838
rect 8760 25774 8812 25780
rect 7748 25356 7800 25362
rect 7748 25298 7800 25304
rect 7472 25220 7524 25226
rect 7472 25162 7524 25168
rect 7104 25152 7156 25158
rect 7104 25094 7156 25100
rect 7116 22642 7144 25094
rect 7484 24954 7512 25162
rect 7760 24954 7788 25298
rect 9324 25294 9352 26386
rect 9508 26042 9536 26930
rect 9680 26920 9732 26926
rect 9680 26862 9732 26868
rect 9496 26036 9548 26042
rect 9496 25978 9548 25984
rect 9312 25288 9364 25294
rect 9312 25230 9364 25236
rect 9508 25226 9536 25978
rect 9692 25974 9720 26862
rect 9864 26580 9916 26586
rect 9864 26522 9916 26528
rect 9680 25968 9732 25974
rect 9680 25910 9732 25916
rect 9496 25220 9548 25226
rect 9496 25162 9548 25168
rect 7896 25052 8204 25061
rect 7896 25050 7902 25052
rect 7958 25050 7982 25052
rect 8038 25050 8062 25052
rect 8118 25050 8142 25052
rect 8198 25050 8204 25052
rect 7958 24998 7960 25050
rect 8140 24998 8142 25050
rect 7896 24996 7902 24998
rect 7958 24996 7982 24998
rect 8038 24996 8062 24998
rect 8118 24996 8142 24998
rect 8198 24996 8204 24998
rect 7896 24987 8204 24996
rect 7472 24948 7524 24954
rect 7472 24890 7524 24896
rect 7748 24948 7800 24954
rect 7748 24890 7800 24896
rect 9496 24880 9548 24886
rect 9496 24822 9548 24828
rect 7748 24744 7800 24750
rect 7748 24686 7800 24692
rect 7288 23792 7340 23798
rect 7288 23734 7340 23740
rect 7300 23186 7328 23734
rect 7288 23180 7340 23186
rect 7288 23122 7340 23128
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 6932 22066 7052 22094
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 6748 21146 6776 21490
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6368 20868 6420 20874
rect 6368 20810 6420 20816
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 5908 19780 5960 19786
rect 5908 19722 5960 19728
rect 5920 19514 5948 19722
rect 5908 19508 5960 19514
rect 5908 19450 5960 19456
rect 6012 19378 6040 20402
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6656 19514 6684 19790
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 5908 18828 5960 18834
rect 5908 18770 5960 18776
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5828 18358 5856 18702
rect 5816 18352 5868 18358
rect 5816 18294 5868 18300
rect 5828 17202 5856 18294
rect 5920 17202 5948 18770
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 6368 17604 6420 17610
rect 6368 17546 6420 17552
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 5552 16454 5580 17002
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5080 15020 5132 15026
rect 5080 14962 5132 14968
rect 5552 14550 5580 15438
rect 5736 15434 5764 16934
rect 5828 16114 5856 17138
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5724 15428 5776 15434
rect 5724 15370 5776 15376
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 5092 13258 5120 14214
rect 5552 14074 5580 14350
rect 5908 14340 5960 14346
rect 5908 14282 5960 14288
rect 5920 14074 5948 14282
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 5828 13394 5856 13806
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 6092 12912 6144 12918
rect 6092 12854 6144 12860
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1596 10266 1624 11086
rect 2332 11082 2360 11630
rect 2964 11280 3016 11286
rect 2964 11222 3016 11228
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 2320 11076 2372 11082
rect 2320 11018 2372 11024
rect 1872 10810 1900 11018
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 2976 10674 3004 11222
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 2976 10198 3004 10610
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 4172 10130 4200 11698
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2792 9586 2820 9998
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2332 8090 2360 8366
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 7478 2452 7686
rect 2412 7472 2464 7478
rect 2412 7414 2464 7420
rect 2136 7336 2188 7342
rect 2136 7278 2188 7284
rect 2148 6458 2176 7278
rect 2516 6798 2544 8910
rect 2608 8566 2636 9318
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 2700 6866 2728 8978
rect 4080 8906 4108 9522
rect 4172 9042 4200 10066
rect 4264 10062 4292 11630
rect 4423 11452 4731 11461
rect 4423 11450 4429 11452
rect 4485 11450 4509 11452
rect 4565 11450 4589 11452
rect 4645 11450 4669 11452
rect 4725 11450 4731 11452
rect 4485 11398 4487 11450
rect 4667 11398 4669 11450
rect 4423 11396 4429 11398
rect 4485 11396 4509 11398
rect 4565 11396 4589 11398
rect 4645 11396 4669 11398
rect 4725 11396 4731 11398
rect 4423 11387 4731 11396
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4264 8974 4292 9998
rect 4356 9654 4384 10542
rect 4423 10364 4731 10373
rect 4423 10362 4429 10364
rect 4485 10362 4509 10364
rect 4565 10362 4589 10364
rect 4645 10362 4669 10364
rect 4725 10362 4731 10364
rect 4485 10310 4487 10362
rect 4667 10310 4669 10362
rect 4423 10308 4429 10310
rect 4485 10308 4509 10310
rect 4565 10308 4589 10310
rect 4645 10308 4669 10310
rect 4725 10308 4731 10310
rect 4423 10299 4731 10308
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4423 9276 4731 9285
rect 4423 9274 4429 9276
rect 4485 9274 4509 9276
rect 4565 9274 4589 9276
rect 4645 9274 4669 9276
rect 4725 9274 4731 9276
rect 4485 9222 4487 9274
rect 4667 9222 4669 9274
rect 4423 9220 4429 9222
rect 4485 9220 4509 9222
rect 4565 9220 4589 9222
rect 4645 9220 4669 9222
rect 4725 9220 4731 9222
rect 4423 9211 4731 9220
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3344 8566 3372 8774
rect 4080 8634 4108 8842
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 4423 8188 4731 8197
rect 4423 8186 4429 8188
rect 4485 8186 4509 8188
rect 4565 8186 4589 8188
rect 4645 8186 4669 8188
rect 4725 8186 4731 8188
rect 4485 8134 4487 8186
rect 4667 8134 4669 8186
rect 4423 8132 4429 8134
rect 4485 8132 4509 8134
rect 4565 8132 4589 8134
rect 4645 8132 4669 8134
rect 4725 8132 4731 8134
rect 4423 8123 4731 8132
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3344 7546 3372 7822
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3436 6866 3464 7414
rect 4423 7100 4731 7109
rect 4423 7098 4429 7100
rect 4485 7098 4509 7100
rect 4565 7098 4589 7100
rect 4645 7098 4669 7100
rect 4725 7098 4731 7100
rect 4485 7046 4487 7098
rect 4667 7046 4669 7098
rect 4423 7044 4429 7046
rect 4485 7044 4509 7046
rect 4565 7044 4589 7046
rect 4645 7044 4669 7046
rect 4725 7044 4731 7046
rect 4423 7035 4731 7044
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2516 5710 2544 6734
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2516 3534 2544 5646
rect 2608 5370 2636 6258
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 3344 4146 3372 5646
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3436 5302 3464 5510
rect 4080 5302 4108 6054
rect 4423 6012 4731 6021
rect 4423 6010 4429 6012
rect 4485 6010 4509 6012
rect 4565 6010 4589 6012
rect 4645 6010 4669 6012
rect 4725 6010 4731 6012
rect 4485 5958 4487 6010
rect 4667 5958 4669 6010
rect 4423 5956 4429 5958
rect 4485 5956 4509 5958
rect 4565 5956 4589 5958
rect 4645 5956 4669 5958
rect 4725 5956 4731 5958
rect 4423 5947 4731 5956
rect 4816 5914 4844 12106
rect 4908 9518 4936 12174
rect 5460 11150 5488 12582
rect 5736 12306 5764 12786
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 5000 10130 5028 10610
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 5460 8838 5488 11086
rect 5644 10470 5672 11086
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5552 9042 5580 9930
rect 5644 9586 5672 10406
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 4908 7002 4936 7414
rect 5000 7410 5028 8434
rect 5552 8090 5580 8978
rect 5736 8498 5764 12242
rect 6104 10130 6132 12854
rect 6380 11762 6408 17546
rect 6564 16658 6592 18022
rect 6748 17678 6776 18226
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 6748 17338 6776 17614
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6736 17332 6788 17338
rect 6736 17274 6788 17280
rect 6840 16658 6868 17478
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 7024 16454 7052 22066
rect 7116 20398 7144 22578
rect 7668 22234 7696 22578
rect 7656 22228 7708 22234
rect 7656 22170 7708 22176
rect 7760 22166 7788 24686
rect 9404 24200 9456 24206
rect 9404 24142 9456 24148
rect 7896 23964 8204 23973
rect 7896 23962 7902 23964
rect 7958 23962 7982 23964
rect 8038 23962 8062 23964
rect 8118 23962 8142 23964
rect 8198 23962 8204 23964
rect 7958 23910 7960 23962
rect 8140 23910 8142 23962
rect 7896 23908 7902 23910
rect 7958 23908 7982 23910
rect 8038 23908 8062 23910
rect 8118 23908 8142 23910
rect 8198 23908 8204 23910
rect 7896 23899 8204 23908
rect 7840 23860 7892 23866
rect 7840 23802 7892 23808
rect 7852 23118 7880 23802
rect 8208 23180 8260 23186
rect 8208 23122 8260 23128
rect 7840 23112 7892 23118
rect 7840 23054 7892 23060
rect 8220 22964 8248 23122
rect 8220 22936 8340 22964
rect 7896 22876 8204 22885
rect 7896 22874 7902 22876
rect 7958 22874 7982 22876
rect 8038 22874 8062 22876
rect 8118 22874 8142 22876
rect 8198 22874 8204 22876
rect 7958 22822 7960 22874
rect 8140 22822 8142 22874
rect 7896 22820 7902 22822
rect 7958 22820 7982 22822
rect 8038 22820 8062 22822
rect 8118 22820 8142 22822
rect 8198 22820 8204 22822
rect 7896 22811 8204 22820
rect 8312 22778 8340 22936
rect 8300 22772 8352 22778
rect 8220 22732 8300 22760
rect 7748 22160 7800 22166
rect 7748 22102 7800 22108
rect 8220 22098 8248 22732
rect 8300 22714 8352 22720
rect 9416 22642 9444 24142
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 8208 22092 8260 22098
rect 8208 22034 8260 22040
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 7896 21788 8204 21797
rect 7896 21786 7902 21788
rect 7958 21786 7982 21788
rect 8038 21786 8062 21788
rect 8118 21786 8142 21788
rect 8198 21786 8204 21788
rect 7958 21734 7960 21786
rect 8140 21734 8142 21786
rect 7896 21732 7902 21734
rect 7958 21732 7982 21734
rect 8038 21732 8062 21734
rect 8118 21732 8142 21734
rect 8198 21732 8204 21734
rect 7896 21723 8204 21732
rect 9416 21146 9444 21830
rect 9404 21140 9456 21146
rect 9404 21082 9456 21088
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7668 20466 7696 20878
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 7116 19446 7144 20334
rect 7564 20256 7616 20262
rect 7564 20198 7616 20204
rect 7472 19780 7524 19786
rect 7472 19722 7524 19728
rect 7104 19440 7156 19446
rect 7104 19382 7156 19388
rect 7116 19310 7144 19382
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7484 18834 7512 19722
rect 7576 19446 7604 20198
rect 7668 20058 7696 20402
rect 7760 20398 7788 20946
rect 7896 20700 8204 20709
rect 7896 20698 7902 20700
rect 7958 20698 7982 20700
rect 8038 20698 8062 20700
rect 8118 20698 8142 20700
rect 8198 20698 8204 20700
rect 7958 20646 7960 20698
rect 8140 20646 8142 20698
rect 7896 20644 7902 20646
rect 7958 20644 7982 20646
rect 8038 20644 8062 20646
rect 8118 20644 8142 20646
rect 8198 20644 8204 20646
rect 7896 20635 8204 20644
rect 9416 20482 9444 21082
rect 9232 20454 9444 20482
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7760 19514 7788 20334
rect 7896 19612 8204 19621
rect 7896 19610 7902 19612
rect 7958 19610 7982 19612
rect 8038 19610 8062 19612
rect 8118 19610 8142 19612
rect 8198 19610 8204 19612
rect 7958 19558 7960 19610
rect 8140 19558 8142 19610
rect 7896 19556 7902 19558
rect 7958 19556 7982 19558
rect 8038 19556 8062 19558
rect 8118 19556 8142 19558
rect 8198 19556 8204 19558
rect 7896 19547 8204 19556
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7564 19440 7616 19446
rect 7564 19382 7616 19388
rect 7656 19440 7708 19446
rect 7656 19382 7708 19388
rect 7564 19168 7616 19174
rect 7668 19122 7696 19382
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 7616 19116 7696 19122
rect 7564 19110 7696 19116
rect 7576 19094 7696 19110
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6564 15434 6592 15982
rect 7300 15706 7328 17614
rect 7380 17604 7432 17610
rect 7380 17546 7432 17552
rect 7392 17134 7420 17546
rect 7668 17202 7696 19094
rect 7896 18524 8204 18533
rect 7896 18522 7902 18524
rect 7958 18522 7982 18524
rect 8038 18522 8062 18524
rect 8118 18522 8142 18524
rect 8198 18522 8204 18524
rect 7958 18470 7960 18522
rect 8140 18470 8142 18522
rect 7896 18468 7902 18470
rect 7958 18468 7982 18470
rect 8038 18468 8062 18470
rect 8118 18468 8142 18470
rect 8198 18468 8204 18470
rect 7896 18459 8204 18468
rect 8312 17746 8340 19314
rect 9232 19258 9260 20454
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9324 19378 9352 19790
rect 9416 19394 9444 20334
rect 9508 19514 9536 24822
rect 9772 23180 9824 23186
rect 9772 23122 9824 23128
rect 9680 22636 9732 22642
rect 9680 22578 9732 22584
rect 9588 21956 9640 21962
rect 9588 21898 9640 21904
rect 9600 20874 9628 21898
rect 9692 21690 9720 22578
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9588 20868 9640 20874
rect 9588 20810 9640 20816
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9312 19372 9364 19378
rect 9416 19366 9536 19394
rect 9312 19314 9364 19320
rect 9508 19310 9536 19366
rect 9496 19304 9548 19310
rect 9232 19230 9352 19258
rect 9496 19246 9548 19252
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9232 18766 9260 19110
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 7896 17436 8204 17445
rect 7896 17434 7902 17436
rect 7958 17434 7982 17436
rect 8038 17434 8062 17436
rect 8118 17434 8142 17436
rect 8198 17434 8204 17436
rect 7958 17382 7960 17434
rect 8140 17382 8142 17434
rect 7896 17380 7902 17382
rect 7958 17380 7982 17382
rect 8038 17380 8062 17382
rect 8118 17380 8142 17382
rect 8198 17380 8204 17382
rect 7896 17371 8204 17380
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7392 16046 7420 17070
rect 8312 16794 8340 17682
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 9220 16516 9272 16522
rect 9220 16458 9272 16464
rect 7896 16348 8204 16357
rect 7896 16346 7902 16348
rect 7958 16346 7982 16348
rect 8038 16346 8062 16348
rect 8118 16346 8142 16348
rect 8198 16346 8204 16348
rect 7958 16294 7960 16346
rect 8140 16294 8142 16346
rect 7896 16292 7902 16294
rect 7958 16292 7982 16294
rect 8038 16292 8062 16294
rect 8118 16292 8142 16294
rect 8198 16292 8204 16294
rect 7896 16283 8204 16292
rect 9232 16250 9260 16458
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9324 16182 9352 19230
rect 9508 18170 9536 19246
rect 9600 18358 9628 20810
rect 9692 20262 9720 20946
rect 9784 20398 9812 23122
rect 9876 21894 9904 26522
rect 10428 26382 10456 26930
rect 10508 26784 10560 26790
rect 10508 26726 10560 26732
rect 10784 26784 10836 26790
rect 10784 26726 10836 26732
rect 10520 26450 10548 26726
rect 10796 26450 10824 26726
rect 11369 26684 11677 26693
rect 11369 26682 11375 26684
rect 11431 26682 11455 26684
rect 11511 26682 11535 26684
rect 11591 26682 11615 26684
rect 11671 26682 11677 26684
rect 11431 26630 11433 26682
rect 11613 26630 11615 26682
rect 11369 26628 11375 26630
rect 11431 26628 11455 26630
rect 11511 26628 11535 26630
rect 11591 26628 11615 26630
rect 11671 26628 11677 26630
rect 11369 26619 11677 26628
rect 10508 26444 10560 26450
rect 10508 26386 10560 26392
rect 10784 26444 10836 26450
rect 10784 26386 10836 26392
rect 10140 26376 10192 26382
rect 10140 26318 10192 26324
rect 10416 26376 10468 26382
rect 10416 26318 10468 26324
rect 10152 26042 10180 26318
rect 11796 26308 11848 26314
rect 11796 26250 11848 26256
rect 10140 26036 10192 26042
rect 10140 25978 10192 25984
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 9772 20392 9824 20398
rect 9772 20334 9824 20340
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9876 20058 9904 20402
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9784 19378 9812 19858
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9784 18970 9812 19314
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9588 18352 9640 18358
rect 9588 18294 9640 18300
rect 9508 18142 9628 18170
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9416 16402 9444 17682
rect 9496 16448 9548 16454
rect 9416 16396 9496 16402
rect 9416 16390 9548 16396
rect 9416 16374 9536 16390
rect 9416 16250 9444 16374
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9312 16176 9364 16182
rect 9312 16118 9364 16124
rect 9600 16046 9628 18142
rect 9968 17542 9996 25230
rect 10152 21690 10180 25978
rect 11369 25596 11677 25605
rect 11369 25594 11375 25596
rect 11431 25594 11455 25596
rect 11511 25594 11535 25596
rect 11591 25594 11615 25596
rect 11671 25594 11677 25596
rect 11431 25542 11433 25594
rect 11613 25542 11615 25594
rect 11369 25540 11375 25542
rect 11431 25540 11455 25542
rect 11511 25540 11535 25542
rect 11591 25540 11615 25542
rect 11671 25540 11677 25542
rect 11369 25531 11677 25540
rect 11808 25362 11836 26250
rect 12268 26246 12296 26930
rect 12532 26920 12584 26926
rect 12532 26862 12584 26868
rect 12072 26240 12124 26246
rect 12072 26182 12124 26188
rect 12256 26240 12308 26246
rect 12256 26182 12308 26188
rect 12084 25906 12112 26182
rect 12544 26042 12572 26862
rect 12532 26036 12584 26042
rect 12532 25978 12584 25984
rect 12072 25900 12124 25906
rect 12072 25842 12124 25848
rect 11244 25356 11296 25362
rect 11244 25298 11296 25304
rect 11796 25356 11848 25362
rect 11796 25298 11848 25304
rect 11256 24138 11284 25298
rect 12084 24818 12112 25842
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 11796 24744 11848 24750
rect 11796 24686 11848 24692
rect 12348 24744 12400 24750
rect 12348 24686 12400 24692
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 11369 24508 11677 24517
rect 11369 24506 11375 24508
rect 11431 24506 11455 24508
rect 11511 24506 11535 24508
rect 11591 24506 11615 24508
rect 11671 24506 11677 24508
rect 11431 24454 11433 24506
rect 11613 24454 11615 24506
rect 11369 24452 11375 24454
rect 11431 24452 11455 24454
rect 11511 24452 11535 24454
rect 11591 24452 11615 24454
rect 11671 24452 11677 24454
rect 11369 24443 11677 24452
rect 11716 24206 11744 24550
rect 11808 24410 11836 24686
rect 11796 24404 11848 24410
rect 11796 24346 11848 24352
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 11244 24132 11296 24138
rect 11244 24074 11296 24080
rect 12164 24064 12216 24070
rect 12164 24006 12216 24012
rect 11369 23420 11677 23429
rect 11369 23418 11375 23420
rect 11431 23418 11455 23420
rect 11511 23418 11535 23420
rect 11591 23418 11615 23420
rect 11671 23418 11677 23420
rect 11431 23366 11433 23418
rect 11613 23366 11615 23418
rect 11369 23364 11375 23366
rect 11431 23364 11455 23366
rect 11511 23364 11535 23366
rect 11591 23364 11615 23366
rect 11671 23364 11677 23366
rect 11369 23355 11677 23364
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 10416 22160 10468 22166
rect 10416 22102 10468 22108
rect 10428 22030 10456 22102
rect 10416 22024 10468 22030
rect 10416 21966 10468 21972
rect 10140 21684 10192 21690
rect 10140 21626 10192 21632
rect 10140 21548 10192 21554
rect 10140 21490 10192 21496
rect 10152 20942 10180 21490
rect 10428 21486 10456 21966
rect 10416 21480 10468 21486
rect 10416 21422 10468 21428
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 10152 20602 10180 20878
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10520 20058 10548 23122
rect 11060 22704 11112 22710
rect 11060 22646 11112 22652
rect 10968 22432 11020 22438
rect 10968 22374 11020 22380
rect 10876 21616 10928 21622
rect 10876 21558 10928 21564
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10704 20466 10732 21490
rect 10888 20466 10916 21558
rect 10980 21554 11008 22374
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 11072 20602 11100 22646
rect 11152 22636 11204 22642
rect 11152 22578 11204 22584
rect 11164 21690 11192 22578
rect 11244 22568 11296 22574
rect 11244 22510 11296 22516
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10508 20052 10560 20058
rect 10508 19994 10560 20000
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10612 19242 10640 19790
rect 10600 19236 10652 19242
rect 10600 19178 10652 19184
rect 10612 18698 10640 19178
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10612 17746 10640 18634
rect 11256 17882 11284 22510
rect 11980 22432 12032 22438
rect 11980 22374 12032 22380
rect 11369 22332 11677 22341
rect 11369 22330 11375 22332
rect 11431 22330 11455 22332
rect 11511 22330 11535 22332
rect 11591 22330 11615 22332
rect 11671 22330 11677 22332
rect 11431 22278 11433 22330
rect 11613 22278 11615 22330
rect 11369 22276 11375 22278
rect 11431 22276 11455 22278
rect 11511 22276 11535 22278
rect 11591 22276 11615 22278
rect 11671 22276 11677 22278
rect 11369 22267 11677 22276
rect 11369 21244 11677 21253
rect 11369 21242 11375 21244
rect 11431 21242 11455 21244
rect 11511 21242 11535 21244
rect 11591 21242 11615 21244
rect 11671 21242 11677 21244
rect 11431 21190 11433 21242
rect 11613 21190 11615 21242
rect 11369 21188 11375 21190
rect 11431 21188 11455 21190
rect 11511 21188 11535 21190
rect 11591 21188 11615 21190
rect 11671 21188 11677 21190
rect 11369 21179 11677 21188
rect 11992 20466 12020 22374
rect 12176 20466 12204 24006
rect 12256 22976 12308 22982
rect 12256 22918 12308 22924
rect 12268 22642 12296 22918
rect 12256 22636 12308 22642
rect 12256 22578 12308 22584
rect 12360 22522 12388 24686
rect 12440 24676 12492 24682
rect 12440 24618 12492 24624
rect 12452 24206 12480 24618
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 12532 24200 12584 24206
rect 12532 24142 12584 24148
rect 12544 23322 12572 24142
rect 12636 23338 12664 27338
rect 12808 26920 12860 26926
rect 12808 26862 12860 26868
rect 12820 26586 12848 26862
rect 13176 26784 13228 26790
rect 13176 26726 13228 26732
rect 12808 26580 12860 26586
rect 12808 26522 12860 26528
rect 13188 26382 13216 26726
rect 13176 26376 13228 26382
rect 13176 26318 13228 26324
rect 13188 25294 13216 26318
rect 13176 25288 13228 25294
rect 13176 25230 13228 25236
rect 12716 24608 12768 24614
rect 12716 24550 12768 24556
rect 12728 24410 12756 24550
rect 12716 24404 12768 24410
rect 12716 24346 12768 24352
rect 12532 23316 12584 23322
rect 12636 23310 12756 23338
rect 12532 23258 12584 23264
rect 12624 23180 12676 23186
rect 12624 23122 12676 23128
rect 12440 22704 12492 22710
rect 12440 22646 12492 22652
rect 12268 22494 12388 22522
rect 12268 22030 12296 22494
rect 12452 22098 12480 22646
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12636 22030 12664 23122
rect 12256 22024 12308 22030
rect 12256 21966 12308 21972
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12268 21350 12296 21966
rect 12532 21956 12584 21962
rect 12532 21898 12584 21904
rect 12348 21480 12400 21486
rect 12348 21422 12400 21428
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 12164 20460 12216 20466
rect 12164 20402 12216 20408
rect 11369 20156 11677 20165
rect 11369 20154 11375 20156
rect 11431 20154 11455 20156
rect 11511 20154 11535 20156
rect 11591 20154 11615 20156
rect 11671 20154 11677 20156
rect 11431 20102 11433 20154
rect 11613 20102 11615 20154
rect 11369 20100 11375 20102
rect 11431 20100 11455 20102
rect 11511 20100 11535 20102
rect 11591 20100 11615 20102
rect 11671 20100 11677 20102
rect 11369 20091 11677 20100
rect 12164 20052 12216 20058
rect 12164 19994 12216 20000
rect 11612 19780 11664 19786
rect 11612 19722 11664 19728
rect 11624 19514 11652 19722
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 12176 19446 12204 19994
rect 12360 19922 12388 21422
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12164 19440 12216 19446
rect 12164 19382 12216 19388
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 11369 19068 11677 19077
rect 11369 19066 11375 19068
rect 11431 19066 11455 19068
rect 11511 19066 11535 19068
rect 11591 19066 11615 19068
rect 11671 19066 11677 19068
rect 11431 19014 11433 19066
rect 11613 19014 11615 19066
rect 11369 19012 11375 19014
rect 11431 19012 11455 19014
rect 11511 19012 11535 19014
rect 11591 19012 11615 19014
rect 11671 19012 11677 19014
rect 11369 19003 11677 19012
rect 11369 17980 11677 17989
rect 11369 17978 11375 17980
rect 11431 17978 11455 17980
rect 11511 17978 11535 17980
rect 11591 17978 11615 17980
rect 11671 17978 11677 17980
rect 11431 17926 11433 17978
rect 11613 17926 11615 17978
rect 11369 17924 11375 17926
rect 11431 17924 11455 17926
rect 11511 17924 11535 17926
rect 11591 17924 11615 17926
rect 11671 17924 11677 17926
rect 11369 17915 11677 17924
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 10600 17740 10652 17746
rect 10600 17682 10652 17688
rect 9956 17536 10008 17542
rect 9956 17478 10008 17484
rect 10612 17202 10640 17682
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 9692 15502 9720 16934
rect 10612 16794 10640 17138
rect 11369 16892 11677 16901
rect 11369 16890 11375 16892
rect 11431 16890 11455 16892
rect 11511 16890 11535 16892
rect 11591 16890 11615 16892
rect 11671 16890 11677 16892
rect 11431 16838 11433 16890
rect 11613 16838 11615 16890
rect 11369 16836 11375 16838
rect 11431 16836 11455 16838
rect 11511 16836 11535 16838
rect 11591 16836 11615 16838
rect 11671 16836 11677 16838
rect 11369 16827 11677 16836
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11716 16046 11744 16594
rect 11808 16250 11836 17138
rect 12084 16454 12112 19314
rect 12544 18970 12572 21898
rect 12728 21434 12756 23310
rect 13188 23186 13216 25230
rect 13176 23180 13228 23186
rect 13176 23122 13228 23128
rect 12808 23112 12860 23118
rect 12808 23054 12860 23060
rect 12820 22030 12848 23054
rect 13360 22568 13412 22574
rect 13360 22510 13412 22516
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 13268 22024 13320 22030
rect 13268 21966 13320 21972
rect 12820 21690 12848 21966
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 12728 21406 12848 21434
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12728 19922 12756 21286
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12820 18290 12848 21406
rect 13004 21146 13032 21490
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 13176 20324 13228 20330
rect 13176 20266 13228 20272
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 13004 19378 13032 19790
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 13188 18698 13216 20266
rect 13280 19514 13308 21966
rect 13372 21146 13400 22510
rect 13544 21956 13596 21962
rect 13544 21898 13596 21904
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 13372 20806 13400 21082
rect 13464 21010 13492 21626
rect 13556 21622 13584 21898
rect 13544 21616 13596 21622
rect 13544 21558 13596 21564
rect 13452 21004 13504 21010
rect 13452 20946 13504 20952
rect 13360 20800 13412 20806
rect 13360 20742 13412 20748
rect 13556 20466 13584 21558
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13268 19372 13320 19378
rect 13372 19360 13400 19654
rect 13320 19332 13400 19360
rect 13268 19314 13320 19320
rect 13176 18692 13228 18698
rect 13176 18634 13228 18640
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 13096 18086 13124 18226
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 12348 17604 12400 17610
rect 12348 17546 12400 17552
rect 12360 16794 12388 17546
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 13004 17066 13032 17478
rect 13096 17354 13124 18022
rect 13188 17746 13216 18634
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 13096 17326 13216 17354
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 12992 17060 13044 17066
rect 12992 17002 13044 17008
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 13004 16590 13032 17002
rect 13096 16998 13124 17138
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 13096 16658 13124 16934
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 11060 16040 11112 16046
rect 10980 15988 11060 15994
rect 10980 15982 11112 15988
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 10980 15966 11100 15982
rect 10980 15910 11008 15966
rect 11992 15910 12020 16050
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 10980 15570 11008 15846
rect 11369 15804 11677 15813
rect 11369 15802 11375 15804
rect 11431 15802 11455 15804
rect 11511 15802 11535 15804
rect 11591 15802 11615 15804
rect 11671 15802 11677 15804
rect 11431 15750 11433 15802
rect 11613 15750 11615 15802
rect 11369 15748 11375 15750
rect 11431 15748 11455 15750
rect 11511 15748 11535 15750
rect 11591 15748 11615 15750
rect 11671 15748 11677 15750
rect 11369 15739 11677 15748
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 6552 15428 6604 15434
rect 6552 15370 6604 15376
rect 9956 15428 10008 15434
rect 9956 15370 10008 15376
rect 7896 15260 8204 15269
rect 7896 15258 7902 15260
rect 7958 15258 7982 15260
rect 8038 15258 8062 15260
rect 8118 15258 8142 15260
rect 8198 15258 8204 15260
rect 7958 15206 7960 15258
rect 8140 15206 8142 15258
rect 7896 15204 7902 15206
rect 7958 15204 7982 15206
rect 8038 15204 8062 15206
rect 8118 15204 8142 15206
rect 8198 15204 8204 15206
rect 7896 15195 8204 15204
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 6564 14482 6592 14962
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6564 13326 6592 14418
rect 6656 14346 6684 14758
rect 7484 14346 7512 14962
rect 9968 14822 9996 15370
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 6644 14340 6696 14346
rect 6644 14282 6696 14288
rect 7472 14340 7524 14346
rect 7472 14282 7524 14288
rect 7484 13938 7512 14282
rect 7576 13938 7604 14758
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9600 14414 9628 14554
rect 9968 14414 9996 14758
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 8208 14272 8260 14278
rect 8260 14232 8340 14260
rect 8208 14214 8260 14220
rect 7896 14172 8204 14181
rect 7896 14170 7902 14172
rect 7958 14170 7982 14172
rect 8038 14170 8062 14172
rect 8118 14170 8142 14172
rect 8198 14170 8204 14172
rect 7958 14118 7960 14170
rect 8140 14118 8142 14170
rect 7896 14116 7902 14118
rect 7958 14116 7982 14118
rect 8038 14116 8062 14118
rect 8118 14116 8142 14118
rect 8198 14116 8204 14118
rect 7896 14107 8204 14116
rect 8208 14000 8260 14006
rect 8312 13988 8340 14232
rect 9600 14074 9628 14350
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 8260 13960 8340 13988
rect 9864 14000 9916 14006
rect 8208 13942 8260 13948
rect 9864 13942 9916 13948
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 9876 13462 9904 13942
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6564 12850 6592 13262
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 7196 13252 7248 13258
rect 7196 13194 7248 13200
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 6656 12986 6684 13194
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 7024 12986 7052 13126
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 7208 12782 7236 13194
rect 7896 13084 8204 13093
rect 7896 13082 7902 13084
rect 7958 13082 7982 13084
rect 8038 13082 8062 13084
rect 8118 13082 8142 13084
rect 8198 13082 8204 13084
rect 7958 13030 7960 13082
rect 8140 13030 8142 13082
rect 7896 13028 7902 13030
rect 7958 13028 7982 13030
rect 8038 13028 8062 13030
rect 8118 13028 8142 13030
rect 8198 13028 8204 13030
rect 7896 13019 8204 13028
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 6552 12164 6604 12170
rect 6552 12106 6604 12112
rect 6564 11898 6592 12106
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7024 11898 7052 12038
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6380 11354 6408 11698
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 7024 11286 7052 11834
rect 7208 11694 7236 12718
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8496 12238 8524 12582
rect 9324 12306 9352 13194
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9784 12442 9812 12786
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 7896 11996 8204 12005
rect 7896 11994 7902 11996
rect 7958 11994 7982 11996
rect 8038 11994 8062 11996
rect 8118 11994 8142 11996
rect 8198 11994 8204 11996
rect 7958 11942 7960 11994
rect 8140 11942 8142 11994
rect 7896 11940 7902 11942
rect 7958 11940 7982 11942
rect 8038 11940 8062 11942
rect 8118 11940 8142 11942
rect 8198 11940 8204 11942
rect 7896 11931 8204 11940
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7116 10674 7144 10950
rect 7668 10742 7696 10950
rect 7896 10908 8204 10917
rect 7896 10906 7902 10908
rect 7958 10906 7982 10908
rect 8038 10906 8062 10908
rect 8118 10906 8142 10908
rect 8198 10906 8204 10908
rect 7958 10854 7960 10906
rect 8140 10854 8142 10906
rect 7896 10852 7902 10854
rect 7958 10852 7982 10854
rect 8038 10852 8062 10854
rect 8118 10852 8142 10854
rect 8198 10852 8204 10854
rect 7896 10843 8204 10852
rect 7656 10736 7708 10742
rect 7656 10678 7708 10684
rect 8116 10736 8168 10742
rect 8116 10678 8168 10684
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 8128 10130 8156 10678
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 7896 9820 8204 9829
rect 7896 9818 7902 9820
rect 7958 9818 7982 9820
rect 8038 9818 8062 9820
rect 8118 9818 8142 9820
rect 8198 9818 8204 9820
rect 7958 9766 7960 9818
rect 8140 9766 8142 9818
rect 7896 9764 7902 9766
rect 7958 9764 7982 9766
rect 8038 9764 8062 9766
rect 8118 9764 8142 9766
rect 8198 9764 8204 9766
rect 7896 9755 8204 9764
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 6932 7970 6960 8910
rect 7024 8634 7052 8978
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 6932 7942 7052 7970
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 5000 5778 5028 7346
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5828 6798 5856 7142
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5828 6254 5856 6734
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 6104 5710 6132 6598
rect 6472 6458 6500 6598
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6564 6390 6592 6598
rect 6552 6384 6604 6390
rect 6552 6326 6604 6332
rect 6564 5914 6592 6326
rect 6748 6186 6776 6802
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 3424 5296 3476 5302
rect 3424 5238 3476 5244
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 4172 4690 4200 5578
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4356 5234 4384 5510
rect 6564 5234 6592 5850
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6840 5166 6868 6258
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 4423 4924 4731 4933
rect 4423 4922 4429 4924
rect 4485 4922 4509 4924
rect 4565 4922 4589 4924
rect 4645 4922 4669 4924
rect 4725 4922 4731 4924
rect 4485 4870 4487 4922
rect 4667 4870 4669 4922
rect 4423 4868 4429 4870
rect 4485 4868 4509 4870
rect 4565 4868 4589 4870
rect 4645 4868 4669 4870
rect 4725 4868 4731 4870
rect 4423 4859 4731 4868
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3344 3942 3372 4082
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 4172 3602 4200 4626
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4356 4214 4384 4422
rect 4344 4208 4396 4214
rect 4344 4150 4396 4156
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 4423 3836 4731 3845
rect 4423 3834 4429 3836
rect 4485 3834 4509 3836
rect 4565 3834 4589 3836
rect 4645 3834 4669 3836
rect 4725 3834 4731 3836
rect 4485 3782 4487 3834
rect 4667 3782 4669 3834
rect 4423 3780 4429 3782
rect 4485 3780 4509 3782
rect 4565 3780 4589 3782
rect 4645 3780 4669 3782
rect 4725 3780 4731 3782
rect 4423 3771 4731 3780
rect 5092 3602 5120 4150
rect 5552 3942 5580 5102
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6656 4146 6684 4490
rect 6748 4282 6776 4558
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 6656 3738 6684 4082
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6748 3670 6776 4218
rect 6840 4146 6868 4626
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 4172 3126 4200 3538
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 6196 3194 6224 3334
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 6932 2990 6960 7754
rect 7024 7546 7052 7942
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 7024 6798 7052 7210
rect 7300 7002 7328 8978
rect 7896 8732 8204 8741
rect 7896 8730 7902 8732
rect 7958 8730 7982 8732
rect 8038 8730 8062 8732
rect 8118 8730 8142 8732
rect 8198 8730 8204 8732
rect 7958 8678 7960 8730
rect 8140 8678 8142 8730
rect 7896 8676 7902 8678
rect 7958 8676 7982 8678
rect 8038 8676 8062 8678
rect 8118 8676 8142 8678
rect 8198 8676 8204 8678
rect 7896 8667 8204 8676
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7392 7546 7420 8434
rect 7760 7546 7788 8570
rect 8496 7886 8524 11494
rect 9232 11218 9260 12174
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9048 7886 9076 11154
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9140 10742 9168 11086
rect 9128 10736 9180 10742
rect 9128 10678 9180 10684
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 9324 8090 9352 10134
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9416 8498 9444 8910
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 7896 7644 8204 7653
rect 7896 7642 7902 7644
rect 7958 7642 7982 7644
rect 8038 7642 8062 7644
rect 8118 7642 8142 7644
rect 8198 7642 8204 7644
rect 7958 7590 7960 7642
rect 8140 7590 8142 7642
rect 7896 7588 7902 7590
rect 7958 7588 7982 7590
rect 8038 7588 8062 7590
rect 8118 7588 8142 7590
rect 8198 7588 8204 7590
rect 7896 7579 8204 7588
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 9140 6866 9168 7686
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 7024 3602 7052 3878
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 7116 3398 7144 6258
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7668 5710 7696 6054
rect 7760 5914 7788 6666
rect 7896 6556 8204 6565
rect 7896 6554 7902 6556
rect 7958 6554 7982 6556
rect 8038 6554 8062 6556
rect 8118 6554 8142 6556
rect 8198 6554 8204 6556
rect 7958 6502 7960 6554
rect 8140 6502 8142 6554
rect 7896 6500 7902 6502
rect 7958 6500 7982 6502
rect 8038 6500 8062 6502
rect 8118 6500 8142 6502
rect 8198 6500 8204 6502
rect 7896 6491 8204 6500
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 8496 5710 8524 6054
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 7300 5370 7328 5646
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7576 5370 7604 5578
rect 7896 5468 8204 5477
rect 7896 5466 7902 5468
rect 7958 5466 7982 5468
rect 8038 5466 8062 5468
rect 8118 5466 8142 5468
rect 8198 5466 8204 5468
rect 7958 5414 7960 5466
rect 8140 5414 8142 5466
rect 7896 5412 7902 5414
rect 7958 5412 7982 5414
rect 8038 5412 8062 5414
rect 8118 5412 8142 5414
rect 8198 5412 8204 5414
rect 7896 5403 8204 5412
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 8312 5234 8340 5646
rect 8496 5302 8524 5646
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8312 4622 8340 5170
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 7288 3460 7340 3466
rect 7288 3402 7340 3408
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 7116 2922 7144 3334
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 4423 2748 4731 2757
rect 4423 2746 4429 2748
rect 4485 2746 4509 2748
rect 4565 2746 4589 2748
rect 4645 2746 4669 2748
rect 4725 2746 4731 2748
rect 4485 2694 4487 2746
rect 4667 2694 4669 2746
rect 4423 2692 4429 2694
rect 4485 2692 4509 2694
rect 4565 2692 4589 2694
rect 4645 2692 4669 2694
rect 4725 2692 4731 2694
rect 4423 2683 4731 2692
rect 7116 2446 7144 2858
rect 7300 2650 7328 3402
rect 7392 3126 7420 4422
rect 7896 4380 8204 4389
rect 7896 4378 7902 4380
rect 7958 4378 7982 4380
rect 8038 4378 8062 4380
rect 8118 4378 8142 4380
rect 8198 4378 8204 4380
rect 7958 4326 7960 4378
rect 8140 4326 8142 4378
rect 7896 4324 7902 4326
rect 7958 4324 7982 4326
rect 8038 4324 8062 4326
rect 8118 4324 8142 4326
rect 8198 4324 8204 4326
rect 7896 4315 8204 4324
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8312 3534 8340 4014
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 7896 3292 8204 3301
rect 7896 3290 7902 3292
rect 7958 3290 7982 3292
rect 8038 3290 8062 3292
rect 8118 3290 8142 3292
rect 8198 3290 8204 3292
rect 7958 3238 7960 3290
rect 8140 3238 8142 3290
rect 7896 3236 7902 3238
rect 7958 3236 7982 3238
rect 8038 3236 8062 3238
rect 8118 3236 8142 3238
rect 8198 3236 8204 3238
rect 7896 3227 8204 3236
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 8404 3058 8432 4422
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9324 3738 9352 4014
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9416 3670 9444 8434
rect 9508 7546 9536 12038
rect 9876 11830 9904 13398
rect 9968 13326 9996 14350
rect 10428 14074 10456 14962
rect 10520 14482 10548 15302
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 10888 14074 10916 14758
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 9968 12714 9996 13262
rect 10796 12918 10824 13874
rect 10980 13870 11008 15506
rect 11072 15366 11100 15574
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 9956 12708 10008 12714
rect 9956 12650 10008 12656
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 10704 11762 10732 12582
rect 10796 12374 10824 12854
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10888 12170 10916 12650
rect 10980 12306 11008 13262
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10876 12164 10928 12170
rect 10876 12106 10928 12112
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9600 8906 9628 9522
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9508 6662 9536 7278
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9508 6322 9536 6598
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9600 6254 9628 7754
rect 9692 6798 9720 11698
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9784 9586 9812 10202
rect 10244 9586 10272 11154
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 9784 8974 9812 9522
rect 10520 9178 10548 9522
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10612 9110 10640 9590
rect 10796 9450 10824 11630
rect 10888 9994 10916 12106
rect 11072 11898 11100 15302
rect 11256 15026 11284 15302
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11256 14618 11284 14962
rect 11369 14716 11677 14725
rect 11369 14714 11375 14716
rect 11431 14714 11455 14716
rect 11511 14714 11535 14716
rect 11591 14714 11615 14716
rect 11671 14714 11677 14716
rect 11431 14662 11433 14714
rect 11613 14662 11615 14714
rect 11369 14660 11375 14662
rect 11431 14660 11455 14662
rect 11511 14660 11535 14662
rect 11591 14660 11615 14662
rect 11671 14660 11677 14662
rect 11369 14651 11677 14660
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11369 13628 11677 13637
rect 11369 13626 11375 13628
rect 11431 13626 11455 13628
rect 11511 13626 11535 13628
rect 11591 13626 11615 13628
rect 11671 13626 11677 13628
rect 11431 13574 11433 13626
rect 11613 13574 11615 13626
rect 11369 13572 11375 13574
rect 11431 13572 11455 13574
rect 11511 13572 11535 13574
rect 11591 13572 11615 13574
rect 11671 13572 11677 13574
rect 11369 13563 11677 13572
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 11072 11218 11100 11834
rect 11164 11762 11192 13126
rect 11369 12540 11677 12549
rect 11369 12538 11375 12540
rect 11431 12538 11455 12540
rect 11511 12538 11535 12540
rect 11591 12538 11615 12540
rect 11671 12538 11677 12540
rect 11431 12486 11433 12538
rect 11613 12486 11615 12538
rect 11369 12484 11375 12486
rect 11431 12484 11455 12486
rect 11511 12484 11535 12486
rect 11591 12484 11615 12486
rect 11671 12484 11677 12486
rect 11369 12475 11677 12484
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11256 11150 11284 12174
rect 11369 11452 11677 11461
rect 11369 11450 11375 11452
rect 11431 11450 11455 11452
rect 11511 11450 11535 11452
rect 11591 11450 11615 11452
rect 11671 11450 11677 11452
rect 11431 11398 11433 11450
rect 11613 11398 11615 11450
rect 11369 11396 11375 11398
rect 11431 11396 11455 11398
rect 11511 11396 11535 11398
rect 11591 11396 11615 11398
rect 11671 11396 11677 11398
rect 11369 11387 11677 11396
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11369 10364 11677 10373
rect 11369 10362 11375 10364
rect 11431 10362 11455 10364
rect 11511 10362 11535 10364
rect 11591 10362 11615 10364
rect 11671 10362 11677 10364
rect 11431 10310 11433 10362
rect 11613 10310 11615 10362
rect 11369 10308 11375 10310
rect 11431 10308 11455 10310
rect 11511 10308 11535 10310
rect 11591 10308 11615 10310
rect 11671 10308 11677 10310
rect 11369 10299 11677 10308
rect 10876 9988 10928 9994
rect 10876 9930 10928 9936
rect 10888 9738 10916 9930
rect 10888 9710 11008 9738
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 10796 8498 10824 9386
rect 10888 8634 10916 9522
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10980 7970 11008 9710
rect 11369 9276 11677 9285
rect 11369 9274 11375 9276
rect 11431 9274 11455 9276
rect 11511 9274 11535 9276
rect 11591 9274 11615 9276
rect 11671 9274 11677 9276
rect 11431 9222 11433 9274
rect 11613 9222 11615 9274
rect 11369 9220 11375 9222
rect 11431 9220 11455 9222
rect 11511 9220 11535 9222
rect 11591 9220 11615 9222
rect 11671 9220 11677 9222
rect 11369 9211 11677 9220
rect 11716 9042 11744 13262
rect 11992 12186 12020 15846
rect 12084 13138 12112 16390
rect 12268 16182 12296 16526
rect 12900 16516 12952 16522
rect 12900 16458 12952 16464
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12452 15570 12480 15914
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12636 15434 12664 16050
rect 12912 15978 12940 16458
rect 13096 16250 13124 16594
rect 13188 16590 13216 17326
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 13188 16114 13216 16526
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 12900 15972 12952 15978
rect 12900 15914 12952 15920
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12360 14414 12388 14962
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12636 14346 12664 15370
rect 12820 14618 12848 15370
rect 12912 14958 12940 15914
rect 13280 15434 13308 19314
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13464 16250 13492 18770
rect 13556 18766 13584 19246
rect 13648 19242 13676 20334
rect 13636 19236 13688 19242
rect 13636 19178 13688 19184
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13556 18154 13584 18702
rect 13648 18630 13676 19178
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 13740 18290 13768 27338
rect 16948 27328 17000 27334
rect 16948 27270 17000 27276
rect 14842 27228 15150 27237
rect 14842 27226 14848 27228
rect 14904 27226 14928 27228
rect 14984 27226 15008 27228
rect 15064 27226 15088 27228
rect 15144 27226 15150 27228
rect 14904 27174 14906 27226
rect 15086 27174 15088 27226
rect 14842 27172 14848 27174
rect 14904 27172 14928 27174
rect 14984 27172 15008 27174
rect 15064 27172 15088 27174
rect 15144 27172 15150 27174
rect 14842 27163 15150 27172
rect 16960 27062 16988 27270
rect 16948 27056 17000 27062
rect 16948 26998 17000 27004
rect 15292 26988 15344 26994
rect 15292 26930 15344 26936
rect 15304 26450 15332 26930
rect 16764 26852 16816 26858
rect 16764 26794 16816 26800
rect 15292 26444 15344 26450
rect 15292 26386 15344 26392
rect 14372 26376 14424 26382
rect 14372 26318 14424 26324
rect 14556 26376 14608 26382
rect 14556 26318 14608 26324
rect 16304 26376 16356 26382
rect 16304 26318 16356 26324
rect 14096 25832 14148 25838
rect 14096 25774 14148 25780
rect 14108 25498 14136 25774
rect 14096 25492 14148 25498
rect 14096 25434 14148 25440
rect 14384 25294 14412 26318
rect 14568 25362 14596 26318
rect 14842 26140 15150 26149
rect 14842 26138 14848 26140
rect 14904 26138 14928 26140
rect 14984 26138 15008 26140
rect 15064 26138 15088 26140
rect 15144 26138 15150 26140
rect 14904 26086 14906 26138
rect 15086 26086 15088 26138
rect 14842 26084 14848 26086
rect 14904 26084 14928 26086
rect 14984 26084 15008 26086
rect 15064 26084 15088 26086
rect 15144 26084 15150 26086
rect 14842 26075 15150 26084
rect 15384 25968 15436 25974
rect 15384 25910 15436 25916
rect 15396 25362 15424 25910
rect 15660 25696 15712 25702
rect 15660 25638 15712 25644
rect 14556 25356 14608 25362
rect 14556 25298 14608 25304
rect 15384 25356 15436 25362
rect 15384 25298 15436 25304
rect 14372 25288 14424 25294
rect 14372 25230 14424 25236
rect 14280 24880 14332 24886
rect 14280 24822 14332 24828
rect 14292 24070 14320 24822
rect 14568 24562 14596 25298
rect 14842 25052 15150 25061
rect 14842 25050 14848 25052
rect 14904 25050 14928 25052
rect 14984 25050 15008 25052
rect 15064 25050 15088 25052
rect 15144 25050 15150 25052
rect 14904 24998 14906 25050
rect 15086 24998 15088 25050
rect 14842 24996 14848 24998
rect 14904 24996 14928 24998
rect 14984 24996 15008 24998
rect 15064 24996 15088 24998
rect 15144 24996 15150 24998
rect 14842 24987 15150 24996
rect 15672 24818 15700 25638
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 14740 24744 14792 24750
rect 14740 24686 14792 24692
rect 15016 24744 15068 24750
rect 15016 24686 15068 24692
rect 14476 24534 14596 24562
rect 14372 24132 14424 24138
rect 14372 24074 14424 24080
rect 14280 24064 14332 24070
rect 14280 24006 14332 24012
rect 14292 23730 14320 24006
rect 14280 23724 14332 23730
rect 14280 23666 14332 23672
rect 14384 23322 14412 24074
rect 14372 23316 14424 23322
rect 14372 23258 14424 23264
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 13832 20534 13860 21286
rect 13820 20528 13872 20534
rect 13820 20470 13872 20476
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13544 18148 13596 18154
rect 13544 18090 13596 18096
rect 13740 17610 13768 18226
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13832 17678 13860 18158
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13728 17604 13780 17610
rect 13728 17546 13780 17552
rect 13740 17134 13768 17546
rect 13832 17202 13860 17614
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13740 16590 13768 17070
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 14108 16522 14136 22918
rect 14188 22568 14240 22574
rect 14188 22510 14240 22516
rect 14200 21554 14228 22510
rect 14476 22030 14504 24534
rect 14556 23656 14608 23662
rect 14556 23598 14608 23604
rect 14568 22982 14596 23598
rect 14752 23186 14780 24686
rect 15028 24410 15056 24686
rect 15016 24404 15068 24410
rect 15016 24346 15068 24352
rect 14842 23964 15150 23973
rect 14842 23962 14848 23964
rect 14904 23962 14928 23964
rect 14984 23962 15008 23964
rect 15064 23962 15088 23964
rect 15144 23962 15150 23964
rect 14904 23910 14906 23962
rect 15086 23910 15088 23962
rect 14842 23908 14848 23910
rect 14904 23908 14928 23910
rect 14984 23908 15008 23910
rect 15064 23908 15088 23910
rect 15144 23908 15150 23910
rect 14842 23899 15150 23908
rect 14740 23180 14792 23186
rect 14740 23122 14792 23128
rect 15672 23118 15700 24754
rect 14648 23112 14700 23118
rect 14648 23054 14700 23060
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14476 20942 14504 21966
rect 14660 21010 14688 23054
rect 16212 22976 16264 22982
rect 16212 22918 16264 22924
rect 14842 22876 15150 22885
rect 14842 22874 14848 22876
rect 14904 22874 14928 22876
rect 14984 22874 15008 22876
rect 15064 22874 15088 22876
rect 15144 22874 15150 22876
rect 14904 22822 14906 22874
rect 15086 22822 15088 22874
rect 14842 22820 14848 22822
rect 14904 22820 14928 22822
rect 14984 22820 15008 22822
rect 15064 22820 15088 22822
rect 15144 22820 15150 22822
rect 14842 22811 15150 22820
rect 15292 22704 15344 22710
rect 15292 22646 15344 22652
rect 15304 22098 15332 22646
rect 16224 22642 16252 22918
rect 16212 22636 16264 22642
rect 16212 22578 16264 22584
rect 15936 22568 15988 22574
rect 15936 22510 15988 22516
rect 15292 22092 15344 22098
rect 15292 22034 15344 22040
rect 14842 21788 15150 21797
rect 14842 21786 14848 21788
rect 14904 21786 14928 21788
rect 14984 21786 15008 21788
rect 15064 21786 15088 21788
rect 15144 21786 15150 21788
rect 14904 21734 14906 21786
rect 15086 21734 15088 21786
rect 14842 21732 14848 21734
rect 14904 21732 14928 21734
rect 14984 21732 15008 21734
rect 15064 21732 15088 21734
rect 15144 21732 15150 21734
rect 14842 21723 15150 21732
rect 15948 21690 15976 22510
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 14740 21480 14792 21486
rect 14740 21422 14792 21428
rect 14648 21004 14700 21010
rect 14648 20946 14700 20952
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14556 20868 14608 20874
rect 14556 20810 14608 20816
rect 14280 20800 14332 20806
rect 14280 20742 14332 20748
rect 14292 20534 14320 20742
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 14568 19922 14596 20810
rect 14556 19916 14608 19922
rect 14476 19876 14556 19904
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14200 16658 14228 19314
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14292 18222 14320 18634
rect 14280 18216 14332 18222
rect 14280 18158 14332 18164
rect 14292 17066 14320 18158
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14384 17542 14412 18022
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14384 17338 14412 17478
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 14280 17060 14332 17066
rect 14280 17002 14332 17008
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 13820 16516 13872 16522
rect 13820 16458 13872 16464
rect 14096 16516 14148 16522
rect 14096 16458 14148 16464
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 12992 15428 13044 15434
rect 12992 15370 13044 15376
rect 13268 15428 13320 15434
rect 13268 15370 13320 15376
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12176 13326 12204 13874
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12084 13110 12204 13138
rect 11900 12158 12020 12186
rect 11900 12102 11928 12158
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 12084 11898 12112 12038
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11532 8838 11560 8978
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10888 7942 11008 7970
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9968 5914 9996 6258
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 10244 5642 10272 6734
rect 10520 5778 10548 7278
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10612 6798 10640 7142
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10704 5914 10732 7890
rect 10888 7886 10916 7942
rect 11072 7886 11100 8774
rect 11532 8566 11560 8774
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11369 8188 11677 8197
rect 11369 8186 11375 8188
rect 11431 8186 11455 8188
rect 11511 8186 11535 8188
rect 11591 8186 11615 8188
rect 11671 8186 11677 8188
rect 11431 8134 11433 8186
rect 11613 8134 11615 8186
rect 11369 8132 11375 8134
rect 11431 8132 11455 8134
rect 11511 8132 11535 8134
rect 11591 8132 11615 8134
rect 11671 8132 11677 8134
rect 11369 8123 11677 8132
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10888 6866 10916 7822
rect 11716 7342 11744 8978
rect 11808 8498 11836 11494
rect 11992 11354 12020 11630
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 12176 11014 12204 13110
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12268 11830 12296 12038
rect 12256 11824 12308 11830
rect 12256 11766 12308 11772
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12176 9926 12204 10950
rect 12636 10130 12664 13806
rect 12820 13258 12848 14554
rect 12912 14482 12940 14894
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 13004 13326 13032 15370
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13464 15026 13492 15302
rect 13740 15026 13768 16050
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13464 14822 13492 14962
rect 13740 14822 13768 14962
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13464 14618 13492 14758
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13464 14278 13492 14554
rect 13832 14346 13860 16458
rect 14108 15638 14136 16458
rect 14096 15632 14148 15638
rect 14096 15574 14148 15580
rect 14200 14482 14228 16594
rect 14292 14890 14320 17002
rect 14476 15910 14504 19876
rect 14556 19858 14608 19864
rect 14660 19310 14688 20946
rect 14752 20806 14780 21422
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14752 20602 14780 20742
rect 14842 20700 15150 20709
rect 14842 20698 14848 20700
rect 14904 20698 14928 20700
rect 14984 20698 15008 20700
rect 15064 20698 15088 20700
rect 15144 20698 15150 20700
rect 14904 20646 14906 20698
rect 15086 20646 15088 20698
rect 14842 20644 14848 20646
rect 14904 20644 14928 20646
rect 14984 20644 15008 20646
rect 15064 20644 15088 20646
rect 15144 20644 15150 20646
rect 14842 20635 15150 20644
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14842 19612 15150 19621
rect 14842 19610 14848 19612
rect 14904 19610 14928 19612
rect 14984 19610 15008 19612
rect 15064 19610 15088 19612
rect 15144 19610 15150 19612
rect 14904 19558 14906 19610
rect 15086 19558 15088 19610
rect 14842 19556 14848 19558
rect 14904 19556 14928 19558
rect 14984 19556 15008 19558
rect 15064 19556 15088 19558
rect 15144 19556 15150 19558
rect 14842 19547 15150 19556
rect 14648 19304 14700 19310
rect 14648 19246 14700 19252
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14752 18426 14780 18702
rect 14842 18524 15150 18533
rect 14842 18522 14848 18524
rect 14904 18522 14928 18524
rect 14984 18522 15008 18524
rect 15064 18522 15088 18524
rect 15144 18522 15150 18524
rect 14904 18470 14906 18522
rect 15086 18470 15088 18522
rect 14842 18468 14848 18470
rect 14904 18468 14928 18470
rect 14984 18468 15008 18470
rect 15064 18468 15088 18470
rect 15144 18468 15150 18470
rect 14842 18459 15150 18468
rect 14740 18420 14792 18426
rect 14740 18362 14792 18368
rect 14648 18284 14700 18290
rect 14648 18226 14700 18232
rect 14660 17610 14688 18226
rect 15212 17610 15240 19246
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15304 18086 15332 18702
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 14648 17604 14700 17610
rect 14648 17546 14700 17552
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 14660 17270 14688 17546
rect 14842 17436 15150 17445
rect 14842 17434 14848 17436
rect 14904 17434 14928 17436
rect 14984 17434 15008 17436
rect 15064 17434 15088 17436
rect 15144 17434 15150 17436
rect 14904 17382 14906 17434
rect 15086 17382 15088 17434
rect 14842 17380 14848 17382
rect 14904 17380 14928 17382
rect 14984 17380 15008 17382
rect 15064 17380 15088 17382
rect 15144 17380 15150 17382
rect 14842 17371 15150 17380
rect 14648 17264 14700 17270
rect 14648 17206 14700 17212
rect 15212 17202 15240 17546
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 14740 17128 14792 17134
rect 14740 17070 14792 17076
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14280 14884 14332 14890
rect 14280 14826 14332 14832
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 14292 14074 14320 14826
rect 14568 14414 14596 16934
rect 14648 16652 14700 16658
rect 14648 16594 14700 16600
rect 14556 14408 14608 14414
rect 14556 14350 14608 14356
rect 14372 14340 14424 14346
rect 14372 14282 14424 14288
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 13372 12782 13400 13670
rect 13464 12986 13492 13942
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13464 12238 13492 12922
rect 14200 12442 14228 13874
rect 14384 13326 14412 14282
rect 14660 13462 14688 16594
rect 14752 16590 14780 17070
rect 15028 17066 15056 17138
rect 15016 17060 15068 17066
rect 15016 17002 15068 17008
rect 15212 16998 15240 17138
rect 15304 17134 15332 18022
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15212 16590 15240 16934
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 14842 16348 15150 16357
rect 14842 16346 14848 16348
rect 14904 16346 14928 16348
rect 14984 16346 15008 16348
rect 15064 16346 15088 16348
rect 15144 16346 15150 16348
rect 14904 16294 14906 16346
rect 15086 16294 15088 16346
rect 14842 16292 14848 16294
rect 14904 16292 14928 16294
rect 14984 16292 15008 16294
rect 15064 16292 15088 16294
rect 15144 16292 15150 16294
rect 14842 16283 15150 16292
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 14752 15366 14780 16050
rect 15764 16046 15792 16934
rect 15948 16182 15976 21082
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 16040 19378 16068 19790
rect 16316 19514 16344 26318
rect 16776 26314 16804 26794
rect 16764 26308 16816 26314
rect 16764 26250 16816 26256
rect 16776 21078 16804 26250
rect 16856 24744 16908 24750
rect 16856 24686 16908 24692
rect 16868 24206 16896 24686
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 16868 22030 16896 24142
rect 16960 22778 16988 26998
rect 17696 26586 17724 27474
rect 20640 27470 20668 29294
rect 24122 29200 24178 30000
rect 27802 29322 27858 30000
rect 27724 29294 27858 29322
rect 24136 27470 24164 29200
rect 27526 27840 27582 27849
rect 25261 27772 25569 27781
rect 27526 27775 27582 27784
rect 25261 27770 25267 27772
rect 25323 27770 25347 27772
rect 25403 27770 25427 27772
rect 25483 27770 25507 27772
rect 25563 27770 25569 27772
rect 25323 27718 25325 27770
rect 25505 27718 25507 27770
rect 25261 27716 25267 27718
rect 25323 27716 25347 27718
rect 25403 27716 25427 27718
rect 25483 27716 25507 27718
rect 25563 27716 25569 27718
rect 25261 27707 25569 27716
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 22284 27464 22336 27470
rect 22284 27406 22336 27412
rect 24124 27464 24176 27470
rect 24124 27406 24176 27412
rect 20904 27328 20956 27334
rect 20904 27270 20956 27276
rect 22192 27328 22244 27334
rect 22192 27270 22244 27276
rect 19800 26988 19852 26994
rect 19800 26930 19852 26936
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 18315 26684 18623 26693
rect 18315 26682 18321 26684
rect 18377 26682 18401 26684
rect 18457 26682 18481 26684
rect 18537 26682 18561 26684
rect 18617 26682 18623 26684
rect 18377 26630 18379 26682
rect 18559 26630 18561 26682
rect 18315 26628 18321 26630
rect 18377 26628 18401 26630
rect 18457 26628 18481 26630
rect 18537 26628 18561 26630
rect 18617 26628 18623 26630
rect 18315 26619 18623 26628
rect 19812 26586 19840 26930
rect 17684 26580 17736 26586
rect 17684 26522 17736 26528
rect 19800 26580 19852 26586
rect 19800 26522 19852 26528
rect 18144 26376 18196 26382
rect 18144 26318 18196 26324
rect 18156 26042 18184 26318
rect 18788 26240 18840 26246
rect 18788 26182 18840 26188
rect 19708 26240 19760 26246
rect 19708 26182 19760 26188
rect 18144 26036 18196 26042
rect 18144 25978 18196 25984
rect 18156 24818 18184 25978
rect 18800 25974 18828 26182
rect 18236 25968 18288 25974
rect 18236 25910 18288 25916
rect 18788 25968 18840 25974
rect 18788 25910 18840 25916
rect 18248 25362 18276 25910
rect 19720 25906 19748 26182
rect 19708 25900 19760 25906
rect 19708 25842 19760 25848
rect 18315 25596 18623 25605
rect 18315 25594 18321 25596
rect 18377 25594 18401 25596
rect 18457 25594 18481 25596
rect 18537 25594 18561 25596
rect 18617 25594 18623 25596
rect 18377 25542 18379 25594
rect 18559 25542 18561 25594
rect 18315 25540 18321 25542
rect 18377 25540 18401 25542
rect 18457 25540 18481 25542
rect 18537 25540 18561 25542
rect 18617 25540 18623 25542
rect 18315 25531 18623 25540
rect 18236 25356 18288 25362
rect 18236 25298 18288 25304
rect 17132 24812 17184 24818
rect 17132 24754 17184 24760
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 17144 24410 17172 24754
rect 17500 24608 17552 24614
rect 17500 24550 17552 24556
rect 17132 24404 17184 24410
rect 17132 24346 17184 24352
rect 17512 24274 17540 24550
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 16948 22772 17000 22778
rect 16948 22714 17000 22720
rect 17696 22506 17724 24210
rect 18156 24206 18184 24754
rect 18315 24508 18623 24517
rect 18315 24506 18321 24508
rect 18377 24506 18401 24508
rect 18457 24506 18481 24508
rect 18537 24506 18561 24508
rect 18617 24506 18623 24508
rect 18377 24454 18379 24506
rect 18559 24454 18561 24506
rect 18315 24452 18321 24454
rect 18377 24452 18401 24454
rect 18457 24452 18481 24454
rect 18537 24452 18561 24454
rect 18617 24452 18623 24454
rect 18315 24443 18623 24452
rect 18144 24200 18196 24206
rect 18144 24142 18196 24148
rect 19616 24200 19668 24206
rect 19616 24142 19668 24148
rect 18604 24064 18656 24070
rect 18604 24006 18656 24012
rect 18880 24064 18932 24070
rect 18880 24006 18932 24012
rect 18616 23730 18644 24006
rect 18892 23798 18920 24006
rect 18880 23792 18932 23798
rect 18880 23734 18932 23740
rect 19432 23792 19484 23798
rect 19432 23734 19484 23740
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18315 23420 18623 23429
rect 18315 23418 18321 23420
rect 18377 23418 18401 23420
rect 18457 23418 18481 23420
rect 18537 23418 18561 23420
rect 18617 23418 18623 23420
rect 18377 23366 18379 23418
rect 18559 23366 18561 23418
rect 18315 23364 18321 23366
rect 18377 23364 18401 23366
rect 18457 23364 18481 23366
rect 18537 23364 18561 23366
rect 18617 23364 18623 23366
rect 18315 23355 18623 23364
rect 19444 22778 19472 23734
rect 19628 23662 19656 24142
rect 19616 23656 19668 23662
rect 19616 23598 19668 23604
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 17776 22636 17828 22642
rect 17776 22578 17828 22584
rect 17684 22500 17736 22506
rect 17684 22442 17736 22448
rect 17500 22432 17552 22438
rect 17500 22374 17552 22380
rect 17512 22030 17540 22374
rect 16856 22024 16908 22030
rect 16856 21966 16908 21972
rect 17316 22024 17368 22030
rect 17316 21966 17368 21972
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17328 21622 17356 21966
rect 17316 21616 17368 21622
rect 17316 21558 17368 21564
rect 17500 21616 17552 21622
rect 17500 21558 17552 21564
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 17236 21146 17264 21490
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 16764 21072 16816 21078
rect 16764 21014 16816 21020
rect 17132 21072 17184 21078
rect 17132 21014 17184 21020
rect 17144 20942 17172 21014
rect 17132 20936 17184 20942
rect 17132 20878 17184 20884
rect 17144 20534 17172 20878
rect 17132 20528 17184 20534
rect 17132 20470 17184 20476
rect 16856 20392 16908 20398
rect 16856 20334 16908 20340
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16776 19922 16804 20198
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16488 19780 16540 19786
rect 16540 19740 16620 19768
rect 16488 19722 16540 19728
rect 16304 19508 16356 19514
rect 16304 19450 16356 19456
rect 16592 19446 16620 19740
rect 16868 19514 16896 20334
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 15936 16176 15988 16182
rect 15936 16118 15988 16124
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 13912 12300 13964 12306
rect 14660 12288 14688 13126
rect 14752 12918 14780 15302
rect 14842 15260 15150 15269
rect 14842 15258 14848 15260
rect 14904 15258 14928 15260
rect 14984 15258 15008 15260
rect 15064 15258 15088 15260
rect 15144 15258 15150 15260
rect 14904 15206 14906 15258
rect 15086 15206 15088 15258
rect 14842 15204 14848 15206
rect 14904 15204 14928 15206
rect 14984 15204 15008 15206
rect 15064 15204 15088 15206
rect 15144 15204 15150 15206
rect 14842 15195 15150 15204
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14844 14414 14872 14826
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14842 14172 15150 14181
rect 14842 14170 14848 14172
rect 14904 14170 14928 14172
rect 14984 14170 15008 14172
rect 15064 14170 15088 14172
rect 15144 14170 15150 14172
rect 14904 14118 14906 14170
rect 15086 14118 15088 14170
rect 14842 14116 14848 14118
rect 14904 14116 14928 14118
rect 14984 14116 15008 14118
rect 15064 14116 15088 14118
rect 15144 14116 15150 14118
rect 14842 14107 15150 14116
rect 15304 13326 15332 14894
rect 15580 14618 15608 14962
rect 16040 14958 16068 19314
rect 16580 18148 16632 18154
rect 16580 18090 16632 18096
rect 16592 16726 16620 18090
rect 16960 18086 16988 19790
rect 17040 19712 17092 19718
rect 17040 19654 17092 19660
rect 17052 19378 17080 19654
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 17512 19310 17540 21558
rect 17788 20534 17816 22578
rect 17960 22568 18012 22574
rect 17960 22510 18012 22516
rect 17868 22500 17920 22506
rect 17868 22442 17920 22448
rect 17880 21010 17908 22442
rect 17972 22234 18000 22510
rect 18315 22332 18623 22341
rect 18315 22330 18321 22332
rect 18377 22330 18401 22332
rect 18457 22330 18481 22332
rect 18537 22330 18561 22332
rect 18617 22330 18623 22332
rect 18377 22278 18379 22330
rect 18559 22278 18561 22330
rect 18315 22276 18321 22278
rect 18377 22276 18401 22278
rect 18457 22276 18481 22278
rect 18537 22276 18561 22278
rect 18617 22276 18623 22278
rect 18315 22267 18623 22276
rect 17960 22228 18012 22234
rect 17960 22170 18012 22176
rect 19628 22030 19656 23598
rect 19616 22024 19668 22030
rect 19616 21966 19668 21972
rect 19720 21554 19748 25842
rect 19812 25430 19840 26522
rect 19996 25838 20024 26930
rect 20916 26926 20944 27270
rect 21788 27228 22096 27237
rect 21788 27226 21794 27228
rect 21850 27226 21874 27228
rect 21930 27226 21954 27228
rect 22010 27226 22034 27228
rect 22090 27226 22096 27228
rect 21850 27174 21852 27226
rect 22032 27174 22034 27226
rect 21788 27172 21794 27174
rect 21850 27172 21874 27174
rect 21930 27172 21954 27174
rect 22010 27172 22034 27174
rect 22090 27172 22096 27174
rect 21788 27163 22096 27172
rect 20352 26920 20404 26926
rect 20352 26862 20404 26868
rect 20904 26920 20956 26926
rect 20904 26862 20956 26868
rect 20364 26314 20392 26862
rect 20352 26308 20404 26314
rect 20352 26250 20404 26256
rect 20720 26308 20772 26314
rect 20720 26250 20772 26256
rect 20732 26042 20760 26250
rect 20720 26036 20772 26042
rect 20720 25978 20772 25984
rect 19984 25832 20036 25838
rect 19984 25774 20036 25780
rect 19800 25424 19852 25430
rect 19852 25372 19932 25378
rect 19800 25366 19932 25372
rect 19812 25350 19932 25366
rect 19800 25288 19852 25294
rect 19800 25230 19852 25236
rect 19812 23050 19840 25230
rect 19800 23044 19852 23050
rect 19800 22986 19852 22992
rect 19812 22642 19840 22986
rect 19904 22642 19932 25350
rect 19996 25294 20024 25774
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 20916 24138 20944 26862
rect 21732 26784 21784 26790
rect 21732 26726 21784 26732
rect 21744 26450 21772 26726
rect 22204 26602 22232 27270
rect 22296 26994 22324 27406
rect 24952 27328 25004 27334
rect 24952 27270 25004 27276
rect 22836 27056 22888 27062
rect 22836 26998 22888 27004
rect 22284 26988 22336 26994
rect 22284 26930 22336 26936
rect 22112 26574 22232 26602
rect 22112 26450 22140 26574
rect 21732 26444 21784 26450
rect 21732 26386 21784 26392
rect 22100 26444 22152 26450
rect 22100 26386 22152 26392
rect 21272 26376 21324 26382
rect 21272 26318 21324 26324
rect 21284 26042 21312 26318
rect 21788 26140 22096 26149
rect 21788 26138 21794 26140
rect 21850 26138 21874 26140
rect 21930 26138 21954 26140
rect 22010 26138 22034 26140
rect 22090 26138 22096 26140
rect 21850 26086 21852 26138
rect 22032 26086 22034 26138
rect 21788 26084 21794 26086
rect 21850 26084 21874 26086
rect 21930 26084 21954 26086
rect 22010 26084 22034 26086
rect 22090 26084 22096 26086
rect 21788 26075 22096 26084
rect 22296 26042 22324 26930
rect 22376 26852 22428 26858
rect 22376 26794 22428 26800
rect 21272 26036 21324 26042
rect 21272 25978 21324 25984
rect 22284 26036 22336 26042
rect 22284 25978 22336 25984
rect 21788 25052 22096 25061
rect 21788 25050 21794 25052
rect 21850 25050 21874 25052
rect 21930 25050 21954 25052
rect 22010 25050 22034 25052
rect 22090 25050 22096 25052
rect 21850 24998 21852 25050
rect 22032 24998 22034 25050
rect 21788 24996 21794 24998
rect 21850 24996 21874 24998
rect 21930 24996 21954 24998
rect 22010 24996 22034 24998
rect 22090 24996 22096 24998
rect 21788 24987 22096 24996
rect 22388 24206 22416 26794
rect 22468 26580 22520 26586
rect 22468 26522 22520 26528
rect 22480 25906 22508 26522
rect 22468 25900 22520 25906
rect 22468 25842 22520 25848
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22756 24750 22784 25230
rect 22744 24744 22796 24750
rect 22744 24686 22796 24692
rect 22468 24268 22520 24274
rect 22468 24210 22520 24216
rect 22376 24200 22428 24206
rect 22376 24142 22428 24148
rect 20904 24132 20956 24138
rect 20904 24074 20956 24080
rect 22284 24064 22336 24070
rect 22284 24006 22336 24012
rect 21788 23964 22096 23973
rect 21788 23962 21794 23964
rect 21850 23962 21874 23964
rect 21930 23962 21954 23964
rect 22010 23962 22034 23964
rect 22090 23962 22096 23964
rect 21850 23910 21852 23962
rect 22032 23910 22034 23962
rect 21788 23908 21794 23910
rect 21850 23908 21874 23910
rect 21930 23908 21954 23910
rect 22010 23908 22034 23910
rect 22090 23908 22096 23910
rect 21788 23899 22096 23908
rect 22296 23798 22324 24006
rect 22284 23792 22336 23798
rect 22284 23734 22336 23740
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 19800 22636 19852 22642
rect 19800 22578 19852 22584
rect 19892 22636 19944 22642
rect 19892 22578 19944 22584
rect 19708 21548 19760 21554
rect 19708 21490 19760 21496
rect 17960 21412 18012 21418
rect 17960 21354 18012 21360
rect 17868 21004 17920 21010
rect 17868 20946 17920 20952
rect 17776 20528 17828 20534
rect 17776 20470 17828 20476
rect 17788 19446 17816 20470
rect 17880 20058 17908 20946
rect 17972 20942 18000 21354
rect 18315 21244 18623 21253
rect 18315 21242 18321 21244
rect 18377 21242 18401 21244
rect 18457 21242 18481 21244
rect 18537 21242 18561 21244
rect 18617 21242 18623 21244
rect 18377 21190 18379 21242
rect 18559 21190 18561 21242
rect 18315 21188 18321 21190
rect 18377 21188 18401 21190
rect 18457 21188 18481 21190
rect 18537 21188 18561 21190
rect 18617 21188 18623 21190
rect 18315 21179 18623 21188
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 18315 20156 18623 20165
rect 18315 20154 18321 20156
rect 18377 20154 18401 20156
rect 18457 20154 18481 20156
rect 18537 20154 18561 20156
rect 18617 20154 18623 20156
rect 18377 20102 18379 20154
rect 18559 20102 18561 20154
rect 18315 20100 18321 20102
rect 18377 20100 18401 20102
rect 18457 20100 18481 20102
rect 18537 20100 18561 20102
rect 18617 20100 18623 20102
rect 18315 20091 18623 20100
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 19616 19780 19668 19786
rect 19616 19722 19668 19728
rect 17776 19440 17828 19446
rect 17776 19382 17828 19388
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17420 18426 17448 18702
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17512 18358 17540 19246
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16856 17604 16908 17610
rect 16856 17546 16908 17552
rect 16868 17338 16896 17546
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 17236 17270 17264 17478
rect 17224 17264 17276 17270
rect 17224 17206 17276 17212
rect 16580 16720 16632 16726
rect 16580 16662 16632 16668
rect 16488 16176 16540 16182
rect 16488 16118 16540 16124
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 14842 13084 15150 13093
rect 14842 13082 14848 13084
rect 14904 13082 14928 13084
rect 14984 13082 15008 13084
rect 15064 13082 15088 13084
rect 15144 13082 15150 13084
rect 14904 13030 14906 13082
rect 15086 13030 15088 13082
rect 14842 13028 14848 13030
rect 14904 13028 14928 13030
rect 14984 13028 15008 13030
rect 15064 13028 15088 13030
rect 15144 13028 15150 13030
rect 14842 13019 15150 13028
rect 15396 12918 15424 14010
rect 15672 13938 15700 14214
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15488 13326 15516 13874
rect 16500 13410 16528 16118
rect 17512 16046 17540 18294
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17500 16040 17552 16046
rect 17500 15982 17552 15988
rect 16672 15972 16724 15978
rect 16672 15914 16724 15920
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 16592 15502 16620 15846
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16500 13382 16620 13410
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 15384 12912 15436 12918
rect 15384 12854 15436 12860
rect 15396 12434 15424 12854
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15212 12406 15424 12434
rect 14832 12300 14884 12306
rect 14660 12260 14832 12288
rect 13912 12242 13964 12248
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13740 11150 13768 11766
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12176 8974 12204 9862
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11369 7100 11677 7109
rect 11369 7098 11375 7100
rect 11431 7098 11455 7100
rect 11511 7098 11535 7100
rect 11591 7098 11615 7100
rect 11671 7098 11677 7100
rect 11431 7046 11433 7098
rect 11613 7046 11615 7098
rect 11369 7044 11375 7046
rect 11431 7044 11455 7046
rect 11511 7044 11535 7046
rect 11591 7044 11615 7046
rect 11671 7044 11677 7046
rect 11369 7035 11677 7044
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10888 6322 10916 6802
rect 11716 6798 11744 7278
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11808 6730 11836 8434
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 11369 6012 11677 6021
rect 11369 6010 11375 6012
rect 11431 6010 11455 6012
rect 11511 6010 11535 6012
rect 11591 6010 11615 6012
rect 11671 6010 11677 6012
rect 11431 5958 11433 6010
rect 11613 5958 11615 6010
rect 11369 5956 11375 5958
rect 11431 5956 11455 5958
rect 11511 5956 11535 5958
rect 11591 5956 11615 5958
rect 11671 5956 11677 5958
rect 11369 5947 11677 5956
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 11369 4924 11677 4933
rect 11369 4922 11375 4924
rect 11431 4922 11455 4924
rect 11511 4922 11535 4924
rect 11591 4922 11615 4924
rect 11671 4922 11677 4924
rect 11431 4870 11433 4922
rect 11613 4870 11615 4922
rect 11369 4868 11375 4870
rect 11431 4868 11455 4870
rect 11511 4868 11535 4870
rect 11591 4868 11615 4870
rect 11671 4868 11677 4870
rect 11369 4859 11677 4868
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 10600 4548 10652 4554
rect 10600 4490 10652 4496
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9692 4078 9720 4422
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9784 3942 9812 4490
rect 10612 4282 10640 4490
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9784 3058 9812 3878
rect 10704 3058 10732 4558
rect 11072 4282 11100 4626
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10888 3194 10916 4150
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 11072 3738 11100 4082
rect 11369 3836 11677 3845
rect 11369 3834 11375 3836
rect 11431 3834 11455 3836
rect 11511 3834 11535 3836
rect 11591 3834 11615 3836
rect 11671 3834 11677 3836
rect 11431 3782 11433 3834
rect 11613 3782 11615 3834
rect 11369 3780 11375 3782
rect 11431 3780 11455 3782
rect 11511 3780 11535 3782
rect 11591 3780 11615 3782
rect 11671 3780 11677 3782
rect 11369 3771 11677 3780
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11716 3466 11744 4422
rect 11900 3738 11928 8298
rect 12176 8090 12204 8774
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12360 7274 12388 10066
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12728 6746 12756 6802
rect 13096 6798 13124 11018
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13648 8090 13676 8434
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13924 7886 13952 12242
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 12636 6718 12756 6746
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12636 6662 12664 6718
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12268 6390 12296 6598
rect 12636 6458 12664 6598
rect 12728 6458 12756 6598
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 12728 5778 12756 6394
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12176 4146 12204 5646
rect 13832 4622 13860 7278
rect 13924 5914 13952 7822
rect 14016 6866 14044 12174
rect 14752 11880 14780 12260
rect 14832 12242 14884 12248
rect 15212 12238 15240 12406
rect 15672 12238 15700 12786
rect 16500 12434 16528 13262
rect 16592 12594 16620 13382
rect 16684 12850 16712 15914
rect 17420 15706 17448 15982
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17236 14006 17264 14214
rect 17224 14000 17276 14006
rect 17224 13942 17276 13948
rect 17420 13938 17448 15642
rect 17512 15434 17540 15982
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 17788 15162 17816 16050
rect 17972 15162 18000 19382
rect 19628 19310 19656 19722
rect 19616 19304 19668 19310
rect 19616 19246 19668 19252
rect 18236 19168 18288 19174
rect 18236 19110 18288 19116
rect 18248 18766 18276 19110
rect 18315 19068 18623 19077
rect 18315 19066 18321 19068
rect 18377 19066 18401 19068
rect 18457 19066 18481 19068
rect 18537 19066 18561 19068
rect 18617 19066 18623 19068
rect 18377 19014 18379 19066
rect 18559 19014 18561 19066
rect 18315 19012 18321 19014
rect 18377 19012 18401 19014
rect 18457 19012 18481 19014
rect 18537 19012 18561 19014
rect 18617 19012 18623 19014
rect 18315 19003 18623 19012
rect 19812 18766 19840 22578
rect 19904 19174 19932 22578
rect 19984 22092 20036 22098
rect 19984 22034 20036 22040
rect 19996 21146 20024 22034
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 20548 20942 20576 23666
rect 21788 22876 22096 22885
rect 21788 22874 21794 22876
rect 21850 22874 21874 22876
rect 21930 22874 21954 22876
rect 22010 22874 22034 22876
rect 22090 22874 22096 22876
rect 21850 22822 21852 22874
rect 22032 22822 22034 22874
rect 21788 22820 21794 22822
rect 21850 22820 21874 22822
rect 21930 22820 21954 22822
rect 22010 22820 22034 22822
rect 22090 22820 22096 22822
rect 21788 22811 22096 22820
rect 21788 21788 22096 21797
rect 21788 21786 21794 21788
rect 21850 21786 21874 21788
rect 21930 21786 21954 21788
rect 22010 21786 22034 21788
rect 22090 21786 22096 21788
rect 21850 21734 21852 21786
rect 22032 21734 22034 21786
rect 21788 21732 21794 21734
rect 21850 21732 21874 21734
rect 21930 21732 21954 21734
rect 22010 21732 22034 21734
rect 22090 21732 22096 21734
rect 21788 21723 22096 21732
rect 21548 21684 21600 21690
rect 21548 21626 21600 21632
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20088 20058 20116 20878
rect 20444 20868 20496 20874
rect 20444 20810 20496 20816
rect 21272 20868 21324 20874
rect 21272 20810 21324 20816
rect 20456 20602 20484 20810
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 21284 20058 21312 20810
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 20088 19446 20116 19994
rect 20904 19780 20956 19786
rect 20904 19722 20956 19728
rect 20916 19514 20944 19722
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 19892 19168 19944 19174
rect 19892 19110 19944 19116
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 19904 18766 19932 19110
rect 21192 18902 21220 19110
rect 21284 18970 21312 19314
rect 21272 18964 21324 18970
rect 21272 18906 21324 18912
rect 21180 18896 21232 18902
rect 21180 18838 21232 18844
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 19800 18760 19852 18766
rect 19800 18702 19852 18708
rect 19892 18760 19944 18766
rect 19892 18702 19944 18708
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 18880 18624 18932 18630
rect 18880 18566 18932 18572
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 18892 18358 18920 18566
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 18880 18352 18932 18358
rect 18880 18294 18932 18300
rect 18696 18216 18748 18222
rect 18696 18158 18748 18164
rect 19708 18216 19760 18222
rect 19708 18158 19760 18164
rect 18315 17980 18623 17989
rect 18315 17978 18321 17980
rect 18377 17978 18401 17980
rect 18457 17978 18481 17980
rect 18537 17978 18561 17980
rect 18617 17978 18623 17980
rect 18377 17926 18379 17978
rect 18559 17926 18561 17978
rect 18315 17924 18321 17926
rect 18377 17924 18401 17926
rect 18457 17924 18481 17926
rect 18537 17924 18561 17926
rect 18617 17924 18623 17926
rect 18315 17915 18623 17924
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 18248 16658 18276 16934
rect 18315 16892 18623 16901
rect 18315 16890 18321 16892
rect 18377 16890 18401 16892
rect 18457 16890 18481 16892
rect 18537 16890 18561 16892
rect 18617 16890 18623 16892
rect 18377 16838 18379 16890
rect 18559 16838 18561 16890
rect 18315 16836 18321 16838
rect 18377 16836 18401 16838
rect 18457 16836 18481 16838
rect 18537 16836 18561 16838
rect 18617 16836 18623 16838
rect 18315 16827 18623 16836
rect 18236 16652 18288 16658
rect 18236 16594 18288 16600
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 18248 14958 18276 16594
rect 18315 15804 18623 15813
rect 18315 15802 18321 15804
rect 18377 15802 18401 15804
rect 18457 15802 18481 15804
rect 18537 15802 18561 15804
rect 18617 15802 18623 15804
rect 18377 15750 18379 15802
rect 18559 15750 18561 15802
rect 18315 15748 18321 15750
rect 18377 15748 18401 15750
rect 18457 15748 18481 15750
rect 18537 15748 18561 15750
rect 18617 15748 18623 15750
rect 18315 15739 18623 15748
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18315 14716 18623 14725
rect 18315 14714 18321 14716
rect 18377 14714 18401 14716
rect 18457 14714 18481 14716
rect 18537 14714 18561 14716
rect 18617 14714 18623 14716
rect 18377 14662 18379 14714
rect 18559 14662 18561 14714
rect 18315 14660 18321 14662
rect 18377 14660 18401 14662
rect 18457 14660 18481 14662
rect 18537 14660 18561 14662
rect 18617 14660 18623 14662
rect 18315 14651 18623 14660
rect 18708 14550 18736 18158
rect 19720 17882 19748 18158
rect 19708 17876 19760 17882
rect 19708 17818 19760 17824
rect 19996 17678 20024 18362
rect 20272 18358 20300 18566
rect 20260 18352 20312 18358
rect 20260 18294 20312 18300
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18892 16182 18920 16390
rect 18880 16176 18932 16182
rect 18880 16118 18932 16124
rect 20640 15978 20668 16594
rect 20628 15972 20680 15978
rect 20628 15914 20680 15920
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18892 14958 18920 15846
rect 20640 15586 20668 15914
rect 20548 15570 20668 15586
rect 20536 15564 20668 15570
rect 20588 15558 20668 15564
rect 20536 15506 20588 15512
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20732 15026 20760 15438
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 17500 14340 17552 14346
rect 17500 14282 17552 14288
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 16856 13252 16908 13258
rect 16856 13194 16908 13200
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 16868 12986 16896 13194
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16960 12986 16988 13126
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16592 12566 16712 12594
rect 16500 12406 16620 12434
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 14842 11996 15150 12005
rect 14842 11994 14848 11996
rect 14904 11994 14928 11996
rect 14984 11994 15008 11996
rect 15064 11994 15088 11996
rect 15144 11994 15150 11996
rect 14904 11942 14906 11994
rect 15086 11942 15088 11994
rect 14842 11940 14848 11942
rect 14904 11940 14928 11942
rect 14984 11940 15008 11942
rect 15064 11940 15088 11942
rect 15144 11940 15150 11942
rect 14842 11931 15150 11940
rect 14752 11852 14872 11880
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14188 11280 14240 11286
rect 14188 11222 14240 11228
rect 14200 8974 14228 11222
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 10742 14320 10950
rect 14280 10736 14332 10742
rect 14280 10678 14332 10684
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14568 10062 14596 10610
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14200 7342 14228 8910
rect 14384 8566 14412 9318
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 13924 5166 13952 5850
rect 14568 5778 14596 9998
rect 14660 9586 14688 11698
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14752 11218 14780 11630
rect 14844 11218 14872 11852
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14752 10810 14780 11154
rect 14842 10908 15150 10917
rect 14842 10906 14848 10908
rect 14904 10906 14928 10908
rect 14984 10906 15008 10908
rect 15064 10906 15088 10908
rect 15144 10906 15150 10908
rect 14904 10854 14906 10906
rect 15086 10854 15088 10906
rect 14842 10852 14848 10854
rect 14904 10852 14928 10854
rect 14984 10852 15008 10854
rect 15064 10852 15088 10854
rect 15144 10852 15150 10854
rect 14842 10843 15150 10852
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 14842 9820 15150 9829
rect 14842 9818 14848 9820
rect 14904 9818 14928 9820
rect 14984 9818 15008 9820
rect 15064 9818 15088 9820
rect 15144 9818 15150 9820
rect 14904 9766 14906 9818
rect 15086 9766 15088 9818
rect 14842 9764 14848 9766
rect 14904 9764 14928 9766
rect 14984 9764 15008 9766
rect 15064 9764 15088 9766
rect 15144 9764 15150 9766
rect 14842 9755 15150 9764
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15120 8974 15148 9522
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 14660 7954 14688 8910
rect 15384 8900 15436 8906
rect 15384 8842 15436 8848
rect 14842 8732 15150 8741
rect 14842 8730 14848 8732
rect 14904 8730 14928 8732
rect 14984 8730 15008 8732
rect 15064 8730 15088 8732
rect 15144 8730 15150 8732
rect 14904 8678 14906 8730
rect 15086 8678 15088 8730
rect 14842 8676 14848 8678
rect 14904 8676 14928 8678
rect 14984 8676 15008 8678
rect 15064 8676 15088 8678
rect 15144 8676 15150 8678
rect 14842 8667 15150 8676
rect 15396 8566 15424 8842
rect 15384 8560 15436 8566
rect 15384 8502 15436 8508
rect 15672 8090 15700 12174
rect 16592 11914 16620 12406
rect 16684 12170 16712 12566
rect 16960 12306 16988 12922
rect 17052 12442 17080 13194
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16592 11886 16712 11914
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15856 8634 15884 8910
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 14660 7410 14688 7890
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 14842 7644 15150 7653
rect 14842 7642 14848 7644
rect 14904 7642 14928 7644
rect 14984 7642 15008 7644
rect 15064 7642 15088 7644
rect 15144 7642 15150 7644
rect 14904 7590 14906 7642
rect 15086 7590 15088 7642
rect 14842 7588 14848 7590
rect 14904 7588 14928 7590
rect 14984 7588 15008 7590
rect 15064 7588 15088 7590
rect 15144 7588 15150 7590
rect 14842 7579 15150 7588
rect 15212 7478 15240 7754
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14842 6556 15150 6565
rect 14842 6554 14848 6556
rect 14904 6554 14928 6556
rect 14984 6554 15008 6556
rect 15064 6554 15088 6556
rect 15144 6554 15150 6556
rect 14904 6502 14906 6554
rect 15086 6502 15088 6554
rect 14842 6500 14848 6502
rect 14904 6500 14928 6502
rect 14984 6500 15008 6502
rect 15064 6500 15088 6502
rect 15144 6500 15150 6502
rect 14842 6491 15150 6500
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 15120 5710 15148 5850
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 14842 5468 15150 5477
rect 14842 5466 14848 5468
rect 14904 5466 14928 5468
rect 14984 5466 15008 5468
rect 15064 5466 15088 5468
rect 15144 5466 15150 5468
rect 14904 5414 14906 5466
rect 15086 5414 15088 5466
rect 14842 5412 14848 5414
rect 14904 5412 14928 5414
rect 14984 5412 15008 5414
rect 15064 5412 15088 5414
rect 15144 5412 15150 5414
rect 14842 5403 15150 5412
rect 15304 5302 15332 5510
rect 15764 5370 15792 5646
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13636 4548 13688 4554
rect 13636 4490 13688 4496
rect 13648 4214 13676 4490
rect 13636 4208 13688 4214
rect 13636 4150 13688 4156
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 12268 3602 12296 3878
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12636 3534 12664 4014
rect 13924 3534 13952 5102
rect 14292 4078 14320 5102
rect 14842 4380 15150 4389
rect 14842 4378 14848 4380
rect 14904 4378 14928 4380
rect 14984 4378 15008 4380
rect 15064 4378 15088 4380
rect 15144 4378 15150 4380
rect 14904 4326 14906 4378
rect 15086 4326 15088 4378
rect 14842 4324 14848 4326
rect 14904 4324 14928 4326
rect 14984 4324 15008 4326
rect 15064 4324 15088 4326
rect 15144 4324 15150 4326
rect 14842 4315 15150 4324
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 11369 2748 11677 2757
rect 11369 2746 11375 2748
rect 11431 2746 11455 2748
rect 11511 2746 11535 2748
rect 11591 2746 11615 2748
rect 11671 2746 11677 2748
rect 11431 2694 11433 2746
rect 11613 2694 11615 2746
rect 11369 2692 11375 2694
rect 11431 2692 11455 2694
rect 11511 2692 11535 2694
rect 11591 2692 11615 2694
rect 11671 2692 11677 2694
rect 11369 2683 11677 2692
rect 12452 2650 12480 2994
rect 12636 2990 12664 3470
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 13740 2514 13768 3470
rect 14016 3194 14044 4014
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 14660 2378 14688 3878
rect 16132 3738 16160 4014
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16592 3602 16620 11766
rect 16684 11762 16712 11886
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16684 10266 16712 11698
rect 16776 11150 16804 11834
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17144 11354 17172 11698
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 17236 10674 17264 12786
rect 17512 12782 17540 14282
rect 17604 13938 17816 13954
rect 17604 13932 17828 13938
rect 17604 13926 17776 13932
rect 17604 13870 17632 13926
rect 17776 13874 17828 13880
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 17972 13326 18000 13806
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18248 13326 18276 13670
rect 18315 13628 18623 13637
rect 18315 13626 18321 13628
rect 18377 13626 18401 13628
rect 18457 13626 18481 13628
rect 18537 13626 18561 13628
rect 18617 13626 18623 13628
rect 18377 13574 18379 13626
rect 18559 13574 18561 13626
rect 18315 13572 18321 13574
rect 18377 13572 18401 13574
rect 18457 13572 18481 13574
rect 18537 13572 18561 13574
rect 18617 13572 18623 13574
rect 18315 13563 18623 13572
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17604 12442 17632 13262
rect 17696 12918 17724 13262
rect 19444 13190 19472 13806
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 18315 12540 18623 12549
rect 18315 12538 18321 12540
rect 18377 12538 18401 12540
rect 18457 12538 18481 12540
rect 18537 12538 18561 12540
rect 18617 12538 18623 12540
rect 18377 12486 18379 12538
rect 18559 12486 18561 12538
rect 18315 12484 18321 12486
rect 18377 12484 18401 12486
rect 18457 12484 18481 12486
rect 18537 12484 18561 12486
rect 18617 12484 18623 12486
rect 18315 12475 18623 12484
rect 19444 12442 19472 12786
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19536 11558 19564 13262
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17420 10606 17448 11154
rect 18156 11150 18184 11494
rect 18315 11452 18623 11461
rect 18315 11450 18321 11452
rect 18377 11450 18401 11452
rect 18457 11450 18481 11452
rect 18537 11450 18561 11452
rect 18617 11450 18623 11452
rect 18377 11398 18379 11450
rect 18559 11398 18561 11450
rect 18315 11396 18321 11398
rect 18377 11396 18401 11398
rect 18457 11396 18481 11398
rect 18537 11396 18561 11398
rect 18617 11396 18623 11398
rect 18315 11387 18623 11396
rect 19352 11218 19380 11494
rect 19628 11354 19656 14758
rect 20364 14482 20392 14758
rect 20352 14476 20404 14482
rect 20352 14418 20404 14424
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19800 12640 19852 12646
rect 19800 12582 19852 12588
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 19812 12374 19840 12582
rect 19800 12368 19852 12374
rect 19800 12310 19852 12316
rect 19904 12306 19932 12582
rect 19892 12300 19944 12306
rect 19892 12242 19944 12248
rect 19904 11694 19932 12242
rect 19892 11688 19944 11694
rect 19892 11630 19944 11636
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19904 11354 19932 11494
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 19708 11280 19760 11286
rect 19708 11222 19760 11228
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 17408 10600 17460 10606
rect 17408 10542 17460 10548
rect 17868 10532 17920 10538
rect 17868 10474 17920 10480
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16776 10062 16804 10406
rect 17880 10266 17908 10474
rect 18315 10364 18623 10373
rect 18315 10362 18321 10364
rect 18377 10362 18401 10364
rect 18457 10362 18481 10364
rect 18537 10362 18561 10364
rect 18617 10362 18623 10364
rect 18377 10310 18379 10362
rect 18559 10310 18561 10362
rect 18315 10308 18321 10310
rect 18377 10308 18401 10310
rect 18457 10308 18481 10310
rect 18537 10308 18561 10310
rect 18617 10308 18623 10310
rect 18315 10299 18623 10308
rect 19444 10266 19472 11018
rect 19720 10742 19748 11222
rect 19708 10736 19760 10742
rect 19708 10678 19760 10684
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18524 9586 18552 9998
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19352 9654 19380 9862
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 18512 9580 18564 9586
rect 18564 9540 18736 9568
rect 18512 9522 18564 9528
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16684 7886 16712 8842
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16868 8498 16896 8774
rect 17144 8566 17172 9318
rect 18315 9276 18623 9285
rect 18315 9274 18321 9276
rect 18377 9274 18401 9276
rect 18457 9274 18481 9276
rect 18537 9274 18561 9276
rect 18617 9274 18623 9276
rect 18377 9222 18379 9274
rect 18559 9222 18561 9274
rect 18315 9220 18321 9222
rect 18377 9220 18401 9222
rect 18457 9220 18481 9222
rect 18537 9220 18561 9222
rect 18617 9220 18623 9222
rect 18315 9211 18623 9220
rect 18708 8974 18736 9540
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18800 9178 18828 9454
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18708 8634 18736 8910
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 18156 7954 18184 8502
rect 18315 8188 18623 8197
rect 18315 8186 18321 8188
rect 18377 8186 18401 8188
rect 18457 8186 18481 8188
rect 18537 8186 18561 8188
rect 18617 8186 18623 8188
rect 18377 8134 18379 8186
rect 18559 8134 18561 8186
rect 18315 8132 18321 8134
rect 18377 8132 18401 8134
rect 18457 8132 18481 8134
rect 18537 8132 18561 8134
rect 18617 8132 18623 8134
rect 18315 8123 18623 8132
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19352 7546 19380 7822
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19720 7478 19748 10678
rect 19800 9512 19852 9518
rect 19800 9454 19852 9460
rect 19812 9042 19840 9454
rect 19800 9036 19852 9042
rect 19800 8978 19852 8984
rect 19996 7954 20024 13126
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 20088 11898 20116 12242
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 20168 11756 20220 11762
rect 20168 11698 20220 11704
rect 20180 8974 20208 11698
rect 20640 11694 20668 13806
rect 20628 11688 20680 11694
rect 20628 11630 20680 11636
rect 20536 11008 20588 11014
rect 20536 10950 20588 10956
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20272 10130 20300 10406
rect 20548 10130 20576 10950
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20536 10124 20588 10130
rect 20536 10066 20588 10072
rect 20640 9654 20668 11630
rect 20732 11150 20760 14214
rect 20824 13870 20852 18702
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20916 12646 20944 15506
rect 21364 15020 21416 15026
rect 21364 14962 21416 14968
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21284 14482 21312 14758
rect 21376 14482 21404 14962
rect 21272 14476 21324 14482
rect 21272 14418 21324 14424
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21180 14340 21232 14346
rect 21180 14282 21232 14288
rect 21192 14006 21220 14282
rect 21180 14000 21232 14006
rect 21180 13942 21232 13948
rect 21560 13938 21588 21626
rect 21640 21548 21692 21554
rect 21640 21490 21692 21496
rect 21652 20806 21680 21490
rect 21824 21344 21876 21350
rect 21824 21286 21876 21292
rect 22284 21344 22336 21350
rect 22284 21286 22336 21292
rect 21836 20942 21864 21286
rect 22296 20942 22324 21286
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 22100 20936 22152 20942
rect 22284 20936 22336 20942
rect 22152 20896 22232 20924
rect 22100 20878 22152 20884
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21652 20534 21680 20742
rect 21788 20700 22096 20709
rect 21788 20698 21794 20700
rect 21850 20698 21874 20700
rect 21930 20698 21954 20700
rect 22010 20698 22034 20700
rect 22090 20698 22096 20700
rect 21850 20646 21852 20698
rect 22032 20646 22034 20698
rect 21788 20644 21794 20646
rect 21850 20644 21874 20646
rect 21930 20644 21954 20646
rect 22010 20644 22034 20646
rect 22090 20644 22096 20646
rect 21788 20635 22096 20644
rect 21640 20528 21692 20534
rect 21640 20470 21692 20476
rect 21788 19612 22096 19621
rect 21788 19610 21794 19612
rect 21850 19610 21874 19612
rect 21930 19610 21954 19612
rect 22010 19610 22034 19612
rect 22090 19610 22096 19612
rect 21850 19558 21852 19610
rect 22032 19558 22034 19610
rect 21788 19556 21794 19558
rect 21850 19556 21874 19558
rect 21930 19556 21954 19558
rect 22010 19556 22034 19558
rect 22090 19556 22096 19558
rect 21788 19547 22096 19556
rect 22204 19514 22232 20896
rect 22284 20878 22336 20884
rect 22376 20868 22428 20874
rect 22376 20810 22428 20816
rect 22388 20602 22416 20810
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22480 20398 22508 24210
rect 22560 23044 22612 23050
rect 22560 22986 22612 22992
rect 22572 22778 22600 22986
rect 22560 22772 22612 22778
rect 22560 22714 22612 22720
rect 22652 22636 22704 22642
rect 22652 22578 22704 22584
rect 22664 22094 22692 22578
rect 22572 22066 22692 22094
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22284 19780 22336 19786
rect 22284 19722 22336 19728
rect 22192 19508 22244 19514
rect 22192 19450 22244 19456
rect 21732 19440 21784 19446
rect 22296 19394 22324 19722
rect 21732 19382 21784 19388
rect 21744 18834 21772 19382
rect 22204 19378 22324 19394
rect 22192 19372 22324 19378
rect 22244 19366 22324 19372
rect 22192 19314 22244 19320
rect 22204 18902 22232 19314
rect 22572 19242 22600 22066
rect 22756 22030 22784 24686
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22756 21690 22784 21966
rect 22744 21684 22796 21690
rect 22744 21626 22796 21632
rect 22848 21554 22876 26998
rect 23020 26988 23072 26994
rect 23020 26930 23072 26936
rect 22928 26920 22980 26926
rect 22928 26862 22980 26868
rect 22940 25498 22968 26862
rect 23032 26586 23060 26930
rect 23940 26852 23992 26858
rect 23940 26794 23992 26800
rect 23388 26784 23440 26790
rect 23388 26726 23440 26732
rect 23020 26580 23072 26586
rect 23020 26522 23072 26528
rect 23112 26376 23164 26382
rect 23112 26318 23164 26324
rect 23124 26042 23152 26318
rect 23112 26036 23164 26042
rect 23112 25978 23164 25984
rect 22928 25492 22980 25498
rect 22928 25434 22980 25440
rect 23400 24886 23428 26726
rect 23952 26042 23980 26794
rect 23940 26036 23992 26042
rect 23940 25978 23992 25984
rect 24032 25832 24084 25838
rect 24032 25774 24084 25780
rect 23664 25764 23716 25770
rect 23664 25706 23716 25712
rect 23572 25696 23624 25702
rect 23572 25638 23624 25644
rect 23480 25152 23532 25158
rect 23480 25094 23532 25100
rect 23492 24954 23520 25094
rect 23480 24948 23532 24954
rect 23480 24890 23532 24896
rect 23388 24880 23440 24886
rect 23388 24822 23440 24828
rect 23584 24818 23612 25638
rect 23676 25362 23704 25706
rect 24044 25362 24072 25774
rect 23664 25356 23716 25362
rect 23664 25298 23716 25304
rect 24032 25356 24084 25362
rect 24032 25298 24084 25304
rect 23572 24812 23624 24818
rect 23572 24754 23624 24760
rect 23676 24274 23704 25298
rect 23756 25152 23808 25158
rect 23756 25094 23808 25100
rect 23664 24268 23716 24274
rect 23664 24210 23716 24216
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 23492 23866 23520 24006
rect 23480 23860 23532 23866
rect 23480 23802 23532 23808
rect 23492 23202 23520 23802
rect 23664 23248 23716 23254
rect 23492 23186 23612 23202
rect 23664 23190 23716 23196
rect 23492 23180 23624 23186
rect 23492 23174 23572 23180
rect 23572 23122 23624 23128
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 23204 21956 23256 21962
rect 23204 21898 23256 21904
rect 23216 21690 23244 21898
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 22836 21548 22888 21554
rect 22836 21490 22888 21496
rect 22848 20534 22876 21490
rect 23400 20534 23428 22714
rect 23480 21616 23532 21622
rect 23480 21558 23532 21564
rect 22836 20528 22888 20534
rect 22836 20470 22888 20476
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 22652 19916 22704 19922
rect 22652 19858 22704 19864
rect 22664 19378 22692 19858
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22928 19372 22980 19378
rect 22928 19314 22980 19320
rect 22560 19236 22612 19242
rect 22560 19178 22612 19184
rect 22192 18896 22244 18902
rect 22192 18838 22244 18844
rect 21732 18828 21784 18834
rect 21732 18770 21784 18776
rect 21640 18624 21692 18630
rect 21640 18566 21692 18572
rect 21652 17610 21680 18566
rect 21788 18524 22096 18533
rect 21788 18522 21794 18524
rect 21850 18522 21874 18524
rect 21930 18522 21954 18524
rect 22010 18522 22034 18524
rect 22090 18522 22096 18524
rect 21850 18470 21852 18522
rect 22032 18470 22034 18522
rect 21788 18468 21794 18470
rect 21850 18468 21874 18470
rect 21930 18468 21954 18470
rect 22010 18468 22034 18470
rect 22090 18468 22096 18470
rect 21788 18459 22096 18468
rect 22204 18426 22232 18838
rect 22192 18420 22244 18426
rect 22192 18362 22244 18368
rect 21640 17604 21692 17610
rect 21640 17546 21692 17552
rect 21652 15910 21680 17546
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 21788 17436 22096 17445
rect 21788 17434 21794 17436
rect 21850 17434 21874 17436
rect 21930 17434 21954 17436
rect 22010 17434 22034 17436
rect 22090 17434 22096 17436
rect 21850 17382 21852 17434
rect 22032 17382 22034 17434
rect 21788 17380 21794 17382
rect 21850 17380 21874 17382
rect 21930 17380 21954 17382
rect 22010 17380 22034 17382
rect 22090 17380 22096 17382
rect 21788 17371 22096 17380
rect 22296 17270 22324 17478
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 22664 17134 22692 19314
rect 22940 18970 22968 19314
rect 22928 18964 22980 18970
rect 22928 18906 22980 18912
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 22744 17264 22796 17270
rect 22744 17206 22796 17212
rect 22284 17128 22336 17134
rect 22284 17070 22336 17076
rect 22652 17128 22704 17134
rect 22652 17070 22704 17076
rect 22296 16658 22324 17070
rect 22284 16652 22336 16658
rect 22284 16594 22336 16600
rect 21788 16348 22096 16357
rect 21788 16346 21794 16348
rect 21850 16346 21874 16348
rect 21930 16346 21954 16348
rect 22010 16346 22034 16348
rect 22090 16346 22096 16348
rect 21850 16294 21852 16346
rect 22032 16294 22034 16346
rect 21788 16292 21794 16294
rect 21850 16292 21874 16294
rect 21930 16292 21954 16294
rect 22010 16292 22034 16294
rect 22090 16292 22096 16294
rect 21788 16283 22096 16292
rect 22296 16046 22324 16594
rect 22468 16516 22520 16522
rect 22468 16458 22520 16464
rect 22480 16182 22508 16458
rect 22756 16250 22784 17206
rect 22836 16516 22888 16522
rect 22836 16458 22888 16464
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 22468 16176 22520 16182
rect 22468 16118 22520 16124
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 22388 15502 22416 16050
rect 22848 15706 22876 16458
rect 22928 16448 22980 16454
rect 22928 16390 22980 16396
rect 22940 16250 22968 16390
rect 22928 16244 22980 16250
rect 22928 16186 22980 16192
rect 23032 16114 23060 18566
rect 23112 17740 23164 17746
rect 23112 17682 23164 17688
rect 23124 16794 23152 17682
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 22928 16108 22980 16114
rect 22928 16050 22980 16056
rect 23020 16108 23072 16114
rect 23020 16050 23072 16056
rect 22836 15700 22888 15706
rect 22836 15642 22888 15648
rect 22940 15502 22968 16050
rect 22376 15496 22428 15502
rect 22376 15438 22428 15444
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 21788 15260 22096 15269
rect 21788 15258 21794 15260
rect 21850 15258 21874 15260
rect 21930 15258 21954 15260
rect 22010 15258 22034 15260
rect 22090 15258 22096 15260
rect 21850 15206 21852 15258
rect 22032 15206 22034 15258
rect 21788 15204 21794 15206
rect 21850 15204 21874 15206
rect 21930 15204 21954 15206
rect 22010 15204 22034 15206
rect 22090 15204 22096 15206
rect 21788 15195 22096 15204
rect 21788 14172 22096 14181
rect 21788 14170 21794 14172
rect 21850 14170 21874 14172
rect 21930 14170 21954 14172
rect 22010 14170 22034 14172
rect 22090 14170 22096 14172
rect 21850 14118 21852 14170
rect 22032 14118 22034 14170
rect 21788 14116 21794 14118
rect 21850 14116 21874 14118
rect 21930 14116 21954 14118
rect 22010 14116 22034 14118
rect 22090 14116 22096 14118
rect 21788 14107 22096 14116
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 21088 13796 21140 13802
rect 21088 13738 21140 13744
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 21008 12986 21036 13262
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 21100 12918 21128 13738
rect 21088 12912 21140 12918
rect 21088 12854 21140 12860
rect 21272 12776 21324 12782
rect 21272 12718 21324 12724
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 21284 12442 21312 12718
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20824 10674 20852 12174
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 20904 11620 20956 11626
rect 20904 11562 20956 11568
rect 20916 11218 20944 11562
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20812 10668 20864 10674
rect 20812 10610 20864 10616
rect 20824 9994 20852 10610
rect 20916 10266 20944 11154
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 21284 9994 21312 11630
rect 21468 10606 21496 13874
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 21788 13084 22096 13093
rect 21788 13082 21794 13084
rect 21850 13082 21874 13084
rect 21930 13082 21954 13084
rect 22010 13082 22034 13084
rect 22090 13082 22096 13084
rect 21850 13030 21852 13082
rect 22032 13030 22034 13082
rect 21788 13028 21794 13030
rect 21850 13028 21874 13030
rect 21930 13028 21954 13030
rect 22010 13028 22034 13030
rect 22090 13028 22096 13030
rect 21788 13019 22096 13028
rect 22388 12850 22416 13126
rect 22468 12912 22520 12918
rect 22468 12854 22520 12860
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22388 12434 22416 12786
rect 22296 12406 22416 12434
rect 21788 11996 22096 12005
rect 21788 11994 21794 11996
rect 21850 11994 21874 11996
rect 21930 11994 21954 11996
rect 22010 11994 22034 11996
rect 22090 11994 22096 11996
rect 21850 11942 21852 11994
rect 22032 11942 22034 11994
rect 21788 11940 21794 11942
rect 21850 11940 21874 11942
rect 21930 11940 21954 11942
rect 22010 11940 22034 11942
rect 22090 11940 22096 11942
rect 21788 11931 22096 11940
rect 21788 10908 22096 10917
rect 21788 10906 21794 10908
rect 21850 10906 21874 10908
rect 21930 10906 21954 10908
rect 22010 10906 22034 10908
rect 22090 10906 22096 10908
rect 21850 10854 21852 10906
rect 22032 10854 22034 10906
rect 21788 10852 21794 10854
rect 21850 10852 21874 10854
rect 21930 10852 21954 10854
rect 22010 10852 22034 10854
rect 22090 10852 22096 10854
rect 21788 10843 22096 10852
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21824 10600 21876 10606
rect 21824 10542 21876 10548
rect 21836 9994 21864 10542
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 21272 9988 21324 9994
rect 21272 9930 21324 9936
rect 21824 9988 21876 9994
rect 21824 9930 21876 9936
rect 20628 9648 20680 9654
rect 20628 9590 20680 9596
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20272 8974 20300 9318
rect 20364 9042 20392 9522
rect 20824 9518 20852 9930
rect 21788 9820 22096 9829
rect 21788 9818 21794 9820
rect 21850 9818 21874 9820
rect 21930 9818 21954 9820
rect 22010 9818 22034 9820
rect 22090 9818 22096 9820
rect 21850 9766 21852 9818
rect 22032 9766 22034 9818
rect 21788 9764 21794 9766
rect 21850 9764 21874 9766
rect 21930 9764 21954 9766
rect 22010 9764 22034 9766
rect 22090 9764 22096 9766
rect 21788 9755 22096 9764
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 22296 9042 22324 12406
rect 22480 11694 22508 12854
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22572 12442 22600 12786
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 23032 12238 23060 16050
rect 23124 16046 23152 16730
rect 23112 16040 23164 16046
rect 23112 15982 23164 15988
rect 23112 13932 23164 13938
rect 23112 13874 23164 13880
rect 23124 13530 23152 13874
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 23492 13326 23520 21558
rect 23572 21344 23624 21350
rect 23572 21286 23624 21292
rect 23584 20942 23612 21286
rect 23676 21010 23704 23190
rect 23768 21622 23796 25094
rect 24044 24954 24072 25298
rect 24032 24948 24084 24954
rect 24032 24890 24084 24896
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24032 23180 24084 23186
rect 24032 23122 24084 23128
rect 24044 22234 24072 23122
rect 24032 22228 24084 22234
rect 24032 22170 24084 22176
rect 24044 21690 24072 22170
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 23756 21616 23808 21622
rect 23756 21558 23808 21564
rect 24688 21010 24716 24550
rect 24768 21412 24820 21418
rect 24768 21354 24820 21360
rect 23664 21004 23716 21010
rect 23664 20946 23716 20952
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 23572 20936 23624 20942
rect 23572 20878 23624 20884
rect 23848 20936 23900 20942
rect 23848 20878 23900 20884
rect 23860 19310 23888 20878
rect 24780 19922 24808 21354
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24768 19916 24820 19922
rect 24768 19858 24820 19864
rect 23848 19304 23900 19310
rect 23848 19246 23900 19252
rect 24032 19236 24084 19242
rect 24032 19178 24084 19184
rect 24044 18766 24072 19178
rect 24032 18760 24084 18766
rect 24032 18702 24084 18708
rect 24676 18352 24728 18358
rect 24676 18294 24728 18300
rect 24688 18170 24716 18294
rect 24872 18170 24900 20742
rect 24964 20466 24992 27270
rect 27540 27062 27568 27775
rect 27724 27470 27752 29294
rect 27802 29200 27858 29294
rect 27896 27532 27948 27538
rect 27896 27474 27948 27480
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 27528 27056 27580 27062
rect 27528 26998 27580 27004
rect 27908 26994 27936 27474
rect 28080 27396 28132 27402
rect 28080 27338 28132 27344
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 27712 26988 27764 26994
rect 27712 26930 27764 26936
rect 27896 26988 27948 26994
rect 27896 26930 27948 26936
rect 25261 26684 25569 26693
rect 25261 26682 25267 26684
rect 25323 26682 25347 26684
rect 25403 26682 25427 26684
rect 25483 26682 25507 26684
rect 25563 26682 25569 26684
rect 25323 26630 25325 26682
rect 25505 26630 25507 26682
rect 25261 26628 25267 26630
rect 25323 26628 25347 26630
rect 25403 26628 25427 26630
rect 25483 26628 25507 26630
rect 25563 26628 25569 26630
rect 25261 26619 25569 26628
rect 25792 25906 25820 26930
rect 26056 26920 26108 26926
rect 26056 26862 26108 26868
rect 26700 26920 26752 26926
rect 26700 26862 26752 26868
rect 25780 25900 25832 25906
rect 25780 25842 25832 25848
rect 26068 25838 26096 26862
rect 26712 26314 26740 26862
rect 27252 26784 27304 26790
rect 27252 26726 27304 26732
rect 27264 26450 27292 26726
rect 27724 26586 27752 26930
rect 27712 26580 27764 26586
rect 27712 26522 27764 26528
rect 27252 26444 27304 26450
rect 27252 26386 27304 26392
rect 26148 26308 26200 26314
rect 26148 26250 26200 26256
rect 26700 26308 26752 26314
rect 26700 26250 26752 26256
rect 26160 25906 26188 26250
rect 26148 25900 26200 25906
rect 26148 25842 26200 25848
rect 26056 25832 26108 25838
rect 26056 25774 26108 25780
rect 25261 25596 25569 25605
rect 25261 25594 25267 25596
rect 25323 25594 25347 25596
rect 25403 25594 25427 25596
rect 25483 25594 25507 25596
rect 25563 25594 25569 25596
rect 25323 25542 25325 25594
rect 25505 25542 25507 25594
rect 25261 25540 25267 25542
rect 25323 25540 25347 25542
rect 25403 25540 25427 25542
rect 25483 25540 25507 25542
rect 25563 25540 25569 25542
rect 25261 25531 25569 25540
rect 25044 25356 25096 25362
rect 25044 25298 25096 25304
rect 25056 24614 25084 25298
rect 25136 24812 25188 24818
rect 25136 24754 25188 24760
rect 25044 24608 25096 24614
rect 25044 24550 25096 24556
rect 25148 23322 25176 24754
rect 25261 24508 25569 24517
rect 25261 24506 25267 24508
rect 25323 24506 25347 24508
rect 25403 24506 25427 24508
rect 25483 24506 25507 24508
rect 25563 24506 25569 24508
rect 25323 24454 25325 24506
rect 25505 24454 25507 24506
rect 25261 24452 25267 24454
rect 25323 24452 25347 24454
rect 25403 24452 25427 24454
rect 25483 24452 25507 24454
rect 25563 24452 25569 24454
rect 25261 24443 25569 24452
rect 26068 23798 26096 25774
rect 26160 25362 26188 25842
rect 26516 25832 26568 25838
rect 26516 25774 26568 25780
rect 26148 25356 26200 25362
rect 26148 25298 26200 25304
rect 26528 25226 26556 25774
rect 27436 25764 27488 25770
rect 27436 25706 27488 25712
rect 26516 25220 26568 25226
rect 26516 25162 26568 25168
rect 27252 25220 27304 25226
rect 27252 25162 27304 25168
rect 26148 24812 26200 24818
rect 26148 24754 26200 24760
rect 26056 23792 26108 23798
rect 26056 23734 26108 23740
rect 26160 23730 26188 24754
rect 27264 24750 27292 25162
rect 27252 24744 27304 24750
rect 27252 24686 27304 24692
rect 27448 23730 27476 25706
rect 27528 25696 27580 25702
rect 27528 25638 27580 25644
rect 27540 25362 27568 25638
rect 27528 25356 27580 25362
rect 27528 25298 27580 25304
rect 28092 25158 28120 27338
rect 28734 27228 29042 27237
rect 28734 27226 28740 27228
rect 28796 27226 28820 27228
rect 28876 27226 28900 27228
rect 28956 27226 28980 27228
rect 29036 27226 29042 27228
rect 28796 27174 28798 27226
rect 28978 27174 28980 27226
rect 28734 27172 28740 27174
rect 28796 27172 28820 27174
rect 28876 27172 28900 27174
rect 28956 27172 28980 27174
rect 29036 27172 29042 27174
rect 28734 27163 29042 27172
rect 28734 26140 29042 26149
rect 28734 26138 28740 26140
rect 28796 26138 28820 26140
rect 28876 26138 28900 26140
rect 28956 26138 28980 26140
rect 29036 26138 29042 26140
rect 28796 26086 28798 26138
rect 28978 26086 28980 26138
rect 28734 26084 28740 26086
rect 28796 26084 28820 26086
rect 28876 26084 28900 26086
rect 28956 26084 28980 26086
rect 29036 26084 29042 26086
rect 28734 26075 29042 26084
rect 28080 25152 28132 25158
rect 28080 25094 28132 25100
rect 28734 25052 29042 25061
rect 28734 25050 28740 25052
rect 28796 25050 28820 25052
rect 28876 25050 28900 25052
rect 28956 25050 28980 25052
rect 29036 25050 29042 25052
rect 28796 24998 28798 25050
rect 28978 24998 28980 25050
rect 28734 24996 28740 24998
rect 28796 24996 28820 24998
rect 28876 24996 28900 24998
rect 28956 24996 28980 24998
rect 29036 24996 29042 24998
rect 28734 24987 29042 24996
rect 27620 24200 27672 24206
rect 27620 24142 27672 24148
rect 28170 24168 28226 24177
rect 26148 23724 26200 23730
rect 26148 23666 26200 23672
rect 27436 23724 27488 23730
rect 27436 23666 27488 23672
rect 25261 23420 25569 23429
rect 25261 23418 25267 23420
rect 25323 23418 25347 23420
rect 25403 23418 25427 23420
rect 25483 23418 25507 23420
rect 25563 23418 25569 23420
rect 25323 23366 25325 23418
rect 25505 23366 25507 23418
rect 25261 23364 25267 23366
rect 25323 23364 25347 23366
rect 25403 23364 25427 23366
rect 25483 23364 25507 23366
rect 25563 23364 25569 23366
rect 25261 23355 25569 23364
rect 26160 23322 26188 23666
rect 27344 23656 27396 23662
rect 27344 23598 27396 23604
rect 26700 23520 26752 23526
rect 26700 23462 26752 23468
rect 25136 23316 25188 23322
rect 25136 23258 25188 23264
rect 26148 23316 26200 23322
rect 26148 23258 26200 23264
rect 26712 23186 26740 23462
rect 26700 23180 26752 23186
rect 26700 23122 26752 23128
rect 26240 23112 26292 23118
rect 26240 23054 26292 23060
rect 26424 23112 26476 23118
rect 26424 23054 26476 23060
rect 26252 22642 26280 23054
rect 26436 22778 26464 23054
rect 26424 22772 26476 22778
rect 26424 22714 26476 22720
rect 26240 22636 26292 22642
rect 26240 22578 26292 22584
rect 27252 22432 27304 22438
rect 27252 22374 27304 22380
rect 25261 22332 25569 22341
rect 25261 22330 25267 22332
rect 25323 22330 25347 22332
rect 25403 22330 25427 22332
rect 25483 22330 25507 22332
rect 25563 22330 25569 22332
rect 25323 22278 25325 22330
rect 25505 22278 25507 22330
rect 25261 22276 25267 22278
rect 25323 22276 25347 22278
rect 25403 22276 25427 22278
rect 25483 22276 25507 22278
rect 25563 22276 25569 22278
rect 25261 22267 25569 22276
rect 27264 22234 27292 22374
rect 27252 22228 27304 22234
rect 27252 22170 27304 22176
rect 26240 22024 26292 22030
rect 26240 21966 26292 21972
rect 26252 21690 26280 21966
rect 26240 21684 26292 21690
rect 26240 21626 26292 21632
rect 26424 21548 26476 21554
rect 26424 21490 26476 21496
rect 26240 21480 26292 21486
rect 26240 21422 26292 21428
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 24952 20460 25004 20466
rect 24952 20402 25004 20408
rect 24964 19854 24992 20402
rect 25148 19922 25176 21286
rect 25261 21244 25569 21253
rect 25261 21242 25267 21244
rect 25323 21242 25347 21244
rect 25403 21242 25427 21244
rect 25483 21242 25507 21244
rect 25563 21242 25569 21244
rect 25323 21190 25325 21242
rect 25505 21190 25507 21242
rect 25261 21188 25267 21190
rect 25323 21188 25347 21190
rect 25403 21188 25427 21190
rect 25483 21188 25507 21190
rect 25563 21188 25569 21190
rect 25261 21179 25569 21188
rect 26252 20398 26280 21422
rect 26436 20466 26464 21490
rect 27356 21486 27384 23598
rect 27448 21554 27476 23666
rect 27528 22636 27580 22642
rect 27528 22578 27580 22584
rect 27540 22098 27568 22578
rect 27528 22092 27580 22098
rect 27528 22034 27580 22040
rect 27436 21548 27488 21554
rect 27436 21490 27488 21496
rect 27344 21480 27396 21486
rect 27344 21422 27396 21428
rect 26424 20460 26476 20466
rect 26424 20402 26476 20408
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 26240 20392 26292 20398
rect 26240 20334 26292 20340
rect 25261 20156 25569 20165
rect 25261 20154 25267 20156
rect 25323 20154 25347 20156
rect 25403 20154 25427 20156
rect 25483 20154 25507 20156
rect 25563 20154 25569 20156
rect 25323 20102 25325 20154
rect 25505 20102 25507 20154
rect 25261 20100 25267 20102
rect 25323 20100 25347 20102
rect 25403 20100 25427 20102
rect 25483 20100 25507 20102
rect 25563 20100 25569 20102
rect 25261 20091 25569 20100
rect 25136 19916 25188 19922
rect 25136 19858 25188 19864
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 25148 18698 25176 19858
rect 26252 19310 26280 20334
rect 26792 20256 26844 20262
rect 26792 20198 26844 20204
rect 26804 19922 26832 20198
rect 27356 20058 27384 20402
rect 27344 20052 27396 20058
rect 27344 19994 27396 20000
rect 26792 19916 26844 19922
rect 26792 19858 26844 19864
rect 26332 19780 26384 19786
rect 26332 19722 26384 19728
rect 26344 19378 26372 19722
rect 27448 19378 27476 21490
rect 27632 20330 27660 24142
rect 28170 24103 28172 24112
rect 28224 24103 28226 24112
rect 28172 24074 28224 24080
rect 28734 23964 29042 23973
rect 28734 23962 28740 23964
rect 28796 23962 28820 23964
rect 28876 23962 28900 23964
rect 28956 23962 28980 23964
rect 29036 23962 29042 23964
rect 28796 23910 28798 23962
rect 28978 23910 28980 23962
rect 28734 23908 28740 23910
rect 28796 23908 28820 23910
rect 28876 23908 28900 23910
rect 28956 23908 28980 23910
rect 29036 23908 29042 23910
rect 28734 23899 29042 23908
rect 27988 23656 28040 23662
rect 27988 23598 28040 23604
rect 28000 23050 28028 23598
rect 27988 23044 28040 23050
rect 27988 22986 28040 22992
rect 28734 22876 29042 22885
rect 28734 22874 28740 22876
rect 28796 22874 28820 22876
rect 28876 22874 28900 22876
rect 28956 22874 28980 22876
rect 29036 22874 29042 22876
rect 28796 22822 28798 22874
rect 28978 22822 28980 22874
rect 28734 22820 28740 22822
rect 28796 22820 28820 22822
rect 28876 22820 28900 22822
rect 28956 22820 28980 22822
rect 29036 22820 29042 22822
rect 28734 22811 29042 22820
rect 28264 21956 28316 21962
rect 28264 21898 28316 21904
rect 28276 21690 28304 21898
rect 28734 21788 29042 21797
rect 28734 21786 28740 21788
rect 28796 21786 28820 21788
rect 28876 21786 28900 21788
rect 28956 21786 28980 21788
rect 29036 21786 29042 21788
rect 28796 21734 28798 21786
rect 28978 21734 28980 21786
rect 28734 21732 28740 21734
rect 28796 21732 28820 21734
rect 28876 21732 28900 21734
rect 28956 21732 28980 21734
rect 29036 21732 29042 21734
rect 28734 21723 29042 21732
rect 28264 21684 28316 21690
rect 28264 21626 28316 21632
rect 27896 20936 27948 20942
rect 27896 20878 27948 20884
rect 27620 20324 27672 20330
rect 27620 20266 27672 20272
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 27436 19372 27488 19378
rect 27436 19314 27488 19320
rect 26240 19304 26292 19310
rect 26240 19246 26292 19252
rect 25964 19168 26016 19174
rect 25964 19110 26016 19116
rect 25261 19068 25569 19077
rect 25261 19066 25267 19068
rect 25323 19066 25347 19068
rect 25403 19066 25427 19068
rect 25483 19066 25507 19068
rect 25563 19066 25569 19068
rect 25323 19014 25325 19066
rect 25505 19014 25507 19066
rect 25261 19012 25267 19014
rect 25323 19012 25347 19014
rect 25403 19012 25427 19014
rect 25483 19012 25507 19014
rect 25563 19012 25569 19014
rect 25261 19003 25569 19012
rect 25976 18834 26004 19110
rect 25964 18828 26016 18834
rect 25964 18770 26016 18776
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 26252 18290 26280 19246
rect 26344 18970 26372 19314
rect 26332 18964 26384 18970
rect 26332 18906 26384 18912
rect 26608 18692 26660 18698
rect 26608 18634 26660 18640
rect 26620 18426 26648 18634
rect 26608 18420 26660 18426
rect 26608 18362 26660 18368
rect 25136 18284 25188 18290
rect 25136 18226 25188 18232
rect 25780 18284 25832 18290
rect 25780 18226 25832 18232
rect 26240 18284 26292 18290
rect 26240 18226 26292 18232
rect 24688 18142 24900 18170
rect 24688 17678 24716 18142
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 24872 17678 24900 18022
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 25148 17542 25176 18226
rect 25261 17980 25569 17989
rect 25261 17978 25267 17980
rect 25323 17978 25347 17980
rect 25403 17978 25427 17980
rect 25483 17978 25507 17980
rect 25563 17978 25569 17980
rect 25323 17926 25325 17978
rect 25505 17926 25507 17978
rect 25261 17924 25267 17926
rect 25323 17924 25347 17926
rect 25403 17924 25427 17926
rect 25483 17924 25507 17926
rect 25563 17924 25569 17926
rect 25261 17915 25569 17924
rect 24032 17536 24084 17542
rect 24032 17478 24084 17484
rect 25136 17536 25188 17542
rect 25136 17478 25188 17484
rect 25320 17536 25372 17542
rect 25320 17478 25372 17484
rect 24044 17270 24072 17478
rect 24032 17264 24084 17270
rect 24032 17206 24084 17212
rect 25044 17264 25096 17270
rect 25044 17206 25096 17212
rect 24492 17196 24544 17202
rect 24492 17138 24544 17144
rect 24768 17196 24820 17202
rect 24768 17138 24820 17144
rect 24032 16720 24084 16726
rect 24032 16662 24084 16668
rect 24044 16250 24072 16662
rect 24504 16590 24532 17138
rect 24780 16726 24808 17138
rect 24768 16720 24820 16726
rect 24768 16662 24820 16668
rect 25056 16590 25084 17206
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 25148 16522 25176 17478
rect 25332 17202 25360 17478
rect 25320 17196 25372 17202
rect 25320 17138 25372 17144
rect 25261 16892 25569 16901
rect 25261 16890 25267 16892
rect 25323 16890 25347 16892
rect 25403 16890 25427 16892
rect 25483 16890 25507 16892
rect 25563 16890 25569 16892
rect 25323 16838 25325 16890
rect 25505 16838 25507 16890
rect 25261 16836 25267 16838
rect 25323 16836 25347 16838
rect 25403 16836 25427 16838
rect 25483 16836 25507 16838
rect 25563 16836 25569 16838
rect 25261 16827 25569 16836
rect 25136 16516 25188 16522
rect 25136 16458 25188 16464
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 23572 13728 23624 13734
rect 23572 13670 23624 13676
rect 23584 13394 23612 13670
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 23492 11082 23520 13262
rect 23664 12640 23716 12646
rect 23664 12582 23716 12588
rect 23676 12238 23704 12582
rect 23768 12306 23796 13330
rect 23756 12300 23808 12306
rect 23756 12242 23808 12248
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23676 11694 23704 12174
rect 23664 11688 23716 11694
rect 23664 11630 23716 11636
rect 23480 11076 23532 11082
rect 23480 11018 23532 11024
rect 23664 11076 23716 11082
rect 23664 11018 23716 11024
rect 22836 11008 22888 11014
rect 22836 10950 22888 10956
rect 22848 10674 22876 10950
rect 22836 10668 22888 10674
rect 22836 10610 22888 10616
rect 23572 10464 23624 10470
rect 23572 10406 23624 10412
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 23032 9654 23060 9998
rect 23020 9648 23072 9654
rect 23020 9590 23072 9596
rect 20352 9036 20404 9042
rect 20352 8978 20404 8984
rect 22284 9036 22336 9042
rect 22284 8978 22336 8984
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 20180 7546 20208 8910
rect 21788 8732 22096 8741
rect 21788 8730 21794 8732
rect 21850 8730 21874 8732
rect 21930 8730 21954 8732
rect 22010 8730 22034 8732
rect 22090 8730 22096 8732
rect 21850 8678 21852 8730
rect 22032 8678 22034 8730
rect 21788 8676 21794 8678
rect 21850 8676 21874 8678
rect 21930 8676 21954 8678
rect 22010 8676 22034 8678
rect 22090 8676 22096 8678
rect 21788 8667 22096 8676
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 22192 7948 22244 7954
rect 22296 7936 22324 8978
rect 22756 8498 22784 8978
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 23112 8832 23164 8838
rect 23112 8774 23164 8780
rect 22848 8634 22876 8774
rect 22836 8628 22888 8634
rect 22836 8570 22888 8576
rect 23124 8566 23152 8774
rect 23112 8560 23164 8566
rect 23112 8502 23164 8508
rect 22744 8492 22796 8498
rect 22744 8434 22796 8440
rect 22244 7908 22324 7936
rect 22192 7890 22244 7896
rect 21180 7812 21232 7818
rect 21180 7754 21232 7760
rect 21192 7546 21220 7754
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 19708 7472 19760 7478
rect 19708 7414 19760 7420
rect 18315 7100 18623 7109
rect 18315 7098 18321 7100
rect 18377 7098 18401 7100
rect 18457 7098 18481 7100
rect 18537 7098 18561 7100
rect 18617 7098 18623 7100
rect 18377 7046 18379 7098
rect 18559 7046 18561 7098
rect 18315 7044 18321 7046
rect 18377 7044 18401 7046
rect 18457 7044 18481 7046
rect 18537 7044 18561 7046
rect 18617 7044 18623 7046
rect 18315 7035 18623 7044
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 16776 5370 16804 5578
rect 16868 5556 16896 6190
rect 17052 5778 17080 6258
rect 17144 5914 17172 6802
rect 21652 6798 21680 7890
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 21788 7644 22096 7653
rect 21788 7642 21794 7644
rect 21850 7642 21874 7644
rect 21930 7642 21954 7644
rect 22010 7642 22034 7644
rect 22090 7642 22096 7644
rect 21850 7590 21852 7642
rect 22032 7590 22034 7642
rect 21788 7588 21794 7590
rect 21850 7588 21874 7590
rect 21930 7588 21954 7590
rect 22010 7588 22034 7590
rect 22090 7588 22096 7590
rect 21788 7579 22096 7588
rect 22204 7410 22232 7686
rect 22480 7546 22508 7754
rect 23584 7546 23612 10406
rect 23676 8974 23704 11018
rect 23860 9042 23888 15982
rect 25261 15804 25569 15813
rect 25261 15802 25267 15804
rect 25323 15802 25347 15804
rect 25403 15802 25427 15804
rect 25483 15802 25507 15804
rect 25563 15802 25569 15804
rect 25323 15750 25325 15802
rect 25505 15750 25507 15802
rect 25261 15748 25267 15750
rect 25323 15748 25347 15750
rect 25403 15748 25427 15750
rect 25483 15748 25507 15750
rect 25563 15748 25569 15750
rect 25261 15739 25569 15748
rect 24872 15286 25084 15314
rect 24780 15094 24808 15125
rect 24768 15088 24820 15094
rect 24872 15042 24900 15286
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24820 15036 24900 15042
rect 24768 15030 24900 15036
rect 24780 15014 24900 15030
rect 24780 14074 24808 15014
rect 24964 14482 24992 15098
rect 25056 15094 25084 15286
rect 25044 15088 25096 15094
rect 25044 15030 25096 15036
rect 25261 14716 25569 14725
rect 25261 14714 25267 14716
rect 25323 14714 25347 14716
rect 25403 14714 25427 14716
rect 25483 14714 25507 14716
rect 25563 14714 25569 14716
rect 25323 14662 25325 14714
rect 25505 14662 25507 14714
rect 25261 14660 25267 14662
rect 25323 14660 25347 14662
rect 25403 14660 25427 14662
rect 25483 14660 25507 14662
rect 25563 14660 25569 14662
rect 25261 14651 25569 14660
rect 24952 14476 25004 14482
rect 24952 14418 25004 14424
rect 24768 14068 24820 14074
rect 24768 14010 24820 14016
rect 25261 13628 25569 13637
rect 25261 13626 25267 13628
rect 25323 13626 25347 13628
rect 25403 13626 25427 13628
rect 25483 13626 25507 13628
rect 25563 13626 25569 13628
rect 25323 13574 25325 13626
rect 25505 13574 25507 13626
rect 25261 13572 25267 13574
rect 25323 13572 25347 13574
rect 25403 13572 25427 13574
rect 25483 13572 25507 13574
rect 25563 13572 25569 13574
rect 25261 13563 25569 13572
rect 24584 13388 24636 13394
rect 24584 13330 24636 13336
rect 24596 12986 24624 13330
rect 24584 12980 24636 12986
rect 24584 12922 24636 12928
rect 25261 12540 25569 12549
rect 25261 12538 25267 12540
rect 25323 12538 25347 12540
rect 25403 12538 25427 12540
rect 25483 12538 25507 12540
rect 25563 12538 25569 12540
rect 25323 12486 25325 12538
rect 25505 12486 25507 12538
rect 25261 12484 25267 12486
rect 25323 12484 25347 12486
rect 25403 12484 25427 12486
rect 25483 12484 25507 12486
rect 25563 12484 25569 12486
rect 25261 12475 25569 12484
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 25056 11830 25084 12038
rect 25044 11824 25096 11830
rect 25044 11766 25096 11772
rect 25688 11824 25740 11830
rect 25688 11766 25740 11772
rect 24676 11756 24728 11762
rect 24676 11698 24728 11704
rect 23940 11552 23992 11558
rect 23940 11494 23992 11500
rect 23952 10810 23980 11494
rect 24688 11150 24716 11698
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24780 11354 24808 11630
rect 25261 11452 25569 11461
rect 25261 11450 25267 11452
rect 25323 11450 25347 11452
rect 25403 11450 25427 11452
rect 25483 11450 25507 11452
rect 25563 11450 25569 11452
rect 25323 11398 25325 11450
rect 25505 11398 25507 11450
rect 25261 11396 25267 11398
rect 25323 11396 25347 11398
rect 25403 11396 25427 11398
rect 25483 11396 25507 11398
rect 25563 11396 25569 11398
rect 25261 11387 25569 11396
rect 24768 11348 24820 11354
rect 24768 11290 24820 11296
rect 25700 11218 25728 11766
rect 25688 11212 25740 11218
rect 25688 11154 25740 11160
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24688 10810 24716 11086
rect 23940 10804 23992 10810
rect 23940 10746 23992 10752
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24124 10736 24176 10742
rect 24124 10678 24176 10684
rect 24136 10130 24164 10678
rect 25261 10364 25569 10373
rect 25261 10362 25267 10364
rect 25323 10362 25347 10364
rect 25403 10362 25427 10364
rect 25483 10362 25507 10364
rect 25563 10362 25569 10364
rect 25323 10310 25325 10362
rect 25505 10310 25507 10362
rect 25261 10308 25267 10310
rect 25323 10308 25347 10310
rect 25403 10308 25427 10310
rect 25483 10308 25507 10310
rect 25563 10308 25569 10310
rect 25261 10299 25569 10308
rect 24124 10124 24176 10130
rect 24124 10066 24176 10072
rect 25261 9276 25569 9285
rect 25261 9274 25267 9276
rect 25323 9274 25347 9276
rect 25403 9274 25427 9276
rect 25483 9274 25507 9276
rect 25563 9274 25569 9276
rect 25323 9222 25325 9274
rect 25505 9222 25507 9274
rect 25261 9220 25267 9222
rect 25323 9220 25347 9222
rect 25403 9220 25427 9222
rect 25483 9220 25507 9222
rect 25563 9220 25569 9222
rect 25261 9211 25569 9220
rect 25792 9110 25820 18226
rect 27620 17672 27672 17678
rect 27620 17614 27672 17620
rect 27252 17264 27304 17270
rect 27252 17206 27304 17212
rect 26332 17196 26384 17202
rect 26332 17138 26384 17144
rect 26884 17196 26936 17202
rect 26884 17138 26936 17144
rect 26344 16794 26372 17138
rect 26332 16788 26384 16794
rect 26332 16730 26384 16736
rect 26896 16658 26924 17138
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 26148 15496 26200 15502
rect 26148 15438 26200 15444
rect 25964 15360 26016 15366
rect 25964 15302 26016 15308
rect 25976 14482 26004 15302
rect 26160 14890 26188 15438
rect 26792 15020 26844 15026
rect 26792 14962 26844 14968
rect 26516 14952 26568 14958
rect 26516 14894 26568 14900
rect 26148 14884 26200 14890
rect 26148 14826 26200 14832
rect 26160 14618 26188 14826
rect 26148 14612 26200 14618
rect 26148 14554 26200 14560
rect 25964 14476 26016 14482
rect 25964 14418 26016 14424
rect 26528 14346 26556 14894
rect 26516 14340 26568 14346
rect 26516 14282 26568 14288
rect 26804 13938 26832 14962
rect 26424 13932 26476 13938
rect 26424 13874 26476 13880
rect 26792 13932 26844 13938
rect 26792 13874 26844 13880
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26252 13394 26280 13670
rect 26240 13388 26292 13394
rect 26240 13330 26292 13336
rect 26436 13258 26464 13874
rect 26424 13252 26476 13258
rect 26424 13194 26476 13200
rect 26436 12850 26464 13194
rect 26332 12844 26384 12850
rect 26332 12786 26384 12792
rect 26424 12844 26476 12850
rect 26424 12786 26476 12792
rect 26344 12238 26372 12786
rect 26424 12640 26476 12646
rect 26424 12582 26476 12588
rect 26700 12640 26752 12646
rect 26700 12582 26752 12588
rect 26436 12306 26464 12582
rect 26712 12306 26740 12582
rect 26424 12300 26476 12306
rect 26424 12242 26476 12248
rect 26700 12300 26752 12306
rect 26700 12242 26752 12248
rect 26332 12232 26384 12238
rect 26332 12174 26384 12180
rect 26344 11898 26372 12174
rect 26332 11892 26384 11898
rect 26332 11834 26384 11840
rect 26056 11212 26108 11218
rect 26056 11154 26108 11160
rect 26068 11054 26096 11154
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 25976 11026 26096 11054
rect 25976 9994 26004 11026
rect 26620 10198 26648 11086
rect 26608 10192 26660 10198
rect 26608 10134 26660 10140
rect 26516 10124 26568 10130
rect 26516 10066 26568 10072
rect 25964 9988 26016 9994
rect 25964 9930 26016 9936
rect 26528 9722 26556 10066
rect 26516 9716 26568 9722
rect 26516 9658 26568 9664
rect 26424 9580 26476 9586
rect 26424 9522 26476 9528
rect 26608 9580 26660 9586
rect 26608 9522 26660 9528
rect 25780 9104 25832 9110
rect 25780 9046 25832 9052
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 22468 7540 22520 7546
rect 22468 7482 22520 7488
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22664 6798 22692 7346
rect 23860 7342 23888 8978
rect 26436 8974 26464 9522
rect 26620 9042 26648 9522
rect 26896 9178 26924 16594
rect 27264 16590 27292 17206
rect 27632 16794 27660 17614
rect 27908 17338 27936 20878
rect 28172 20868 28224 20874
rect 28172 20810 28224 20816
rect 28184 20505 28212 20810
rect 28734 20700 29042 20709
rect 28734 20698 28740 20700
rect 28796 20698 28820 20700
rect 28876 20698 28900 20700
rect 28956 20698 28980 20700
rect 29036 20698 29042 20700
rect 28796 20646 28798 20698
rect 28978 20646 28980 20698
rect 28734 20644 28740 20646
rect 28796 20644 28820 20646
rect 28876 20644 28900 20646
rect 28956 20644 28980 20646
rect 29036 20644 29042 20646
rect 28734 20635 29042 20644
rect 28170 20496 28226 20505
rect 28170 20431 28226 20440
rect 28080 19780 28132 19786
rect 28080 19722 28132 19728
rect 28092 19514 28120 19722
rect 28734 19612 29042 19621
rect 28734 19610 28740 19612
rect 28796 19610 28820 19612
rect 28876 19610 28900 19612
rect 28956 19610 28980 19612
rect 29036 19610 29042 19612
rect 28796 19558 28798 19610
rect 28978 19558 28980 19610
rect 28734 19556 28740 19558
rect 28796 19556 28820 19558
rect 28876 19556 28900 19558
rect 28956 19556 28980 19558
rect 29036 19556 29042 19558
rect 28734 19547 29042 19556
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 28734 18524 29042 18533
rect 28734 18522 28740 18524
rect 28796 18522 28820 18524
rect 28876 18522 28900 18524
rect 28956 18522 28980 18524
rect 29036 18522 29042 18524
rect 28796 18470 28798 18522
rect 28978 18470 28980 18522
rect 28734 18468 28740 18470
rect 28796 18468 28820 18470
rect 28876 18468 28900 18470
rect 28956 18468 28980 18470
rect 29036 18468 29042 18470
rect 28734 18459 29042 18468
rect 28172 17604 28224 17610
rect 28172 17546 28224 17552
rect 27896 17332 27948 17338
rect 27896 17274 27948 17280
rect 28184 16833 28212 17546
rect 28734 17436 29042 17445
rect 28734 17434 28740 17436
rect 28796 17434 28820 17436
rect 28876 17434 28900 17436
rect 28956 17434 28980 17436
rect 29036 17434 29042 17436
rect 28796 17382 28798 17434
rect 28978 17382 28980 17434
rect 28734 17380 28740 17382
rect 28796 17380 28820 17382
rect 28876 17380 28900 17382
rect 28956 17380 28980 17382
rect 29036 17380 29042 17382
rect 28734 17371 29042 17380
rect 28170 16824 28226 16833
rect 27620 16788 27672 16794
rect 28170 16759 28226 16768
rect 27620 16730 27672 16736
rect 27252 16584 27304 16590
rect 27252 16526 27304 16532
rect 28734 16348 29042 16357
rect 28734 16346 28740 16348
rect 28796 16346 28820 16348
rect 28876 16346 28900 16348
rect 28956 16346 28980 16348
rect 29036 16346 29042 16348
rect 28796 16294 28798 16346
rect 28978 16294 28980 16346
rect 28734 16292 28740 16294
rect 28796 16292 28820 16294
rect 28876 16292 28900 16294
rect 28956 16292 28980 16294
rect 29036 16292 29042 16294
rect 28734 16283 29042 16292
rect 28734 15260 29042 15269
rect 28734 15258 28740 15260
rect 28796 15258 28820 15260
rect 28876 15258 28900 15260
rect 28956 15258 28980 15260
rect 29036 15258 29042 15260
rect 28796 15206 28798 15258
rect 28978 15206 28980 15258
rect 28734 15204 28740 15206
rect 28796 15204 28820 15206
rect 28876 15204 28900 15206
rect 28956 15204 28980 15206
rect 29036 15204 29042 15206
rect 28734 15195 29042 15204
rect 27988 15020 28040 15026
rect 27988 14962 28040 14968
rect 27436 14884 27488 14890
rect 27436 14826 27488 14832
rect 27252 14816 27304 14822
rect 27252 14758 27304 14764
rect 27264 13394 27292 14758
rect 27344 13932 27396 13938
rect 27344 13874 27396 13880
rect 27252 13388 27304 13394
rect 27252 13330 27304 13336
rect 27356 11762 27384 13874
rect 27448 13870 27476 14826
rect 27804 14000 27856 14006
rect 27804 13942 27856 13948
rect 27436 13864 27488 13870
rect 27436 13806 27488 13812
rect 27448 13682 27476 13806
rect 27448 13654 27568 13682
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 27448 12442 27476 12786
rect 27436 12436 27488 12442
rect 27436 12378 27488 12384
rect 27344 11756 27396 11762
rect 27344 11698 27396 11704
rect 27356 11218 27384 11698
rect 27540 11694 27568 13654
rect 27816 13258 27844 13942
rect 28000 13530 28028 14962
rect 28734 14172 29042 14181
rect 28734 14170 28740 14172
rect 28796 14170 28820 14172
rect 28876 14170 28900 14172
rect 28956 14170 28980 14172
rect 29036 14170 29042 14172
rect 28796 14118 28798 14170
rect 28978 14118 28980 14170
rect 28734 14116 28740 14118
rect 28796 14116 28820 14118
rect 28876 14116 28900 14118
rect 28956 14116 28980 14118
rect 29036 14116 29042 14118
rect 28734 14107 29042 14116
rect 27988 13524 28040 13530
rect 27988 13466 28040 13472
rect 28170 13288 28226 13297
rect 27804 13252 27856 13258
rect 28170 13223 28226 13232
rect 27804 13194 27856 13200
rect 28184 12918 28212 13223
rect 28734 13084 29042 13093
rect 28734 13082 28740 13084
rect 28796 13082 28820 13084
rect 28876 13082 28900 13084
rect 28956 13082 28980 13084
rect 29036 13082 29042 13084
rect 28796 13030 28798 13082
rect 28978 13030 28980 13082
rect 28734 13028 28740 13030
rect 28796 13028 28820 13030
rect 28876 13028 28900 13030
rect 28956 13028 28980 13030
rect 29036 13028 29042 13030
rect 28734 13019 29042 13028
rect 28172 12912 28224 12918
rect 28172 12854 28224 12860
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 27528 11688 27580 11694
rect 27528 11630 27580 11636
rect 27344 11212 27396 11218
rect 27344 11154 27396 11160
rect 27540 11150 27568 11630
rect 27528 11144 27580 11150
rect 27528 11086 27580 11092
rect 27632 10198 27660 12786
rect 27988 12164 28040 12170
rect 27988 12106 28040 12112
rect 28000 11830 28028 12106
rect 28734 11996 29042 12005
rect 28734 11994 28740 11996
rect 28796 11994 28820 11996
rect 28876 11994 28900 11996
rect 28956 11994 28980 11996
rect 29036 11994 29042 11996
rect 28796 11942 28798 11994
rect 28978 11942 28980 11994
rect 28734 11940 28740 11942
rect 28796 11940 28820 11942
rect 28876 11940 28900 11942
rect 28956 11940 28980 11942
rect 29036 11940 29042 11942
rect 28734 11931 29042 11940
rect 27988 11824 28040 11830
rect 27988 11766 28040 11772
rect 28734 10908 29042 10917
rect 28734 10906 28740 10908
rect 28796 10906 28820 10908
rect 28876 10906 28900 10908
rect 28956 10906 28980 10908
rect 29036 10906 29042 10908
rect 28796 10854 28798 10906
rect 28978 10854 28980 10906
rect 28734 10852 28740 10854
rect 28796 10852 28820 10854
rect 28876 10852 28900 10854
rect 28956 10852 28980 10854
rect 29036 10852 29042 10854
rect 28734 10843 29042 10852
rect 27896 10668 27948 10674
rect 27896 10610 27948 10616
rect 27620 10192 27672 10198
rect 27620 10134 27672 10140
rect 27620 10056 27672 10062
rect 27620 9998 27672 10004
rect 27632 9722 27660 9998
rect 27620 9716 27672 9722
rect 27620 9658 27672 9664
rect 27252 9512 27304 9518
rect 27252 9454 27304 9460
rect 26884 9172 26936 9178
rect 26884 9114 26936 9120
rect 26608 9036 26660 9042
rect 26608 8978 26660 8984
rect 27264 8974 27292 9454
rect 27804 9444 27856 9450
rect 27804 9386 27856 9392
rect 27436 9104 27488 9110
rect 27436 9046 27488 9052
rect 26424 8968 26476 8974
rect 26424 8910 26476 8916
rect 27252 8968 27304 8974
rect 27252 8910 27304 8916
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 25148 8634 25176 8774
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 24768 7880 24820 7886
rect 24768 7822 24820 7828
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 17592 6724 17644 6730
rect 17592 6666 17644 6672
rect 17604 6458 17632 6666
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 18156 6254 18184 6598
rect 18524 6322 18552 6598
rect 19444 6458 19472 6734
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19444 6322 19472 6394
rect 19536 6390 19564 6598
rect 19524 6384 19576 6390
rect 19524 6326 19576 6332
rect 20732 6322 20760 6734
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 20720 6316 20772 6322
rect 20720 6258 20772 6264
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 19524 6248 19576 6254
rect 19524 6190 19576 6196
rect 18315 6012 18623 6021
rect 18315 6010 18321 6012
rect 18377 6010 18401 6012
rect 18457 6010 18481 6012
rect 18537 6010 18561 6012
rect 18617 6010 18623 6012
rect 18377 5958 18379 6010
rect 18559 5958 18561 6010
rect 18315 5956 18321 5958
rect 18377 5956 18401 5958
rect 18457 5956 18481 5958
rect 18537 5956 18561 5958
rect 18617 5956 18623 5958
rect 18315 5947 18623 5956
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 16948 5568 17000 5574
rect 16868 5528 16948 5556
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16868 5234 16896 5528
rect 16948 5510 17000 5516
rect 17052 5234 17080 5714
rect 19536 5710 19564 6190
rect 19800 6112 19852 6118
rect 19800 6054 19852 6060
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 19812 5778 19840 6054
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 18315 4924 18623 4933
rect 18315 4922 18321 4924
rect 18377 4922 18401 4924
rect 18457 4922 18481 4924
rect 18537 4922 18561 4924
rect 18617 4922 18623 4924
rect 18377 4870 18379 4922
rect 18559 4870 18561 4922
rect 18315 4868 18321 4870
rect 18377 4868 18401 4870
rect 18457 4868 18481 4870
rect 18537 4868 18561 4870
rect 18617 4868 18623 4870
rect 18315 4859 18623 4868
rect 19536 4622 19564 5646
rect 20548 5642 20576 6054
rect 21284 5914 21312 6258
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 20536 5636 20588 5642
rect 20536 5578 20588 5584
rect 21284 4690 21312 5850
rect 21652 5710 21680 6734
rect 21788 6556 22096 6565
rect 21788 6554 21794 6556
rect 21850 6554 21874 6556
rect 21930 6554 21954 6556
rect 22010 6554 22034 6556
rect 22090 6554 22096 6556
rect 21850 6502 21852 6554
rect 22032 6502 22034 6554
rect 21788 6500 21794 6502
rect 21850 6500 21874 6502
rect 21930 6500 21954 6502
rect 22010 6500 22034 6502
rect 22090 6500 22096 6502
rect 21788 6491 22096 6500
rect 22664 6254 22692 6734
rect 22652 6248 22704 6254
rect 22652 6190 22704 6196
rect 22100 6112 22152 6118
rect 22100 6054 22152 6060
rect 22112 5710 22140 6054
rect 21640 5704 21692 5710
rect 21560 5652 21640 5658
rect 21560 5646 21692 5652
rect 22100 5704 22152 5710
rect 22152 5664 22232 5692
rect 22100 5646 22152 5652
rect 21560 5630 21680 5646
rect 21560 5234 21588 5630
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 21548 5228 21600 5234
rect 21548 5170 21600 5176
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 19524 4616 19576 4622
rect 19524 4558 19576 4564
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 17236 3534 17264 4082
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 18315 3836 18623 3845
rect 18315 3834 18321 3836
rect 18377 3834 18401 3836
rect 18457 3834 18481 3836
rect 18537 3834 18561 3836
rect 18617 3834 18623 3836
rect 18377 3782 18379 3834
rect 18559 3782 18561 3834
rect 18315 3780 18321 3782
rect 18377 3780 18401 3782
rect 18457 3780 18481 3782
rect 18537 3780 18561 3782
rect 18617 3780 18623 3782
rect 18315 3771 18623 3780
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14752 3194 14780 3334
rect 14842 3292 15150 3301
rect 14842 3290 14848 3292
rect 14904 3290 14928 3292
rect 14984 3290 15008 3292
rect 15064 3290 15088 3292
rect 15144 3290 15150 3292
rect 14904 3238 14906 3290
rect 15086 3238 15088 3290
rect 14842 3236 14848 3238
rect 14904 3236 14928 3238
rect 14984 3236 15008 3238
rect 15064 3236 15088 3238
rect 15144 3236 15150 3238
rect 14842 3227 15150 3236
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 16316 2990 16344 3470
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17972 3126 18000 3334
rect 19536 3194 19564 3538
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 19628 3194 19656 3470
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19616 3188 19668 3194
rect 19616 3130 19668 3136
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 19720 2990 19748 3878
rect 19812 3738 19840 3878
rect 19996 3738 20024 4082
rect 20640 4078 20668 4558
rect 21652 4554 21680 5510
rect 21788 5468 22096 5477
rect 21788 5466 21794 5468
rect 21850 5466 21874 5468
rect 21930 5466 21954 5468
rect 22010 5466 22034 5468
rect 22090 5466 22096 5468
rect 21850 5414 21852 5466
rect 22032 5414 22034 5466
rect 21788 5412 21794 5414
rect 21850 5412 21874 5414
rect 21930 5412 21954 5414
rect 22010 5412 22034 5414
rect 22090 5412 22096 5414
rect 21788 5403 22096 5412
rect 22204 5234 22232 5664
rect 22192 5228 22244 5234
rect 22192 5170 22244 5176
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 21640 4548 21692 4554
rect 21640 4490 21692 4496
rect 22192 4480 22244 4486
rect 22192 4422 22244 4428
rect 21788 4380 22096 4389
rect 21788 4378 21794 4380
rect 21850 4378 21874 4380
rect 21930 4378 21954 4380
rect 22010 4378 22034 4380
rect 22090 4378 22096 4380
rect 21850 4326 21852 4378
rect 22032 4326 22034 4378
rect 21788 4324 21794 4326
rect 21850 4324 21874 4326
rect 21930 4324 21954 4326
rect 22010 4324 22034 4326
rect 22090 4324 22096 4326
rect 21788 4315 22096 4324
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 20640 3534 20668 4014
rect 22204 3602 22232 4422
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20640 3058 20668 3470
rect 22296 3466 22324 4966
rect 22664 4622 22692 6190
rect 24780 6118 24808 7822
rect 25044 7472 25096 7478
rect 25044 7414 25096 7420
rect 25056 7206 25084 7414
rect 25148 7410 25176 8570
rect 25261 8188 25569 8197
rect 25261 8186 25267 8188
rect 25323 8186 25347 8188
rect 25403 8186 25427 8188
rect 25483 8186 25507 8188
rect 25563 8186 25569 8188
rect 25323 8134 25325 8186
rect 25505 8134 25507 8186
rect 25261 8132 25267 8134
rect 25323 8132 25347 8134
rect 25403 8132 25427 8134
rect 25483 8132 25507 8134
rect 25563 8132 25569 8134
rect 25261 8123 25569 8132
rect 26436 7868 26464 8910
rect 27264 8090 27292 8910
rect 27448 8430 27476 9046
rect 27816 8974 27844 9386
rect 27804 8968 27856 8974
rect 27804 8910 27856 8916
rect 27528 8492 27580 8498
rect 27528 8434 27580 8440
rect 27436 8424 27488 8430
rect 27436 8366 27488 8372
rect 27252 8084 27304 8090
rect 27252 8026 27304 8032
rect 26436 7840 26556 7868
rect 25964 7812 26016 7818
rect 25964 7754 26016 7760
rect 25412 7744 25464 7750
rect 25412 7686 25464 7692
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25424 7546 25452 7686
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25424 7410 25452 7482
rect 25136 7404 25188 7410
rect 25136 7346 25188 7352
rect 25412 7404 25464 7410
rect 25412 7346 25464 7352
rect 25044 7200 25096 7206
rect 25044 7142 25096 7148
rect 25056 6458 25084 7142
rect 25261 7100 25569 7109
rect 25261 7098 25267 7100
rect 25323 7098 25347 7100
rect 25403 7098 25427 7100
rect 25483 7098 25507 7100
rect 25563 7098 25569 7100
rect 25323 7046 25325 7098
rect 25505 7046 25507 7098
rect 25261 7044 25267 7046
rect 25323 7044 25347 7046
rect 25403 7044 25427 7046
rect 25483 7044 25507 7046
rect 25563 7044 25569 7046
rect 25261 7035 25569 7044
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 25261 6012 25569 6021
rect 25261 6010 25267 6012
rect 25323 6010 25347 6012
rect 25403 6010 25427 6012
rect 25483 6010 25507 6012
rect 25563 6010 25569 6012
rect 25323 5958 25325 6010
rect 25505 5958 25507 6010
rect 25261 5956 25267 5958
rect 25323 5956 25347 5958
rect 25403 5956 25427 5958
rect 25483 5956 25507 5958
rect 25563 5956 25569 5958
rect 25261 5947 25569 5956
rect 25700 5370 25728 7686
rect 25976 7274 26004 7754
rect 26424 7744 26476 7750
rect 26422 7712 26424 7721
rect 26476 7712 26478 7721
rect 26344 7670 26422 7698
rect 26344 7410 26372 7670
rect 26422 7647 26478 7656
rect 26528 7546 26556 7840
rect 26608 7744 26660 7750
rect 26608 7686 26660 7692
rect 26424 7540 26476 7546
rect 26424 7482 26476 7488
rect 26516 7540 26568 7546
rect 26516 7482 26568 7488
rect 26332 7404 26384 7410
rect 26332 7346 26384 7352
rect 25964 7268 26016 7274
rect 25964 7210 26016 7216
rect 25688 5364 25740 5370
rect 25688 5306 25740 5312
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 22652 4616 22704 4622
rect 22652 4558 22704 4564
rect 22284 3460 22336 3466
rect 22284 3402 22336 3408
rect 21788 3292 22096 3301
rect 21788 3290 21794 3292
rect 21850 3290 21874 3292
rect 21930 3290 21954 3292
rect 22010 3290 22034 3292
rect 22090 3290 22096 3292
rect 21850 3238 21852 3290
rect 22032 3238 22034 3290
rect 21788 3236 21794 3238
rect 21850 3236 21874 3238
rect 21930 3236 21954 3238
rect 22010 3236 22034 3238
rect 22090 3236 22096 3238
rect 21788 3227 22096 3236
rect 22756 3126 22784 4966
rect 25261 4924 25569 4933
rect 25261 4922 25267 4924
rect 25323 4922 25347 4924
rect 25403 4922 25427 4924
rect 25483 4922 25507 4924
rect 25563 4922 25569 4924
rect 25323 4870 25325 4922
rect 25505 4870 25507 4922
rect 25261 4868 25267 4870
rect 25323 4868 25347 4870
rect 25403 4868 25427 4870
rect 25483 4868 25507 4870
rect 25563 4868 25569 4870
rect 25261 4859 25569 4868
rect 23296 4616 23348 4622
rect 23296 4558 23348 4564
rect 22928 4548 22980 4554
rect 22928 4490 22980 4496
rect 22940 3738 22968 4490
rect 22928 3732 22980 3738
rect 22928 3674 22980 3680
rect 22744 3120 22796 3126
rect 22744 3062 22796 3068
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 20640 2854 20668 2994
rect 22940 2990 22968 3674
rect 23308 2990 23336 4558
rect 25596 4548 25648 4554
rect 25596 4490 25648 4496
rect 25608 4146 25636 4490
rect 25700 4486 25728 5306
rect 25976 5166 26004 7210
rect 26436 6730 26464 7482
rect 26516 7404 26568 7410
rect 26516 7346 26568 7352
rect 26528 7206 26556 7346
rect 26516 7200 26568 7206
rect 26516 7142 26568 7148
rect 26424 6724 26476 6730
rect 26424 6666 26476 6672
rect 26436 5574 26464 6666
rect 26620 6662 26648 7686
rect 26608 6656 26660 6662
rect 26608 6598 26660 6604
rect 27252 5636 27304 5642
rect 27252 5578 27304 5584
rect 26424 5568 26476 5574
rect 26424 5510 26476 5516
rect 26436 5302 26464 5510
rect 27264 5370 27292 5578
rect 27252 5364 27304 5370
rect 27252 5306 27304 5312
rect 26424 5296 26476 5302
rect 26424 5238 26476 5244
rect 26148 5228 26200 5234
rect 26148 5170 26200 5176
rect 26332 5228 26384 5234
rect 26332 5170 26384 5176
rect 25964 5160 26016 5166
rect 25964 5102 26016 5108
rect 25976 4622 26004 5102
rect 25964 4616 26016 4622
rect 25964 4558 26016 4564
rect 25688 4480 25740 4486
rect 25688 4422 25740 4428
rect 25964 4480 26016 4486
rect 25964 4422 26016 4428
rect 25700 4214 25728 4422
rect 25688 4208 25740 4214
rect 25688 4150 25740 4156
rect 25976 4146 26004 4422
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 25596 4140 25648 4146
rect 25596 4082 25648 4088
rect 25964 4140 26016 4146
rect 25964 4082 26016 4088
rect 24688 3738 24716 4082
rect 25608 3942 25636 4082
rect 25596 3936 25648 3942
rect 25596 3878 25648 3884
rect 25261 3836 25569 3845
rect 25261 3834 25267 3836
rect 25323 3834 25347 3836
rect 25403 3834 25427 3836
rect 25483 3834 25507 3836
rect 25563 3834 25569 3836
rect 25323 3782 25325 3834
rect 25505 3782 25507 3834
rect 25261 3780 25267 3782
rect 25323 3780 25347 3782
rect 25403 3780 25427 3782
rect 25483 3780 25507 3782
rect 25563 3780 25569 3782
rect 25261 3771 25569 3780
rect 24676 3732 24728 3738
rect 24676 3674 24728 3680
rect 25608 3534 25636 3878
rect 25596 3528 25648 3534
rect 25596 3470 25648 3476
rect 25608 3058 25636 3470
rect 25976 3194 26004 4082
rect 26160 4078 26188 5170
rect 26344 4826 26372 5170
rect 26700 5024 26752 5030
rect 26700 4966 26752 4972
rect 26332 4820 26384 4826
rect 26332 4762 26384 4768
rect 26240 4616 26292 4622
rect 26240 4558 26292 4564
rect 26252 4146 26280 4558
rect 26712 4486 26740 4966
rect 27448 4826 27476 8366
rect 27540 7546 27568 8434
rect 27816 8090 27844 8910
rect 27908 8634 27936 10610
rect 28172 10600 28224 10606
rect 28172 10542 28224 10548
rect 28184 9489 28212 10542
rect 28734 9820 29042 9829
rect 28734 9818 28740 9820
rect 28796 9818 28820 9820
rect 28876 9818 28900 9820
rect 28956 9818 28980 9820
rect 29036 9818 29042 9820
rect 28796 9766 28798 9818
rect 28978 9766 28980 9818
rect 28734 9764 28740 9766
rect 28796 9764 28820 9766
rect 28876 9764 28900 9766
rect 28956 9764 28980 9766
rect 29036 9764 29042 9766
rect 28734 9755 29042 9764
rect 28170 9480 28226 9489
rect 28170 9415 28226 9424
rect 28356 8900 28408 8906
rect 28356 8842 28408 8848
rect 27896 8628 27948 8634
rect 27896 8570 27948 8576
rect 28368 8498 28396 8842
rect 28734 8732 29042 8741
rect 28734 8730 28740 8732
rect 28796 8730 28820 8732
rect 28876 8730 28900 8732
rect 28956 8730 28980 8732
rect 29036 8730 29042 8732
rect 28796 8678 28798 8730
rect 28978 8678 28980 8730
rect 28734 8676 28740 8678
rect 28796 8676 28820 8678
rect 28876 8676 28900 8678
rect 28956 8676 28980 8678
rect 29036 8676 29042 8678
rect 28734 8667 29042 8676
rect 28356 8492 28408 8498
rect 28356 8434 28408 8440
rect 27804 8084 27856 8090
rect 27804 8026 27856 8032
rect 27988 7880 28040 7886
rect 27988 7822 28040 7828
rect 27620 7744 27672 7750
rect 27618 7712 27620 7721
rect 27672 7712 27674 7721
rect 27618 7647 27674 7656
rect 27528 7540 27580 7546
rect 27528 7482 27580 7488
rect 28000 7410 28028 7822
rect 28734 7644 29042 7653
rect 28734 7642 28740 7644
rect 28796 7642 28820 7644
rect 28876 7642 28900 7644
rect 28956 7642 28980 7644
rect 29036 7642 29042 7644
rect 28796 7590 28798 7642
rect 28978 7590 28980 7642
rect 28734 7588 28740 7590
rect 28796 7588 28820 7590
rect 28876 7588 28900 7590
rect 28956 7588 28980 7590
rect 29036 7588 29042 7590
rect 28734 7579 29042 7588
rect 27988 7404 28040 7410
rect 27988 7346 28040 7352
rect 28000 7002 28028 7346
rect 28080 7200 28132 7206
rect 28080 7142 28132 7148
rect 27988 6996 28040 7002
rect 27988 6938 28040 6944
rect 28092 6798 28120 7142
rect 28080 6792 28132 6798
rect 28080 6734 28132 6740
rect 28734 6556 29042 6565
rect 28734 6554 28740 6556
rect 28796 6554 28820 6556
rect 28876 6554 28900 6556
rect 28956 6554 28980 6556
rect 29036 6554 29042 6556
rect 28796 6502 28798 6554
rect 28978 6502 28980 6554
rect 28734 6500 28740 6502
rect 28796 6500 28820 6502
rect 28876 6500 28900 6502
rect 28956 6500 28980 6502
rect 29036 6500 29042 6502
rect 28734 6491 29042 6500
rect 27896 6316 27948 6322
rect 27896 6258 27948 6264
rect 27804 5704 27856 5710
rect 27804 5646 27856 5652
rect 27816 5370 27844 5646
rect 27804 5364 27856 5370
rect 27804 5306 27856 5312
rect 27528 5228 27580 5234
rect 27528 5170 27580 5176
rect 27252 4820 27304 4826
rect 27252 4762 27304 4768
rect 27436 4820 27488 4826
rect 27436 4762 27488 4768
rect 26700 4480 26752 4486
rect 26700 4422 26752 4428
rect 27264 4146 27292 4762
rect 27436 4548 27488 4554
rect 27436 4490 27488 4496
rect 26240 4140 26292 4146
rect 26240 4082 26292 4088
rect 27252 4140 27304 4146
rect 27252 4082 27304 4088
rect 26148 4072 26200 4078
rect 26148 4014 26200 4020
rect 26160 3738 26188 4014
rect 27160 3936 27212 3942
rect 27160 3878 27212 3884
rect 26148 3732 26200 3738
rect 26148 3674 26200 3680
rect 25964 3188 26016 3194
rect 25964 3130 26016 3136
rect 27172 3058 27200 3878
rect 27252 3528 27304 3534
rect 27252 3470 27304 3476
rect 27264 3194 27292 3470
rect 27252 3188 27304 3194
rect 27252 3130 27304 3136
rect 27448 3058 27476 4490
rect 27540 4146 27568 5170
rect 27908 4826 27936 6258
rect 28172 6248 28224 6254
rect 28172 6190 28224 6196
rect 28184 5817 28212 6190
rect 28170 5808 28226 5817
rect 28170 5743 28226 5752
rect 28734 5468 29042 5477
rect 28734 5466 28740 5468
rect 28796 5466 28820 5468
rect 28876 5466 28900 5468
rect 28956 5466 28980 5468
rect 29036 5466 29042 5468
rect 28796 5414 28798 5466
rect 28978 5414 28980 5466
rect 28734 5412 28740 5414
rect 28796 5412 28820 5414
rect 28876 5412 28900 5414
rect 28956 5412 28980 5414
rect 29036 5412 29042 5414
rect 28734 5403 29042 5412
rect 27896 4820 27948 4826
rect 27896 4762 27948 4768
rect 28264 4684 28316 4690
rect 28264 4626 28316 4632
rect 27712 4616 27764 4622
rect 27712 4558 27764 4564
rect 27724 4282 27752 4558
rect 28276 4282 28304 4626
rect 28356 4480 28408 4486
rect 28356 4422 28408 4428
rect 27712 4276 27764 4282
rect 27712 4218 27764 4224
rect 28264 4276 28316 4282
rect 28264 4218 28316 4224
rect 28368 4146 28396 4422
rect 28734 4380 29042 4389
rect 28734 4378 28740 4380
rect 28796 4378 28820 4380
rect 28876 4378 28900 4380
rect 28956 4378 28980 4380
rect 29036 4378 29042 4380
rect 28796 4326 28798 4378
rect 28978 4326 28980 4378
rect 28734 4324 28740 4326
rect 28796 4324 28820 4326
rect 28876 4324 28900 4326
rect 28956 4324 28980 4326
rect 29036 4324 29042 4326
rect 28734 4315 29042 4324
rect 27528 4140 27580 4146
rect 27528 4082 27580 4088
rect 28356 4140 28408 4146
rect 28356 4082 28408 4088
rect 27540 3534 27568 4082
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 28734 3292 29042 3301
rect 28734 3290 28740 3292
rect 28796 3290 28820 3292
rect 28876 3290 28900 3292
rect 28956 3290 28980 3292
rect 29036 3290 29042 3292
rect 28796 3238 28798 3290
rect 28978 3238 28980 3290
rect 28734 3236 28740 3238
rect 28796 3236 28820 3238
rect 28876 3236 28900 3238
rect 28956 3236 28980 3238
rect 29036 3236 29042 3238
rect 28734 3227 29042 3236
rect 25596 3052 25648 3058
rect 25596 2994 25648 3000
rect 27160 3052 27212 3058
rect 27160 2994 27212 3000
rect 27436 3052 27488 3058
rect 27436 2994 27488 3000
rect 22928 2984 22980 2990
rect 22928 2926 22980 2932
rect 23296 2984 23348 2990
rect 23296 2926 23348 2932
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 27896 2848 27948 2854
rect 27896 2790 27948 2796
rect 18315 2748 18623 2757
rect 18315 2746 18321 2748
rect 18377 2746 18401 2748
rect 18457 2746 18481 2748
rect 18537 2746 18561 2748
rect 18617 2746 18623 2748
rect 18377 2694 18379 2746
rect 18559 2694 18561 2746
rect 18315 2692 18321 2694
rect 18377 2692 18401 2694
rect 18457 2692 18481 2694
rect 18537 2692 18561 2694
rect 18617 2692 18623 2694
rect 18315 2683 18623 2692
rect 25261 2748 25569 2757
rect 25261 2746 25267 2748
rect 25323 2746 25347 2748
rect 25403 2746 25427 2748
rect 25483 2746 25507 2748
rect 25563 2746 25569 2748
rect 25323 2694 25325 2746
rect 25505 2694 25507 2746
rect 25261 2692 25267 2694
rect 25323 2692 25347 2694
rect 25403 2692 25427 2694
rect 25483 2692 25507 2694
rect 25563 2692 25569 2694
rect 25261 2683 25569 2692
rect 27908 2446 27936 2790
rect 27896 2440 27948 2446
rect 27896 2382 27948 2388
rect 28170 2408 28226 2417
rect 14648 2372 14700 2378
rect 28170 2343 28172 2352
rect 14648 2314 14700 2320
rect 28224 2343 28226 2352
rect 28172 2314 28224 2320
rect 7896 2204 8204 2213
rect 7896 2202 7902 2204
rect 7958 2202 7982 2204
rect 8038 2202 8062 2204
rect 8118 2202 8142 2204
rect 8198 2202 8204 2204
rect 7958 2150 7960 2202
rect 8140 2150 8142 2202
rect 7896 2148 7902 2150
rect 7958 2148 7982 2150
rect 8038 2148 8062 2150
rect 8118 2148 8142 2150
rect 8198 2148 8204 2150
rect 7896 2139 8204 2148
rect 14842 2204 15150 2213
rect 14842 2202 14848 2204
rect 14904 2202 14928 2204
rect 14984 2202 15008 2204
rect 15064 2202 15088 2204
rect 15144 2202 15150 2204
rect 14904 2150 14906 2202
rect 15086 2150 15088 2202
rect 14842 2148 14848 2150
rect 14904 2148 14928 2150
rect 14984 2148 15008 2150
rect 15064 2148 15088 2150
rect 15144 2148 15150 2150
rect 14842 2139 15150 2148
rect 21788 2204 22096 2213
rect 21788 2202 21794 2204
rect 21850 2202 21874 2204
rect 21930 2202 21954 2204
rect 22010 2202 22034 2204
rect 22090 2202 22096 2204
rect 21850 2150 21852 2202
rect 22032 2150 22034 2202
rect 21788 2148 21794 2150
rect 21850 2148 21874 2150
rect 21930 2148 21954 2150
rect 22010 2148 22034 2150
rect 22090 2148 22096 2150
rect 21788 2139 22096 2148
rect 28734 2204 29042 2213
rect 28734 2202 28740 2204
rect 28796 2202 28820 2204
rect 28876 2202 28900 2204
rect 28956 2202 28980 2204
rect 29036 2202 29042 2204
rect 28796 2150 28798 2202
rect 28978 2150 28980 2202
rect 28734 2148 28740 2150
rect 28796 2148 28820 2150
rect 28876 2148 28900 2150
rect 28956 2148 28980 2150
rect 29036 2148 29042 2150
rect 28734 2139 29042 2148
<< via2 >>
rect 4429 27770 4485 27772
rect 4509 27770 4565 27772
rect 4589 27770 4645 27772
rect 4669 27770 4725 27772
rect 4429 27718 4475 27770
rect 4475 27718 4485 27770
rect 4509 27718 4539 27770
rect 4539 27718 4551 27770
rect 4551 27718 4565 27770
rect 4589 27718 4603 27770
rect 4603 27718 4615 27770
rect 4615 27718 4645 27770
rect 4669 27718 4679 27770
rect 4679 27718 4725 27770
rect 4429 27716 4485 27718
rect 4509 27716 4565 27718
rect 4589 27716 4645 27718
rect 4669 27716 4725 27718
rect 11375 27770 11431 27772
rect 11455 27770 11511 27772
rect 11535 27770 11591 27772
rect 11615 27770 11671 27772
rect 11375 27718 11421 27770
rect 11421 27718 11431 27770
rect 11455 27718 11485 27770
rect 11485 27718 11497 27770
rect 11497 27718 11511 27770
rect 11535 27718 11549 27770
rect 11549 27718 11561 27770
rect 11561 27718 11591 27770
rect 11615 27718 11625 27770
rect 11625 27718 11671 27770
rect 11375 27716 11431 27718
rect 11455 27716 11511 27718
rect 11535 27716 11591 27718
rect 11615 27716 11671 27718
rect 18321 27770 18377 27772
rect 18401 27770 18457 27772
rect 18481 27770 18537 27772
rect 18561 27770 18617 27772
rect 18321 27718 18367 27770
rect 18367 27718 18377 27770
rect 18401 27718 18431 27770
rect 18431 27718 18443 27770
rect 18443 27718 18457 27770
rect 18481 27718 18495 27770
rect 18495 27718 18507 27770
rect 18507 27718 18537 27770
rect 18561 27718 18571 27770
rect 18571 27718 18617 27770
rect 18321 27716 18377 27718
rect 18401 27716 18457 27718
rect 18481 27716 18537 27718
rect 18561 27716 18617 27718
rect 4429 26682 4485 26684
rect 4509 26682 4565 26684
rect 4589 26682 4645 26684
rect 4669 26682 4725 26684
rect 4429 26630 4475 26682
rect 4475 26630 4485 26682
rect 4509 26630 4539 26682
rect 4539 26630 4551 26682
rect 4551 26630 4565 26682
rect 4589 26630 4603 26682
rect 4603 26630 4615 26682
rect 4615 26630 4645 26682
rect 4669 26630 4679 26682
rect 4679 26630 4725 26682
rect 4429 26628 4485 26630
rect 4509 26628 4565 26630
rect 4589 26628 4645 26630
rect 4669 26628 4725 26630
rect 4429 25594 4485 25596
rect 4509 25594 4565 25596
rect 4589 25594 4645 25596
rect 4669 25594 4725 25596
rect 4429 25542 4475 25594
rect 4475 25542 4485 25594
rect 4509 25542 4539 25594
rect 4539 25542 4551 25594
rect 4551 25542 4565 25594
rect 4589 25542 4603 25594
rect 4603 25542 4615 25594
rect 4615 25542 4645 25594
rect 4669 25542 4679 25594
rect 4679 25542 4725 25594
rect 4429 25540 4485 25542
rect 4509 25540 4565 25542
rect 4589 25540 4645 25542
rect 4669 25540 4725 25542
rect 7902 27226 7958 27228
rect 7982 27226 8038 27228
rect 8062 27226 8118 27228
rect 8142 27226 8198 27228
rect 7902 27174 7948 27226
rect 7948 27174 7958 27226
rect 7982 27174 8012 27226
rect 8012 27174 8024 27226
rect 8024 27174 8038 27226
rect 8062 27174 8076 27226
rect 8076 27174 8088 27226
rect 8088 27174 8118 27226
rect 8142 27174 8152 27226
rect 8152 27174 8198 27226
rect 7902 27172 7958 27174
rect 7982 27172 8038 27174
rect 8062 27172 8118 27174
rect 8142 27172 8198 27174
rect 4429 24506 4485 24508
rect 4509 24506 4565 24508
rect 4589 24506 4645 24508
rect 4669 24506 4725 24508
rect 4429 24454 4475 24506
rect 4475 24454 4485 24506
rect 4509 24454 4539 24506
rect 4539 24454 4551 24506
rect 4551 24454 4565 24506
rect 4589 24454 4603 24506
rect 4603 24454 4615 24506
rect 4615 24454 4645 24506
rect 4669 24454 4679 24506
rect 4679 24454 4725 24506
rect 4429 24452 4485 24454
rect 4509 24452 4565 24454
rect 4589 24452 4645 24454
rect 4669 24452 4725 24454
rect 4429 23418 4485 23420
rect 4509 23418 4565 23420
rect 4589 23418 4645 23420
rect 4669 23418 4725 23420
rect 4429 23366 4475 23418
rect 4475 23366 4485 23418
rect 4509 23366 4539 23418
rect 4539 23366 4551 23418
rect 4551 23366 4565 23418
rect 4589 23366 4603 23418
rect 4603 23366 4615 23418
rect 4615 23366 4645 23418
rect 4669 23366 4679 23418
rect 4679 23366 4725 23418
rect 4429 23364 4485 23366
rect 4509 23364 4565 23366
rect 4589 23364 4645 23366
rect 4669 23364 4725 23366
rect 4429 22330 4485 22332
rect 4509 22330 4565 22332
rect 4589 22330 4645 22332
rect 4669 22330 4725 22332
rect 4429 22278 4475 22330
rect 4475 22278 4485 22330
rect 4509 22278 4539 22330
rect 4539 22278 4551 22330
rect 4551 22278 4565 22330
rect 4589 22278 4603 22330
rect 4603 22278 4615 22330
rect 4615 22278 4645 22330
rect 4669 22278 4679 22330
rect 4679 22278 4725 22330
rect 4429 22276 4485 22278
rect 4509 22276 4565 22278
rect 4589 22276 4645 22278
rect 4669 22276 4725 22278
rect 4429 21242 4485 21244
rect 4509 21242 4565 21244
rect 4589 21242 4645 21244
rect 4669 21242 4725 21244
rect 4429 21190 4475 21242
rect 4475 21190 4485 21242
rect 4509 21190 4539 21242
rect 4539 21190 4551 21242
rect 4551 21190 4565 21242
rect 4589 21190 4603 21242
rect 4603 21190 4615 21242
rect 4615 21190 4645 21242
rect 4669 21190 4679 21242
rect 4679 21190 4725 21242
rect 4429 21188 4485 21190
rect 4509 21188 4565 21190
rect 4589 21188 4645 21190
rect 4669 21188 4725 21190
rect 4429 20154 4485 20156
rect 4509 20154 4565 20156
rect 4589 20154 4645 20156
rect 4669 20154 4725 20156
rect 4429 20102 4475 20154
rect 4475 20102 4485 20154
rect 4509 20102 4539 20154
rect 4539 20102 4551 20154
rect 4551 20102 4565 20154
rect 4589 20102 4603 20154
rect 4603 20102 4615 20154
rect 4615 20102 4645 20154
rect 4669 20102 4679 20154
rect 4679 20102 4725 20154
rect 4429 20100 4485 20102
rect 4509 20100 4565 20102
rect 4589 20100 4645 20102
rect 4669 20100 4725 20102
rect 4429 19066 4485 19068
rect 4509 19066 4565 19068
rect 4589 19066 4645 19068
rect 4669 19066 4725 19068
rect 4429 19014 4475 19066
rect 4475 19014 4485 19066
rect 4509 19014 4539 19066
rect 4539 19014 4551 19066
rect 4551 19014 4565 19066
rect 4589 19014 4603 19066
rect 4603 19014 4615 19066
rect 4615 19014 4645 19066
rect 4669 19014 4679 19066
rect 4679 19014 4725 19066
rect 4429 19012 4485 19014
rect 4509 19012 4565 19014
rect 4589 19012 4645 19014
rect 4669 19012 4725 19014
rect 4429 17978 4485 17980
rect 4509 17978 4565 17980
rect 4589 17978 4645 17980
rect 4669 17978 4725 17980
rect 4429 17926 4475 17978
rect 4475 17926 4485 17978
rect 4509 17926 4539 17978
rect 4539 17926 4551 17978
rect 4551 17926 4565 17978
rect 4589 17926 4603 17978
rect 4603 17926 4615 17978
rect 4615 17926 4645 17978
rect 4669 17926 4679 17978
rect 4679 17926 4725 17978
rect 4429 17924 4485 17926
rect 4509 17924 4565 17926
rect 4589 17924 4645 17926
rect 4669 17924 4725 17926
rect 4429 16890 4485 16892
rect 4509 16890 4565 16892
rect 4589 16890 4645 16892
rect 4669 16890 4725 16892
rect 4429 16838 4475 16890
rect 4475 16838 4485 16890
rect 4509 16838 4539 16890
rect 4539 16838 4551 16890
rect 4551 16838 4565 16890
rect 4589 16838 4603 16890
rect 4603 16838 4615 16890
rect 4615 16838 4645 16890
rect 4669 16838 4679 16890
rect 4679 16838 4725 16890
rect 4429 16836 4485 16838
rect 4509 16836 4565 16838
rect 4589 16836 4645 16838
rect 4669 16836 4725 16838
rect 4429 15802 4485 15804
rect 4509 15802 4565 15804
rect 4589 15802 4645 15804
rect 4669 15802 4725 15804
rect 4429 15750 4475 15802
rect 4475 15750 4485 15802
rect 4509 15750 4539 15802
rect 4539 15750 4551 15802
rect 4551 15750 4565 15802
rect 4589 15750 4603 15802
rect 4603 15750 4615 15802
rect 4615 15750 4645 15802
rect 4669 15750 4679 15802
rect 4679 15750 4725 15802
rect 4429 15748 4485 15750
rect 4509 15748 4565 15750
rect 4589 15748 4645 15750
rect 4669 15748 4725 15750
rect 4429 14714 4485 14716
rect 4509 14714 4565 14716
rect 4589 14714 4645 14716
rect 4669 14714 4725 14716
rect 4429 14662 4475 14714
rect 4475 14662 4485 14714
rect 4509 14662 4539 14714
rect 4539 14662 4551 14714
rect 4551 14662 4565 14714
rect 4589 14662 4603 14714
rect 4603 14662 4615 14714
rect 4615 14662 4645 14714
rect 4669 14662 4679 14714
rect 4679 14662 4725 14714
rect 4429 14660 4485 14662
rect 4509 14660 4565 14662
rect 4589 14660 4645 14662
rect 4669 14660 4725 14662
rect 4429 13626 4485 13628
rect 4509 13626 4565 13628
rect 4589 13626 4645 13628
rect 4669 13626 4725 13628
rect 4429 13574 4475 13626
rect 4475 13574 4485 13626
rect 4509 13574 4539 13626
rect 4539 13574 4551 13626
rect 4551 13574 4565 13626
rect 4589 13574 4603 13626
rect 4603 13574 4615 13626
rect 4615 13574 4645 13626
rect 4669 13574 4679 13626
rect 4679 13574 4725 13626
rect 4429 13572 4485 13574
rect 4509 13572 4565 13574
rect 4589 13572 4645 13574
rect 4669 13572 4725 13574
rect 4429 12538 4485 12540
rect 4509 12538 4565 12540
rect 4589 12538 4645 12540
rect 4669 12538 4725 12540
rect 4429 12486 4475 12538
rect 4475 12486 4485 12538
rect 4509 12486 4539 12538
rect 4539 12486 4551 12538
rect 4551 12486 4565 12538
rect 4589 12486 4603 12538
rect 4603 12486 4615 12538
rect 4615 12486 4645 12538
rect 4669 12486 4679 12538
rect 4679 12486 4725 12538
rect 4429 12484 4485 12486
rect 4509 12484 4565 12486
rect 4589 12484 4645 12486
rect 4669 12484 4725 12486
rect 7902 26138 7958 26140
rect 7982 26138 8038 26140
rect 8062 26138 8118 26140
rect 8142 26138 8198 26140
rect 7902 26086 7948 26138
rect 7948 26086 7958 26138
rect 7982 26086 8012 26138
rect 8012 26086 8024 26138
rect 8024 26086 8038 26138
rect 8062 26086 8076 26138
rect 8076 26086 8088 26138
rect 8088 26086 8118 26138
rect 8142 26086 8152 26138
rect 8152 26086 8198 26138
rect 7902 26084 7958 26086
rect 7982 26084 8038 26086
rect 8062 26084 8118 26086
rect 8142 26084 8198 26086
rect 7902 25050 7958 25052
rect 7982 25050 8038 25052
rect 8062 25050 8118 25052
rect 8142 25050 8198 25052
rect 7902 24998 7948 25050
rect 7948 24998 7958 25050
rect 7982 24998 8012 25050
rect 8012 24998 8024 25050
rect 8024 24998 8038 25050
rect 8062 24998 8076 25050
rect 8076 24998 8088 25050
rect 8088 24998 8118 25050
rect 8142 24998 8152 25050
rect 8152 24998 8198 25050
rect 7902 24996 7958 24998
rect 7982 24996 8038 24998
rect 8062 24996 8118 24998
rect 8142 24996 8198 24998
rect 4429 11450 4485 11452
rect 4509 11450 4565 11452
rect 4589 11450 4645 11452
rect 4669 11450 4725 11452
rect 4429 11398 4475 11450
rect 4475 11398 4485 11450
rect 4509 11398 4539 11450
rect 4539 11398 4551 11450
rect 4551 11398 4565 11450
rect 4589 11398 4603 11450
rect 4603 11398 4615 11450
rect 4615 11398 4645 11450
rect 4669 11398 4679 11450
rect 4679 11398 4725 11450
rect 4429 11396 4485 11398
rect 4509 11396 4565 11398
rect 4589 11396 4645 11398
rect 4669 11396 4725 11398
rect 4429 10362 4485 10364
rect 4509 10362 4565 10364
rect 4589 10362 4645 10364
rect 4669 10362 4725 10364
rect 4429 10310 4475 10362
rect 4475 10310 4485 10362
rect 4509 10310 4539 10362
rect 4539 10310 4551 10362
rect 4551 10310 4565 10362
rect 4589 10310 4603 10362
rect 4603 10310 4615 10362
rect 4615 10310 4645 10362
rect 4669 10310 4679 10362
rect 4679 10310 4725 10362
rect 4429 10308 4485 10310
rect 4509 10308 4565 10310
rect 4589 10308 4645 10310
rect 4669 10308 4725 10310
rect 4429 9274 4485 9276
rect 4509 9274 4565 9276
rect 4589 9274 4645 9276
rect 4669 9274 4725 9276
rect 4429 9222 4475 9274
rect 4475 9222 4485 9274
rect 4509 9222 4539 9274
rect 4539 9222 4551 9274
rect 4551 9222 4565 9274
rect 4589 9222 4603 9274
rect 4603 9222 4615 9274
rect 4615 9222 4645 9274
rect 4669 9222 4679 9274
rect 4679 9222 4725 9274
rect 4429 9220 4485 9222
rect 4509 9220 4565 9222
rect 4589 9220 4645 9222
rect 4669 9220 4725 9222
rect 4429 8186 4485 8188
rect 4509 8186 4565 8188
rect 4589 8186 4645 8188
rect 4669 8186 4725 8188
rect 4429 8134 4475 8186
rect 4475 8134 4485 8186
rect 4509 8134 4539 8186
rect 4539 8134 4551 8186
rect 4551 8134 4565 8186
rect 4589 8134 4603 8186
rect 4603 8134 4615 8186
rect 4615 8134 4645 8186
rect 4669 8134 4679 8186
rect 4679 8134 4725 8186
rect 4429 8132 4485 8134
rect 4509 8132 4565 8134
rect 4589 8132 4645 8134
rect 4669 8132 4725 8134
rect 4429 7098 4485 7100
rect 4509 7098 4565 7100
rect 4589 7098 4645 7100
rect 4669 7098 4725 7100
rect 4429 7046 4475 7098
rect 4475 7046 4485 7098
rect 4509 7046 4539 7098
rect 4539 7046 4551 7098
rect 4551 7046 4565 7098
rect 4589 7046 4603 7098
rect 4603 7046 4615 7098
rect 4615 7046 4645 7098
rect 4669 7046 4679 7098
rect 4679 7046 4725 7098
rect 4429 7044 4485 7046
rect 4509 7044 4565 7046
rect 4589 7044 4645 7046
rect 4669 7044 4725 7046
rect 4429 6010 4485 6012
rect 4509 6010 4565 6012
rect 4589 6010 4645 6012
rect 4669 6010 4725 6012
rect 4429 5958 4475 6010
rect 4475 5958 4485 6010
rect 4509 5958 4539 6010
rect 4539 5958 4551 6010
rect 4551 5958 4565 6010
rect 4589 5958 4603 6010
rect 4603 5958 4615 6010
rect 4615 5958 4645 6010
rect 4669 5958 4679 6010
rect 4679 5958 4725 6010
rect 4429 5956 4485 5958
rect 4509 5956 4565 5958
rect 4589 5956 4645 5958
rect 4669 5956 4725 5958
rect 7902 23962 7958 23964
rect 7982 23962 8038 23964
rect 8062 23962 8118 23964
rect 8142 23962 8198 23964
rect 7902 23910 7948 23962
rect 7948 23910 7958 23962
rect 7982 23910 8012 23962
rect 8012 23910 8024 23962
rect 8024 23910 8038 23962
rect 8062 23910 8076 23962
rect 8076 23910 8088 23962
rect 8088 23910 8118 23962
rect 8142 23910 8152 23962
rect 8152 23910 8198 23962
rect 7902 23908 7958 23910
rect 7982 23908 8038 23910
rect 8062 23908 8118 23910
rect 8142 23908 8198 23910
rect 7902 22874 7958 22876
rect 7982 22874 8038 22876
rect 8062 22874 8118 22876
rect 8142 22874 8198 22876
rect 7902 22822 7948 22874
rect 7948 22822 7958 22874
rect 7982 22822 8012 22874
rect 8012 22822 8024 22874
rect 8024 22822 8038 22874
rect 8062 22822 8076 22874
rect 8076 22822 8088 22874
rect 8088 22822 8118 22874
rect 8142 22822 8152 22874
rect 8152 22822 8198 22874
rect 7902 22820 7958 22822
rect 7982 22820 8038 22822
rect 8062 22820 8118 22822
rect 8142 22820 8198 22822
rect 7902 21786 7958 21788
rect 7982 21786 8038 21788
rect 8062 21786 8118 21788
rect 8142 21786 8198 21788
rect 7902 21734 7948 21786
rect 7948 21734 7958 21786
rect 7982 21734 8012 21786
rect 8012 21734 8024 21786
rect 8024 21734 8038 21786
rect 8062 21734 8076 21786
rect 8076 21734 8088 21786
rect 8088 21734 8118 21786
rect 8142 21734 8152 21786
rect 8152 21734 8198 21786
rect 7902 21732 7958 21734
rect 7982 21732 8038 21734
rect 8062 21732 8118 21734
rect 8142 21732 8198 21734
rect 7902 20698 7958 20700
rect 7982 20698 8038 20700
rect 8062 20698 8118 20700
rect 8142 20698 8198 20700
rect 7902 20646 7948 20698
rect 7948 20646 7958 20698
rect 7982 20646 8012 20698
rect 8012 20646 8024 20698
rect 8024 20646 8038 20698
rect 8062 20646 8076 20698
rect 8076 20646 8088 20698
rect 8088 20646 8118 20698
rect 8142 20646 8152 20698
rect 8152 20646 8198 20698
rect 7902 20644 7958 20646
rect 7982 20644 8038 20646
rect 8062 20644 8118 20646
rect 8142 20644 8198 20646
rect 7902 19610 7958 19612
rect 7982 19610 8038 19612
rect 8062 19610 8118 19612
rect 8142 19610 8198 19612
rect 7902 19558 7948 19610
rect 7948 19558 7958 19610
rect 7982 19558 8012 19610
rect 8012 19558 8024 19610
rect 8024 19558 8038 19610
rect 8062 19558 8076 19610
rect 8076 19558 8088 19610
rect 8088 19558 8118 19610
rect 8142 19558 8152 19610
rect 8152 19558 8198 19610
rect 7902 19556 7958 19558
rect 7982 19556 8038 19558
rect 8062 19556 8118 19558
rect 8142 19556 8198 19558
rect 7902 18522 7958 18524
rect 7982 18522 8038 18524
rect 8062 18522 8118 18524
rect 8142 18522 8198 18524
rect 7902 18470 7948 18522
rect 7948 18470 7958 18522
rect 7982 18470 8012 18522
rect 8012 18470 8024 18522
rect 8024 18470 8038 18522
rect 8062 18470 8076 18522
rect 8076 18470 8088 18522
rect 8088 18470 8118 18522
rect 8142 18470 8152 18522
rect 8152 18470 8198 18522
rect 7902 18468 7958 18470
rect 7982 18468 8038 18470
rect 8062 18468 8118 18470
rect 8142 18468 8198 18470
rect 7902 17434 7958 17436
rect 7982 17434 8038 17436
rect 8062 17434 8118 17436
rect 8142 17434 8198 17436
rect 7902 17382 7948 17434
rect 7948 17382 7958 17434
rect 7982 17382 8012 17434
rect 8012 17382 8024 17434
rect 8024 17382 8038 17434
rect 8062 17382 8076 17434
rect 8076 17382 8088 17434
rect 8088 17382 8118 17434
rect 8142 17382 8152 17434
rect 8152 17382 8198 17434
rect 7902 17380 7958 17382
rect 7982 17380 8038 17382
rect 8062 17380 8118 17382
rect 8142 17380 8198 17382
rect 7902 16346 7958 16348
rect 7982 16346 8038 16348
rect 8062 16346 8118 16348
rect 8142 16346 8198 16348
rect 7902 16294 7948 16346
rect 7948 16294 7958 16346
rect 7982 16294 8012 16346
rect 8012 16294 8024 16346
rect 8024 16294 8038 16346
rect 8062 16294 8076 16346
rect 8076 16294 8088 16346
rect 8088 16294 8118 16346
rect 8142 16294 8152 16346
rect 8152 16294 8198 16346
rect 7902 16292 7958 16294
rect 7982 16292 8038 16294
rect 8062 16292 8118 16294
rect 8142 16292 8198 16294
rect 11375 26682 11431 26684
rect 11455 26682 11511 26684
rect 11535 26682 11591 26684
rect 11615 26682 11671 26684
rect 11375 26630 11421 26682
rect 11421 26630 11431 26682
rect 11455 26630 11485 26682
rect 11485 26630 11497 26682
rect 11497 26630 11511 26682
rect 11535 26630 11549 26682
rect 11549 26630 11561 26682
rect 11561 26630 11591 26682
rect 11615 26630 11625 26682
rect 11625 26630 11671 26682
rect 11375 26628 11431 26630
rect 11455 26628 11511 26630
rect 11535 26628 11591 26630
rect 11615 26628 11671 26630
rect 11375 25594 11431 25596
rect 11455 25594 11511 25596
rect 11535 25594 11591 25596
rect 11615 25594 11671 25596
rect 11375 25542 11421 25594
rect 11421 25542 11431 25594
rect 11455 25542 11485 25594
rect 11485 25542 11497 25594
rect 11497 25542 11511 25594
rect 11535 25542 11549 25594
rect 11549 25542 11561 25594
rect 11561 25542 11591 25594
rect 11615 25542 11625 25594
rect 11625 25542 11671 25594
rect 11375 25540 11431 25542
rect 11455 25540 11511 25542
rect 11535 25540 11591 25542
rect 11615 25540 11671 25542
rect 11375 24506 11431 24508
rect 11455 24506 11511 24508
rect 11535 24506 11591 24508
rect 11615 24506 11671 24508
rect 11375 24454 11421 24506
rect 11421 24454 11431 24506
rect 11455 24454 11485 24506
rect 11485 24454 11497 24506
rect 11497 24454 11511 24506
rect 11535 24454 11549 24506
rect 11549 24454 11561 24506
rect 11561 24454 11591 24506
rect 11615 24454 11625 24506
rect 11625 24454 11671 24506
rect 11375 24452 11431 24454
rect 11455 24452 11511 24454
rect 11535 24452 11591 24454
rect 11615 24452 11671 24454
rect 11375 23418 11431 23420
rect 11455 23418 11511 23420
rect 11535 23418 11591 23420
rect 11615 23418 11671 23420
rect 11375 23366 11421 23418
rect 11421 23366 11431 23418
rect 11455 23366 11485 23418
rect 11485 23366 11497 23418
rect 11497 23366 11511 23418
rect 11535 23366 11549 23418
rect 11549 23366 11561 23418
rect 11561 23366 11591 23418
rect 11615 23366 11625 23418
rect 11625 23366 11671 23418
rect 11375 23364 11431 23366
rect 11455 23364 11511 23366
rect 11535 23364 11591 23366
rect 11615 23364 11671 23366
rect 11375 22330 11431 22332
rect 11455 22330 11511 22332
rect 11535 22330 11591 22332
rect 11615 22330 11671 22332
rect 11375 22278 11421 22330
rect 11421 22278 11431 22330
rect 11455 22278 11485 22330
rect 11485 22278 11497 22330
rect 11497 22278 11511 22330
rect 11535 22278 11549 22330
rect 11549 22278 11561 22330
rect 11561 22278 11591 22330
rect 11615 22278 11625 22330
rect 11625 22278 11671 22330
rect 11375 22276 11431 22278
rect 11455 22276 11511 22278
rect 11535 22276 11591 22278
rect 11615 22276 11671 22278
rect 11375 21242 11431 21244
rect 11455 21242 11511 21244
rect 11535 21242 11591 21244
rect 11615 21242 11671 21244
rect 11375 21190 11421 21242
rect 11421 21190 11431 21242
rect 11455 21190 11485 21242
rect 11485 21190 11497 21242
rect 11497 21190 11511 21242
rect 11535 21190 11549 21242
rect 11549 21190 11561 21242
rect 11561 21190 11591 21242
rect 11615 21190 11625 21242
rect 11625 21190 11671 21242
rect 11375 21188 11431 21190
rect 11455 21188 11511 21190
rect 11535 21188 11591 21190
rect 11615 21188 11671 21190
rect 11375 20154 11431 20156
rect 11455 20154 11511 20156
rect 11535 20154 11591 20156
rect 11615 20154 11671 20156
rect 11375 20102 11421 20154
rect 11421 20102 11431 20154
rect 11455 20102 11485 20154
rect 11485 20102 11497 20154
rect 11497 20102 11511 20154
rect 11535 20102 11549 20154
rect 11549 20102 11561 20154
rect 11561 20102 11591 20154
rect 11615 20102 11625 20154
rect 11625 20102 11671 20154
rect 11375 20100 11431 20102
rect 11455 20100 11511 20102
rect 11535 20100 11591 20102
rect 11615 20100 11671 20102
rect 11375 19066 11431 19068
rect 11455 19066 11511 19068
rect 11535 19066 11591 19068
rect 11615 19066 11671 19068
rect 11375 19014 11421 19066
rect 11421 19014 11431 19066
rect 11455 19014 11485 19066
rect 11485 19014 11497 19066
rect 11497 19014 11511 19066
rect 11535 19014 11549 19066
rect 11549 19014 11561 19066
rect 11561 19014 11591 19066
rect 11615 19014 11625 19066
rect 11625 19014 11671 19066
rect 11375 19012 11431 19014
rect 11455 19012 11511 19014
rect 11535 19012 11591 19014
rect 11615 19012 11671 19014
rect 11375 17978 11431 17980
rect 11455 17978 11511 17980
rect 11535 17978 11591 17980
rect 11615 17978 11671 17980
rect 11375 17926 11421 17978
rect 11421 17926 11431 17978
rect 11455 17926 11485 17978
rect 11485 17926 11497 17978
rect 11497 17926 11511 17978
rect 11535 17926 11549 17978
rect 11549 17926 11561 17978
rect 11561 17926 11591 17978
rect 11615 17926 11625 17978
rect 11625 17926 11671 17978
rect 11375 17924 11431 17926
rect 11455 17924 11511 17926
rect 11535 17924 11591 17926
rect 11615 17924 11671 17926
rect 11375 16890 11431 16892
rect 11455 16890 11511 16892
rect 11535 16890 11591 16892
rect 11615 16890 11671 16892
rect 11375 16838 11421 16890
rect 11421 16838 11431 16890
rect 11455 16838 11485 16890
rect 11485 16838 11497 16890
rect 11497 16838 11511 16890
rect 11535 16838 11549 16890
rect 11549 16838 11561 16890
rect 11561 16838 11591 16890
rect 11615 16838 11625 16890
rect 11625 16838 11671 16890
rect 11375 16836 11431 16838
rect 11455 16836 11511 16838
rect 11535 16836 11591 16838
rect 11615 16836 11671 16838
rect 11375 15802 11431 15804
rect 11455 15802 11511 15804
rect 11535 15802 11591 15804
rect 11615 15802 11671 15804
rect 11375 15750 11421 15802
rect 11421 15750 11431 15802
rect 11455 15750 11485 15802
rect 11485 15750 11497 15802
rect 11497 15750 11511 15802
rect 11535 15750 11549 15802
rect 11549 15750 11561 15802
rect 11561 15750 11591 15802
rect 11615 15750 11625 15802
rect 11625 15750 11671 15802
rect 11375 15748 11431 15750
rect 11455 15748 11511 15750
rect 11535 15748 11591 15750
rect 11615 15748 11671 15750
rect 7902 15258 7958 15260
rect 7982 15258 8038 15260
rect 8062 15258 8118 15260
rect 8142 15258 8198 15260
rect 7902 15206 7948 15258
rect 7948 15206 7958 15258
rect 7982 15206 8012 15258
rect 8012 15206 8024 15258
rect 8024 15206 8038 15258
rect 8062 15206 8076 15258
rect 8076 15206 8088 15258
rect 8088 15206 8118 15258
rect 8142 15206 8152 15258
rect 8152 15206 8198 15258
rect 7902 15204 7958 15206
rect 7982 15204 8038 15206
rect 8062 15204 8118 15206
rect 8142 15204 8198 15206
rect 7902 14170 7958 14172
rect 7982 14170 8038 14172
rect 8062 14170 8118 14172
rect 8142 14170 8198 14172
rect 7902 14118 7948 14170
rect 7948 14118 7958 14170
rect 7982 14118 8012 14170
rect 8012 14118 8024 14170
rect 8024 14118 8038 14170
rect 8062 14118 8076 14170
rect 8076 14118 8088 14170
rect 8088 14118 8118 14170
rect 8142 14118 8152 14170
rect 8152 14118 8198 14170
rect 7902 14116 7958 14118
rect 7982 14116 8038 14118
rect 8062 14116 8118 14118
rect 8142 14116 8198 14118
rect 7902 13082 7958 13084
rect 7982 13082 8038 13084
rect 8062 13082 8118 13084
rect 8142 13082 8198 13084
rect 7902 13030 7948 13082
rect 7948 13030 7958 13082
rect 7982 13030 8012 13082
rect 8012 13030 8024 13082
rect 8024 13030 8038 13082
rect 8062 13030 8076 13082
rect 8076 13030 8088 13082
rect 8088 13030 8118 13082
rect 8142 13030 8152 13082
rect 8152 13030 8198 13082
rect 7902 13028 7958 13030
rect 7982 13028 8038 13030
rect 8062 13028 8118 13030
rect 8142 13028 8198 13030
rect 7902 11994 7958 11996
rect 7982 11994 8038 11996
rect 8062 11994 8118 11996
rect 8142 11994 8198 11996
rect 7902 11942 7948 11994
rect 7948 11942 7958 11994
rect 7982 11942 8012 11994
rect 8012 11942 8024 11994
rect 8024 11942 8038 11994
rect 8062 11942 8076 11994
rect 8076 11942 8088 11994
rect 8088 11942 8118 11994
rect 8142 11942 8152 11994
rect 8152 11942 8198 11994
rect 7902 11940 7958 11942
rect 7982 11940 8038 11942
rect 8062 11940 8118 11942
rect 8142 11940 8198 11942
rect 7902 10906 7958 10908
rect 7982 10906 8038 10908
rect 8062 10906 8118 10908
rect 8142 10906 8198 10908
rect 7902 10854 7948 10906
rect 7948 10854 7958 10906
rect 7982 10854 8012 10906
rect 8012 10854 8024 10906
rect 8024 10854 8038 10906
rect 8062 10854 8076 10906
rect 8076 10854 8088 10906
rect 8088 10854 8118 10906
rect 8142 10854 8152 10906
rect 8152 10854 8198 10906
rect 7902 10852 7958 10854
rect 7982 10852 8038 10854
rect 8062 10852 8118 10854
rect 8142 10852 8198 10854
rect 7902 9818 7958 9820
rect 7982 9818 8038 9820
rect 8062 9818 8118 9820
rect 8142 9818 8198 9820
rect 7902 9766 7948 9818
rect 7948 9766 7958 9818
rect 7982 9766 8012 9818
rect 8012 9766 8024 9818
rect 8024 9766 8038 9818
rect 8062 9766 8076 9818
rect 8076 9766 8088 9818
rect 8088 9766 8118 9818
rect 8142 9766 8152 9818
rect 8152 9766 8198 9818
rect 7902 9764 7958 9766
rect 7982 9764 8038 9766
rect 8062 9764 8118 9766
rect 8142 9764 8198 9766
rect 4429 4922 4485 4924
rect 4509 4922 4565 4924
rect 4589 4922 4645 4924
rect 4669 4922 4725 4924
rect 4429 4870 4475 4922
rect 4475 4870 4485 4922
rect 4509 4870 4539 4922
rect 4539 4870 4551 4922
rect 4551 4870 4565 4922
rect 4589 4870 4603 4922
rect 4603 4870 4615 4922
rect 4615 4870 4645 4922
rect 4669 4870 4679 4922
rect 4679 4870 4725 4922
rect 4429 4868 4485 4870
rect 4509 4868 4565 4870
rect 4589 4868 4645 4870
rect 4669 4868 4725 4870
rect 4429 3834 4485 3836
rect 4509 3834 4565 3836
rect 4589 3834 4645 3836
rect 4669 3834 4725 3836
rect 4429 3782 4475 3834
rect 4475 3782 4485 3834
rect 4509 3782 4539 3834
rect 4539 3782 4551 3834
rect 4551 3782 4565 3834
rect 4589 3782 4603 3834
rect 4603 3782 4615 3834
rect 4615 3782 4645 3834
rect 4669 3782 4679 3834
rect 4679 3782 4725 3834
rect 4429 3780 4485 3782
rect 4509 3780 4565 3782
rect 4589 3780 4645 3782
rect 4669 3780 4725 3782
rect 7902 8730 7958 8732
rect 7982 8730 8038 8732
rect 8062 8730 8118 8732
rect 8142 8730 8198 8732
rect 7902 8678 7948 8730
rect 7948 8678 7958 8730
rect 7982 8678 8012 8730
rect 8012 8678 8024 8730
rect 8024 8678 8038 8730
rect 8062 8678 8076 8730
rect 8076 8678 8088 8730
rect 8088 8678 8118 8730
rect 8142 8678 8152 8730
rect 8152 8678 8198 8730
rect 7902 8676 7958 8678
rect 7982 8676 8038 8678
rect 8062 8676 8118 8678
rect 8142 8676 8198 8678
rect 7902 7642 7958 7644
rect 7982 7642 8038 7644
rect 8062 7642 8118 7644
rect 8142 7642 8198 7644
rect 7902 7590 7948 7642
rect 7948 7590 7958 7642
rect 7982 7590 8012 7642
rect 8012 7590 8024 7642
rect 8024 7590 8038 7642
rect 8062 7590 8076 7642
rect 8076 7590 8088 7642
rect 8088 7590 8118 7642
rect 8142 7590 8152 7642
rect 8152 7590 8198 7642
rect 7902 7588 7958 7590
rect 7982 7588 8038 7590
rect 8062 7588 8118 7590
rect 8142 7588 8198 7590
rect 7902 6554 7958 6556
rect 7982 6554 8038 6556
rect 8062 6554 8118 6556
rect 8142 6554 8198 6556
rect 7902 6502 7948 6554
rect 7948 6502 7958 6554
rect 7982 6502 8012 6554
rect 8012 6502 8024 6554
rect 8024 6502 8038 6554
rect 8062 6502 8076 6554
rect 8076 6502 8088 6554
rect 8088 6502 8118 6554
rect 8142 6502 8152 6554
rect 8152 6502 8198 6554
rect 7902 6500 7958 6502
rect 7982 6500 8038 6502
rect 8062 6500 8118 6502
rect 8142 6500 8198 6502
rect 7902 5466 7958 5468
rect 7982 5466 8038 5468
rect 8062 5466 8118 5468
rect 8142 5466 8198 5468
rect 7902 5414 7948 5466
rect 7948 5414 7958 5466
rect 7982 5414 8012 5466
rect 8012 5414 8024 5466
rect 8024 5414 8038 5466
rect 8062 5414 8076 5466
rect 8076 5414 8088 5466
rect 8088 5414 8118 5466
rect 8142 5414 8152 5466
rect 8152 5414 8198 5466
rect 7902 5412 7958 5414
rect 7982 5412 8038 5414
rect 8062 5412 8118 5414
rect 8142 5412 8198 5414
rect 4429 2746 4485 2748
rect 4509 2746 4565 2748
rect 4589 2746 4645 2748
rect 4669 2746 4725 2748
rect 4429 2694 4475 2746
rect 4475 2694 4485 2746
rect 4509 2694 4539 2746
rect 4539 2694 4551 2746
rect 4551 2694 4565 2746
rect 4589 2694 4603 2746
rect 4603 2694 4615 2746
rect 4615 2694 4645 2746
rect 4669 2694 4679 2746
rect 4679 2694 4725 2746
rect 4429 2692 4485 2694
rect 4509 2692 4565 2694
rect 4589 2692 4645 2694
rect 4669 2692 4725 2694
rect 7902 4378 7958 4380
rect 7982 4378 8038 4380
rect 8062 4378 8118 4380
rect 8142 4378 8198 4380
rect 7902 4326 7948 4378
rect 7948 4326 7958 4378
rect 7982 4326 8012 4378
rect 8012 4326 8024 4378
rect 8024 4326 8038 4378
rect 8062 4326 8076 4378
rect 8076 4326 8088 4378
rect 8088 4326 8118 4378
rect 8142 4326 8152 4378
rect 8152 4326 8198 4378
rect 7902 4324 7958 4326
rect 7982 4324 8038 4326
rect 8062 4324 8118 4326
rect 8142 4324 8198 4326
rect 7902 3290 7958 3292
rect 7982 3290 8038 3292
rect 8062 3290 8118 3292
rect 8142 3290 8198 3292
rect 7902 3238 7948 3290
rect 7948 3238 7958 3290
rect 7982 3238 8012 3290
rect 8012 3238 8024 3290
rect 8024 3238 8038 3290
rect 8062 3238 8076 3290
rect 8076 3238 8088 3290
rect 8088 3238 8118 3290
rect 8142 3238 8152 3290
rect 8152 3238 8198 3290
rect 7902 3236 7958 3238
rect 7982 3236 8038 3238
rect 8062 3236 8118 3238
rect 8142 3236 8198 3238
rect 11375 14714 11431 14716
rect 11455 14714 11511 14716
rect 11535 14714 11591 14716
rect 11615 14714 11671 14716
rect 11375 14662 11421 14714
rect 11421 14662 11431 14714
rect 11455 14662 11485 14714
rect 11485 14662 11497 14714
rect 11497 14662 11511 14714
rect 11535 14662 11549 14714
rect 11549 14662 11561 14714
rect 11561 14662 11591 14714
rect 11615 14662 11625 14714
rect 11625 14662 11671 14714
rect 11375 14660 11431 14662
rect 11455 14660 11511 14662
rect 11535 14660 11591 14662
rect 11615 14660 11671 14662
rect 11375 13626 11431 13628
rect 11455 13626 11511 13628
rect 11535 13626 11591 13628
rect 11615 13626 11671 13628
rect 11375 13574 11421 13626
rect 11421 13574 11431 13626
rect 11455 13574 11485 13626
rect 11485 13574 11497 13626
rect 11497 13574 11511 13626
rect 11535 13574 11549 13626
rect 11549 13574 11561 13626
rect 11561 13574 11591 13626
rect 11615 13574 11625 13626
rect 11625 13574 11671 13626
rect 11375 13572 11431 13574
rect 11455 13572 11511 13574
rect 11535 13572 11591 13574
rect 11615 13572 11671 13574
rect 11375 12538 11431 12540
rect 11455 12538 11511 12540
rect 11535 12538 11591 12540
rect 11615 12538 11671 12540
rect 11375 12486 11421 12538
rect 11421 12486 11431 12538
rect 11455 12486 11485 12538
rect 11485 12486 11497 12538
rect 11497 12486 11511 12538
rect 11535 12486 11549 12538
rect 11549 12486 11561 12538
rect 11561 12486 11591 12538
rect 11615 12486 11625 12538
rect 11625 12486 11671 12538
rect 11375 12484 11431 12486
rect 11455 12484 11511 12486
rect 11535 12484 11591 12486
rect 11615 12484 11671 12486
rect 11375 11450 11431 11452
rect 11455 11450 11511 11452
rect 11535 11450 11591 11452
rect 11615 11450 11671 11452
rect 11375 11398 11421 11450
rect 11421 11398 11431 11450
rect 11455 11398 11485 11450
rect 11485 11398 11497 11450
rect 11497 11398 11511 11450
rect 11535 11398 11549 11450
rect 11549 11398 11561 11450
rect 11561 11398 11591 11450
rect 11615 11398 11625 11450
rect 11625 11398 11671 11450
rect 11375 11396 11431 11398
rect 11455 11396 11511 11398
rect 11535 11396 11591 11398
rect 11615 11396 11671 11398
rect 11375 10362 11431 10364
rect 11455 10362 11511 10364
rect 11535 10362 11591 10364
rect 11615 10362 11671 10364
rect 11375 10310 11421 10362
rect 11421 10310 11431 10362
rect 11455 10310 11485 10362
rect 11485 10310 11497 10362
rect 11497 10310 11511 10362
rect 11535 10310 11549 10362
rect 11549 10310 11561 10362
rect 11561 10310 11591 10362
rect 11615 10310 11625 10362
rect 11625 10310 11671 10362
rect 11375 10308 11431 10310
rect 11455 10308 11511 10310
rect 11535 10308 11591 10310
rect 11615 10308 11671 10310
rect 11375 9274 11431 9276
rect 11455 9274 11511 9276
rect 11535 9274 11591 9276
rect 11615 9274 11671 9276
rect 11375 9222 11421 9274
rect 11421 9222 11431 9274
rect 11455 9222 11485 9274
rect 11485 9222 11497 9274
rect 11497 9222 11511 9274
rect 11535 9222 11549 9274
rect 11549 9222 11561 9274
rect 11561 9222 11591 9274
rect 11615 9222 11625 9274
rect 11625 9222 11671 9274
rect 11375 9220 11431 9222
rect 11455 9220 11511 9222
rect 11535 9220 11591 9222
rect 11615 9220 11671 9222
rect 14848 27226 14904 27228
rect 14928 27226 14984 27228
rect 15008 27226 15064 27228
rect 15088 27226 15144 27228
rect 14848 27174 14894 27226
rect 14894 27174 14904 27226
rect 14928 27174 14958 27226
rect 14958 27174 14970 27226
rect 14970 27174 14984 27226
rect 15008 27174 15022 27226
rect 15022 27174 15034 27226
rect 15034 27174 15064 27226
rect 15088 27174 15098 27226
rect 15098 27174 15144 27226
rect 14848 27172 14904 27174
rect 14928 27172 14984 27174
rect 15008 27172 15064 27174
rect 15088 27172 15144 27174
rect 14848 26138 14904 26140
rect 14928 26138 14984 26140
rect 15008 26138 15064 26140
rect 15088 26138 15144 26140
rect 14848 26086 14894 26138
rect 14894 26086 14904 26138
rect 14928 26086 14958 26138
rect 14958 26086 14970 26138
rect 14970 26086 14984 26138
rect 15008 26086 15022 26138
rect 15022 26086 15034 26138
rect 15034 26086 15064 26138
rect 15088 26086 15098 26138
rect 15098 26086 15144 26138
rect 14848 26084 14904 26086
rect 14928 26084 14984 26086
rect 15008 26084 15064 26086
rect 15088 26084 15144 26086
rect 14848 25050 14904 25052
rect 14928 25050 14984 25052
rect 15008 25050 15064 25052
rect 15088 25050 15144 25052
rect 14848 24998 14894 25050
rect 14894 24998 14904 25050
rect 14928 24998 14958 25050
rect 14958 24998 14970 25050
rect 14970 24998 14984 25050
rect 15008 24998 15022 25050
rect 15022 24998 15034 25050
rect 15034 24998 15064 25050
rect 15088 24998 15098 25050
rect 15098 24998 15144 25050
rect 14848 24996 14904 24998
rect 14928 24996 14984 24998
rect 15008 24996 15064 24998
rect 15088 24996 15144 24998
rect 14848 23962 14904 23964
rect 14928 23962 14984 23964
rect 15008 23962 15064 23964
rect 15088 23962 15144 23964
rect 14848 23910 14894 23962
rect 14894 23910 14904 23962
rect 14928 23910 14958 23962
rect 14958 23910 14970 23962
rect 14970 23910 14984 23962
rect 15008 23910 15022 23962
rect 15022 23910 15034 23962
rect 15034 23910 15064 23962
rect 15088 23910 15098 23962
rect 15098 23910 15144 23962
rect 14848 23908 14904 23910
rect 14928 23908 14984 23910
rect 15008 23908 15064 23910
rect 15088 23908 15144 23910
rect 14848 22874 14904 22876
rect 14928 22874 14984 22876
rect 15008 22874 15064 22876
rect 15088 22874 15144 22876
rect 14848 22822 14894 22874
rect 14894 22822 14904 22874
rect 14928 22822 14958 22874
rect 14958 22822 14970 22874
rect 14970 22822 14984 22874
rect 15008 22822 15022 22874
rect 15022 22822 15034 22874
rect 15034 22822 15064 22874
rect 15088 22822 15098 22874
rect 15098 22822 15144 22874
rect 14848 22820 14904 22822
rect 14928 22820 14984 22822
rect 15008 22820 15064 22822
rect 15088 22820 15144 22822
rect 14848 21786 14904 21788
rect 14928 21786 14984 21788
rect 15008 21786 15064 21788
rect 15088 21786 15144 21788
rect 14848 21734 14894 21786
rect 14894 21734 14904 21786
rect 14928 21734 14958 21786
rect 14958 21734 14970 21786
rect 14970 21734 14984 21786
rect 15008 21734 15022 21786
rect 15022 21734 15034 21786
rect 15034 21734 15064 21786
rect 15088 21734 15098 21786
rect 15098 21734 15144 21786
rect 14848 21732 14904 21734
rect 14928 21732 14984 21734
rect 15008 21732 15064 21734
rect 15088 21732 15144 21734
rect 11375 8186 11431 8188
rect 11455 8186 11511 8188
rect 11535 8186 11591 8188
rect 11615 8186 11671 8188
rect 11375 8134 11421 8186
rect 11421 8134 11431 8186
rect 11455 8134 11485 8186
rect 11485 8134 11497 8186
rect 11497 8134 11511 8186
rect 11535 8134 11549 8186
rect 11549 8134 11561 8186
rect 11561 8134 11591 8186
rect 11615 8134 11625 8186
rect 11625 8134 11671 8186
rect 11375 8132 11431 8134
rect 11455 8132 11511 8134
rect 11535 8132 11591 8134
rect 11615 8132 11671 8134
rect 14848 20698 14904 20700
rect 14928 20698 14984 20700
rect 15008 20698 15064 20700
rect 15088 20698 15144 20700
rect 14848 20646 14894 20698
rect 14894 20646 14904 20698
rect 14928 20646 14958 20698
rect 14958 20646 14970 20698
rect 14970 20646 14984 20698
rect 15008 20646 15022 20698
rect 15022 20646 15034 20698
rect 15034 20646 15064 20698
rect 15088 20646 15098 20698
rect 15098 20646 15144 20698
rect 14848 20644 14904 20646
rect 14928 20644 14984 20646
rect 15008 20644 15064 20646
rect 15088 20644 15144 20646
rect 14848 19610 14904 19612
rect 14928 19610 14984 19612
rect 15008 19610 15064 19612
rect 15088 19610 15144 19612
rect 14848 19558 14894 19610
rect 14894 19558 14904 19610
rect 14928 19558 14958 19610
rect 14958 19558 14970 19610
rect 14970 19558 14984 19610
rect 15008 19558 15022 19610
rect 15022 19558 15034 19610
rect 15034 19558 15064 19610
rect 15088 19558 15098 19610
rect 15098 19558 15144 19610
rect 14848 19556 14904 19558
rect 14928 19556 14984 19558
rect 15008 19556 15064 19558
rect 15088 19556 15144 19558
rect 14848 18522 14904 18524
rect 14928 18522 14984 18524
rect 15008 18522 15064 18524
rect 15088 18522 15144 18524
rect 14848 18470 14894 18522
rect 14894 18470 14904 18522
rect 14928 18470 14958 18522
rect 14958 18470 14970 18522
rect 14970 18470 14984 18522
rect 15008 18470 15022 18522
rect 15022 18470 15034 18522
rect 15034 18470 15064 18522
rect 15088 18470 15098 18522
rect 15098 18470 15144 18522
rect 14848 18468 14904 18470
rect 14928 18468 14984 18470
rect 15008 18468 15064 18470
rect 15088 18468 15144 18470
rect 14848 17434 14904 17436
rect 14928 17434 14984 17436
rect 15008 17434 15064 17436
rect 15088 17434 15144 17436
rect 14848 17382 14894 17434
rect 14894 17382 14904 17434
rect 14928 17382 14958 17434
rect 14958 17382 14970 17434
rect 14970 17382 14984 17434
rect 15008 17382 15022 17434
rect 15022 17382 15034 17434
rect 15034 17382 15064 17434
rect 15088 17382 15098 17434
rect 15098 17382 15144 17434
rect 14848 17380 14904 17382
rect 14928 17380 14984 17382
rect 15008 17380 15064 17382
rect 15088 17380 15144 17382
rect 14848 16346 14904 16348
rect 14928 16346 14984 16348
rect 15008 16346 15064 16348
rect 15088 16346 15144 16348
rect 14848 16294 14894 16346
rect 14894 16294 14904 16346
rect 14928 16294 14958 16346
rect 14958 16294 14970 16346
rect 14970 16294 14984 16346
rect 15008 16294 15022 16346
rect 15022 16294 15034 16346
rect 15034 16294 15064 16346
rect 15088 16294 15098 16346
rect 15098 16294 15144 16346
rect 14848 16292 14904 16294
rect 14928 16292 14984 16294
rect 15008 16292 15064 16294
rect 15088 16292 15144 16294
rect 27526 27784 27582 27840
rect 25267 27770 25323 27772
rect 25347 27770 25403 27772
rect 25427 27770 25483 27772
rect 25507 27770 25563 27772
rect 25267 27718 25313 27770
rect 25313 27718 25323 27770
rect 25347 27718 25377 27770
rect 25377 27718 25389 27770
rect 25389 27718 25403 27770
rect 25427 27718 25441 27770
rect 25441 27718 25453 27770
rect 25453 27718 25483 27770
rect 25507 27718 25517 27770
rect 25517 27718 25563 27770
rect 25267 27716 25323 27718
rect 25347 27716 25403 27718
rect 25427 27716 25483 27718
rect 25507 27716 25563 27718
rect 18321 26682 18377 26684
rect 18401 26682 18457 26684
rect 18481 26682 18537 26684
rect 18561 26682 18617 26684
rect 18321 26630 18367 26682
rect 18367 26630 18377 26682
rect 18401 26630 18431 26682
rect 18431 26630 18443 26682
rect 18443 26630 18457 26682
rect 18481 26630 18495 26682
rect 18495 26630 18507 26682
rect 18507 26630 18537 26682
rect 18561 26630 18571 26682
rect 18571 26630 18617 26682
rect 18321 26628 18377 26630
rect 18401 26628 18457 26630
rect 18481 26628 18537 26630
rect 18561 26628 18617 26630
rect 18321 25594 18377 25596
rect 18401 25594 18457 25596
rect 18481 25594 18537 25596
rect 18561 25594 18617 25596
rect 18321 25542 18367 25594
rect 18367 25542 18377 25594
rect 18401 25542 18431 25594
rect 18431 25542 18443 25594
rect 18443 25542 18457 25594
rect 18481 25542 18495 25594
rect 18495 25542 18507 25594
rect 18507 25542 18537 25594
rect 18561 25542 18571 25594
rect 18571 25542 18617 25594
rect 18321 25540 18377 25542
rect 18401 25540 18457 25542
rect 18481 25540 18537 25542
rect 18561 25540 18617 25542
rect 18321 24506 18377 24508
rect 18401 24506 18457 24508
rect 18481 24506 18537 24508
rect 18561 24506 18617 24508
rect 18321 24454 18367 24506
rect 18367 24454 18377 24506
rect 18401 24454 18431 24506
rect 18431 24454 18443 24506
rect 18443 24454 18457 24506
rect 18481 24454 18495 24506
rect 18495 24454 18507 24506
rect 18507 24454 18537 24506
rect 18561 24454 18571 24506
rect 18571 24454 18617 24506
rect 18321 24452 18377 24454
rect 18401 24452 18457 24454
rect 18481 24452 18537 24454
rect 18561 24452 18617 24454
rect 18321 23418 18377 23420
rect 18401 23418 18457 23420
rect 18481 23418 18537 23420
rect 18561 23418 18617 23420
rect 18321 23366 18367 23418
rect 18367 23366 18377 23418
rect 18401 23366 18431 23418
rect 18431 23366 18443 23418
rect 18443 23366 18457 23418
rect 18481 23366 18495 23418
rect 18495 23366 18507 23418
rect 18507 23366 18537 23418
rect 18561 23366 18571 23418
rect 18571 23366 18617 23418
rect 18321 23364 18377 23366
rect 18401 23364 18457 23366
rect 18481 23364 18537 23366
rect 18561 23364 18617 23366
rect 14848 15258 14904 15260
rect 14928 15258 14984 15260
rect 15008 15258 15064 15260
rect 15088 15258 15144 15260
rect 14848 15206 14894 15258
rect 14894 15206 14904 15258
rect 14928 15206 14958 15258
rect 14958 15206 14970 15258
rect 14970 15206 14984 15258
rect 15008 15206 15022 15258
rect 15022 15206 15034 15258
rect 15034 15206 15064 15258
rect 15088 15206 15098 15258
rect 15098 15206 15144 15258
rect 14848 15204 14904 15206
rect 14928 15204 14984 15206
rect 15008 15204 15064 15206
rect 15088 15204 15144 15206
rect 14848 14170 14904 14172
rect 14928 14170 14984 14172
rect 15008 14170 15064 14172
rect 15088 14170 15144 14172
rect 14848 14118 14894 14170
rect 14894 14118 14904 14170
rect 14928 14118 14958 14170
rect 14958 14118 14970 14170
rect 14970 14118 14984 14170
rect 15008 14118 15022 14170
rect 15022 14118 15034 14170
rect 15034 14118 15064 14170
rect 15088 14118 15098 14170
rect 15098 14118 15144 14170
rect 14848 14116 14904 14118
rect 14928 14116 14984 14118
rect 15008 14116 15064 14118
rect 15088 14116 15144 14118
rect 18321 22330 18377 22332
rect 18401 22330 18457 22332
rect 18481 22330 18537 22332
rect 18561 22330 18617 22332
rect 18321 22278 18367 22330
rect 18367 22278 18377 22330
rect 18401 22278 18431 22330
rect 18431 22278 18443 22330
rect 18443 22278 18457 22330
rect 18481 22278 18495 22330
rect 18495 22278 18507 22330
rect 18507 22278 18537 22330
rect 18561 22278 18571 22330
rect 18571 22278 18617 22330
rect 18321 22276 18377 22278
rect 18401 22276 18457 22278
rect 18481 22276 18537 22278
rect 18561 22276 18617 22278
rect 21794 27226 21850 27228
rect 21874 27226 21930 27228
rect 21954 27226 22010 27228
rect 22034 27226 22090 27228
rect 21794 27174 21840 27226
rect 21840 27174 21850 27226
rect 21874 27174 21904 27226
rect 21904 27174 21916 27226
rect 21916 27174 21930 27226
rect 21954 27174 21968 27226
rect 21968 27174 21980 27226
rect 21980 27174 22010 27226
rect 22034 27174 22044 27226
rect 22044 27174 22090 27226
rect 21794 27172 21850 27174
rect 21874 27172 21930 27174
rect 21954 27172 22010 27174
rect 22034 27172 22090 27174
rect 21794 26138 21850 26140
rect 21874 26138 21930 26140
rect 21954 26138 22010 26140
rect 22034 26138 22090 26140
rect 21794 26086 21840 26138
rect 21840 26086 21850 26138
rect 21874 26086 21904 26138
rect 21904 26086 21916 26138
rect 21916 26086 21930 26138
rect 21954 26086 21968 26138
rect 21968 26086 21980 26138
rect 21980 26086 22010 26138
rect 22034 26086 22044 26138
rect 22044 26086 22090 26138
rect 21794 26084 21850 26086
rect 21874 26084 21930 26086
rect 21954 26084 22010 26086
rect 22034 26084 22090 26086
rect 21794 25050 21850 25052
rect 21874 25050 21930 25052
rect 21954 25050 22010 25052
rect 22034 25050 22090 25052
rect 21794 24998 21840 25050
rect 21840 24998 21850 25050
rect 21874 24998 21904 25050
rect 21904 24998 21916 25050
rect 21916 24998 21930 25050
rect 21954 24998 21968 25050
rect 21968 24998 21980 25050
rect 21980 24998 22010 25050
rect 22034 24998 22044 25050
rect 22044 24998 22090 25050
rect 21794 24996 21850 24998
rect 21874 24996 21930 24998
rect 21954 24996 22010 24998
rect 22034 24996 22090 24998
rect 21794 23962 21850 23964
rect 21874 23962 21930 23964
rect 21954 23962 22010 23964
rect 22034 23962 22090 23964
rect 21794 23910 21840 23962
rect 21840 23910 21850 23962
rect 21874 23910 21904 23962
rect 21904 23910 21916 23962
rect 21916 23910 21930 23962
rect 21954 23910 21968 23962
rect 21968 23910 21980 23962
rect 21980 23910 22010 23962
rect 22034 23910 22044 23962
rect 22044 23910 22090 23962
rect 21794 23908 21850 23910
rect 21874 23908 21930 23910
rect 21954 23908 22010 23910
rect 22034 23908 22090 23910
rect 18321 21242 18377 21244
rect 18401 21242 18457 21244
rect 18481 21242 18537 21244
rect 18561 21242 18617 21244
rect 18321 21190 18367 21242
rect 18367 21190 18377 21242
rect 18401 21190 18431 21242
rect 18431 21190 18443 21242
rect 18443 21190 18457 21242
rect 18481 21190 18495 21242
rect 18495 21190 18507 21242
rect 18507 21190 18537 21242
rect 18561 21190 18571 21242
rect 18571 21190 18617 21242
rect 18321 21188 18377 21190
rect 18401 21188 18457 21190
rect 18481 21188 18537 21190
rect 18561 21188 18617 21190
rect 18321 20154 18377 20156
rect 18401 20154 18457 20156
rect 18481 20154 18537 20156
rect 18561 20154 18617 20156
rect 18321 20102 18367 20154
rect 18367 20102 18377 20154
rect 18401 20102 18431 20154
rect 18431 20102 18443 20154
rect 18443 20102 18457 20154
rect 18481 20102 18495 20154
rect 18495 20102 18507 20154
rect 18507 20102 18537 20154
rect 18561 20102 18571 20154
rect 18571 20102 18617 20154
rect 18321 20100 18377 20102
rect 18401 20100 18457 20102
rect 18481 20100 18537 20102
rect 18561 20100 18617 20102
rect 14848 13082 14904 13084
rect 14928 13082 14984 13084
rect 15008 13082 15064 13084
rect 15088 13082 15144 13084
rect 14848 13030 14894 13082
rect 14894 13030 14904 13082
rect 14928 13030 14958 13082
rect 14958 13030 14970 13082
rect 14970 13030 14984 13082
rect 15008 13030 15022 13082
rect 15022 13030 15034 13082
rect 15034 13030 15064 13082
rect 15088 13030 15098 13082
rect 15098 13030 15144 13082
rect 14848 13028 14904 13030
rect 14928 13028 14984 13030
rect 15008 13028 15064 13030
rect 15088 13028 15144 13030
rect 11375 7098 11431 7100
rect 11455 7098 11511 7100
rect 11535 7098 11591 7100
rect 11615 7098 11671 7100
rect 11375 7046 11421 7098
rect 11421 7046 11431 7098
rect 11455 7046 11485 7098
rect 11485 7046 11497 7098
rect 11497 7046 11511 7098
rect 11535 7046 11549 7098
rect 11549 7046 11561 7098
rect 11561 7046 11591 7098
rect 11615 7046 11625 7098
rect 11625 7046 11671 7098
rect 11375 7044 11431 7046
rect 11455 7044 11511 7046
rect 11535 7044 11591 7046
rect 11615 7044 11671 7046
rect 11375 6010 11431 6012
rect 11455 6010 11511 6012
rect 11535 6010 11591 6012
rect 11615 6010 11671 6012
rect 11375 5958 11421 6010
rect 11421 5958 11431 6010
rect 11455 5958 11485 6010
rect 11485 5958 11497 6010
rect 11497 5958 11511 6010
rect 11535 5958 11549 6010
rect 11549 5958 11561 6010
rect 11561 5958 11591 6010
rect 11615 5958 11625 6010
rect 11625 5958 11671 6010
rect 11375 5956 11431 5958
rect 11455 5956 11511 5958
rect 11535 5956 11591 5958
rect 11615 5956 11671 5958
rect 11375 4922 11431 4924
rect 11455 4922 11511 4924
rect 11535 4922 11591 4924
rect 11615 4922 11671 4924
rect 11375 4870 11421 4922
rect 11421 4870 11431 4922
rect 11455 4870 11485 4922
rect 11485 4870 11497 4922
rect 11497 4870 11511 4922
rect 11535 4870 11549 4922
rect 11549 4870 11561 4922
rect 11561 4870 11591 4922
rect 11615 4870 11625 4922
rect 11625 4870 11671 4922
rect 11375 4868 11431 4870
rect 11455 4868 11511 4870
rect 11535 4868 11591 4870
rect 11615 4868 11671 4870
rect 11375 3834 11431 3836
rect 11455 3834 11511 3836
rect 11535 3834 11591 3836
rect 11615 3834 11671 3836
rect 11375 3782 11421 3834
rect 11421 3782 11431 3834
rect 11455 3782 11485 3834
rect 11485 3782 11497 3834
rect 11497 3782 11511 3834
rect 11535 3782 11549 3834
rect 11549 3782 11561 3834
rect 11561 3782 11591 3834
rect 11615 3782 11625 3834
rect 11625 3782 11671 3834
rect 11375 3780 11431 3782
rect 11455 3780 11511 3782
rect 11535 3780 11591 3782
rect 11615 3780 11671 3782
rect 18321 19066 18377 19068
rect 18401 19066 18457 19068
rect 18481 19066 18537 19068
rect 18561 19066 18617 19068
rect 18321 19014 18367 19066
rect 18367 19014 18377 19066
rect 18401 19014 18431 19066
rect 18431 19014 18443 19066
rect 18443 19014 18457 19066
rect 18481 19014 18495 19066
rect 18495 19014 18507 19066
rect 18507 19014 18537 19066
rect 18561 19014 18571 19066
rect 18571 19014 18617 19066
rect 18321 19012 18377 19014
rect 18401 19012 18457 19014
rect 18481 19012 18537 19014
rect 18561 19012 18617 19014
rect 21794 22874 21850 22876
rect 21874 22874 21930 22876
rect 21954 22874 22010 22876
rect 22034 22874 22090 22876
rect 21794 22822 21840 22874
rect 21840 22822 21850 22874
rect 21874 22822 21904 22874
rect 21904 22822 21916 22874
rect 21916 22822 21930 22874
rect 21954 22822 21968 22874
rect 21968 22822 21980 22874
rect 21980 22822 22010 22874
rect 22034 22822 22044 22874
rect 22044 22822 22090 22874
rect 21794 22820 21850 22822
rect 21874 22820 21930 22822
rect 21954 22820 22010 22822
rect 22034 22820 22090 22822
rect 21794 21786 21850 21788
rect 21874 21786 21930 21788
rect 21954 21786 22010 21788
rect 22034 21786 22090 21788
rect 21794 21734 21840 21786
rect 21840 21734 21850 21786
rect 21874 21734 21904 21786
rect 21904 21734 21916 21786
rect 21916 21734 21930 21786
rect 21954 21734 21968 21786
rect 21968 21734 21980 21786
rect 21980 21734 22010 21786
rect 22034 21734 22044 21786
rect 22044 21734 22090 21786
rect 21794 21732 21850 21734
rect 21874 21732 21930 21734
rect 21954 21732 22010 21734
rect 22034 21732 22090 21734
rect 18321 17978 18377 17980
rect 18401 17978 18457 17980
rect 18481 17978 18537 17980
rect 18561 17978 18617 17980
rect 18321 17926 18367 17978
rect 18367 17926 18377 17978
rect 18401 17926 18431 17978
rect 18431 17926 18443 17978
rect 18443 17926 18457 17978
rect 18481 17926 18495 17978
rect 18495 17926 18507 17978
rect 18507 17926 18537 17978
rect 18561 17926 18571 17978
rect 18571 17926 18617 17978
rect 18321 17924 18377 17926
rect 18401 17924 18457 17926
rect 18481 17924 18537 17926
rect 18561 17924 18617 17926
rect 18321 16890 18377 16892
rect 18401 16890 18457 16892
rect 18481 16890 18537 16892
rect 18561 16890 18617 16892
rect 18321 16838 18367 16890
rect 18367 16838 18377 16890
rect 18401 16838 18431 16890
rect 18431 16838 18443 16890
rect 18443 16838 18457 16890
rect 18481 16838 18495 16890
rect 18495 16838 18507 16890
rect 18507 16838 18537 16890
rect 18561 16838 18571 16890
rect 18571 16838 18617 16890
rect 18321 16836 18377 16838
rect 18401 16836 18457 16838
rect 18481 16836 18537 16838
rect 18561 16836 18617 16838
rect 18321 15802 18377 15804
rect 18401 15802 18457 15804
rect 18481 15802 18537 15804
rect 18561 15802 18617 15804
rect 18321 15750 18367 15802
rect 18367 15750 18377 15802
rect 18401 15750 18431 15802
rect 18431 15750 18443 15802
rect 18443 15750 18457 15802
rect 18481 15750 18495 15802
rect 18495 15750 18507 15802
rect 18507 15750 18537 15802
rect 18561 15750 18571 15802
rect 18571 15750 18617 15802
rect 18321 15748 18377 15750
rect 18401 15748 18457 15750
rect 18481 15748 18537 15750
rect 18561 15748 18617 15750
rect 18321 14714 18377 14716
rect 18401 14714 18457 14716
rect 18481 14714 18537 14716
rect 18561 14714 18617 14716
rect 18321 14662 18367 14714
rect 18367 14662 18377 14714
rect 18401 14662 18431 14714
rect 18431 14662 18443 14714
rect 18443 14662 18457 14714
rect 18481 14662 18495 14714
rect 18495 14662 18507 14714
rect 18507 14662 18537 14714
rect 18561 14662 18571 14714
rect 18571 14662 18617 14714
rect 18321 14660 18377 14662
rect 18401 14660 18457 14662
rect 18481 14660 18537 14662
rect 18561 14660 18617 14662
rect 14848 11994 14904 11996
rect 14928 11994 14984 11996
rect 15008 11994 15064 11996
rect 15088 11994 15144 11996
rect 14848 11942 14894 11994
rect 14894 11942 14904 11994
rect 14928 11942 14958 11994
rect 14958 11942 14970 11994
rect 14970 11942 14984 11994
rect 15008 11942 15022 11994
rect 15022 11942 15034 11994
rect 15034 11942 15064 11994
rect 15088 11942 15098 11994
rect 15098 11942 15144 11994
rect 14848 11940 14904 11942
rect 14928 11940 14984 11942
rect 15008 11940 15064 11942
rect 15088 11940 15144 11942
rect 14848 10906 14904 10908
rect 14928 10906 14984 10908
rect 15008 10906 15064 10908
rect 15088 10906 15144 10908
rect 14848 10854 14894 10906
rect 14894 10854 14904 10906
rect 14928 10854 14958 10906
rect 14958 10854 14970 10906
rect 14970 10854 14984 10906
rect 15008 10854 15022 10906
rect 15022 10854 15034 10906
rect 15034 10854 15064 10906
rect 15088 10854 15098 10906
rect 15098 10854 15144 10906
rect 14848 10852 14904 10854
rect 14928 10852 14984 10854
rect 15008 10852 15064 10854
rect 15088 10852 15144 10854
rect 14848 9818 14904 9820
rect 14928 9818 14984 9820
rect 15008 9818 15064 9820
rect 15088 9818 15144 9820
rect 14848 9766 14894 9818
rect 14894 9766 14904 9818
rect 14928 9766 14958 9818
rect 14958 9766 14970 9818
rect 14970 9766 14984 9818
rect 15008 9766 15022 9818
rect 15022 9766 15034 9818
rect 15034 9766 15064 9818
rect 15088 9766 15098 9818
rect 15098 9766 15144 9818
rect 14848 9764 14904 9766
rect 14928 9764 14984 9766
rect 15008 9764 15064 9766
rect 15088 9764 15144 9766
rect 14848 8730 14904 8732
rect 14928 8730 14984 8732
rect 15008 8730 15064 8732
rect 15088 8730 15144 8732
rect 14848 8678 14894 8730
rect 14894 8678 14904 8730
rect 14928 8678 14958 8730
rect 14958 8678 14970 8730
rect 14970 8678 14984 8730
rect 15008 8678 15022 8730
rect 15022 8678 15034 8730
rect 15034 8678 15064 8730
rect 15088 8678 15098 8730
rect 15098 8678 15144 8730
rect 14848 8676 14904 8678
rect 14928 8676 14984 8678
rect 15008 8676 15064 8678
rect 15088 8676 15144 8678
rect 14848 7642 14904 7644
rect 14928 7642 14984 7644
rect 15008 7642 15064 7644
rect 15088 7642 15144 7644
rect 14848 7590 14894 7642
rect 14894 7590 14904 7642
rect 14928 7590 14958 7642
rect 14958 7590 14970 7642
rect 14970 7590 14984 7642
rect 15008 7590 15022 7642
rect 15022 7590 15034 7642
rect 15034 7590 15064 7642
rect 15088 7590 15098 7642
rect 15098 7590 15144 7642
rect 14848 7588 14904 7590
rect 14928 7588 14984 7590
rect 15008 7588 15064 7590
rect 15088 7588 15144 7590
rect 14848 6554 14904 6556
rect 14928 6554 14984 6556
rect 15008 6554 15064 6556
rect 15088 6554 15144 6556
rect 14848 6502 14894 6554
rect 14894 6502 14904 6554
rect 14928 6502 14958 6554
rect 14958 6502 14970 6554
rect 14970 6502 14984 6554
rect 15008 6502 15022 6554
rect 15022 6502 15034 6554
rect 15034 6502 15064 6554
rect 15088 6502 15098 6554
rect 15098 6502 15144 6554
rect 14848 6500 14904 6502
rect 14928 6500 14984 6502
rect 15008 6500 15064 6502
rect 15088 6500 15144 6502
rect 14848 5466 14904 5468
rect 14928 5466 14984 5468
rect 15008 5466 15064 5468
rect 15088 5466 15144 5468
rect 14848 5414 14894 5466
rect 14894 5414 14904 5466
rect 14928 5414 14958 5466
rect 14958 5414 14970 5466
rect 14970 5414 14984 5466
rect 15008 5414 15022 5466
rect 15022 5414 15034 5466
rect 15034 5414 15064 5466
rect 15088 5414 15098 5466
rect 15098 5414 15144 5466
rect 14848 5412 14904 5414
rect 14928 5412 14984 5414
rect 15008 5412 15064 5414
rect 15088 5412 15144 5414
rect 14848 4378 14904 4380
rect 14928 4378 14984 4380
rect 15008 4378 15064 4380
rect 15088 4378 15144 4380
rect 14848 4326 14894 4378
rect 14894 4326 14904 4378
rect 14928 4326 14958 4378
rect 14958 4326 14970 4378
rect 14970 4326 14984 4378
rect 15008 4326 15022 4378
rect 15022 4326 15034 4378
rect 15034 4326 15064 4378
rect 15088 4326 15098 4378
rect 15098 4326 15144 4378
rect 14848 4324 14904 4326
rect 14928 4324 14984 4326
rect 15008 4324 15064 4326
rect 15088 4324 15144 4326
rect 11375 2746 11431 2748
rect 11455 2746 11511 2748
rect 11535 2746 11591 2748
rect 11615 2746 11671 2748
rect 11375 2694 11421 2746
rect 11421 2694 11431 2746
rect 11455 2694 11485 2746
rect 11485 2694 11497 2746
rect 11497 2694 11511 2746
rect 11535 2694 11549 2746
rect 11549 2694 11561 2746
rect 11561 2694 11591 2746
rect 11615 2694 11625 2746
rect 11625 2694 11671 2746
rect 11375 2692 11431 2694
rect 11455 2692 11511 2694
rect 11535 2692 11591 2694
rect 11615 2692 11671 2694
rect 18321 13626 18377 13628
rect 18401 13626 18457 13628
rect 18481 13626 18537 13628
rect 18561 13626 18617 13628
rect 18321 13574 18367 13626
rect 18367 13574 18377 13626
rect 18401 13574 18431 13626
rect 18431 13574 18443 13626
rect 18443 13574 18457 13626
rect 18481 13574 18495 13626
rect 18495 13574 18507 13626
rect 18507 13574 18537 13626
rect 18561 13574 18571 13626
rect 18571 13574 18617 13626
rect 18321 13572 18377 13574
rect 18401 13572 18457 13574
rect 18481 13572 18537 13574
rect 18561 13572 18617 13574
rect 18321 12538 18377 12540
rect 18401 12538 18457 12540
rect 18481 12538 18537 12540
rect 18561 12538 18617 12540
rect 18321 12486 18367 12538
rect 18367 12486 18377 12538
rect 18401 12486 18431 12538
rect 18431 12486 18443 12538
rect 18443 12486 18457 12538
rect 18481 12486 18495 12538
rect 18495 12486 18507 12538
rect 18507 12486 18537 12538
rect 18561 12486 18571 12538
rect 18571 12486 18617 12538
rect 18321 12484 18377 12486
rect 18401 12484 18457 12486
rect 18481 12484 18537 12486
rect 18561 12484 18617 12486
rect 18321 11450 18377 11452
rect 18401 11450 18457 11452
rect 18481 11450 18537 11452
rect 18561 11450 18617 11452
rect 18321 11398 18367 11450
rect 18367 11398 18377 11450
rect 18401 11398 18431 11450
rect 18431 11398 18443 11450
rect 18443 11398 18457 11450
rect 18481 11398 18495 11450
rect 18495 11398 18507 11450
rect 18507 11398 18537 11450
rect 18561 11398 18571 11450
rect 18571 11398 18617 11450
rect 18321 11396 18377 11398
rect 18401 11396 18457 11398
rect 18481 11396 18537 11398
rect 18561 11396 18617 11398
rect 18321 10362 18377 10364
rect 18401 10362 18457 10364
rect 18481 10362 18537 10364
rect 18561 10362 18617 10364
rect 18321 10310 18367 10362
rect 18367 10310 18377 10362
rect 18401 10310 18431 10362
rect 18431 10310 18443 10362
rect 18443 10310 18457 10362
rect 18481 10310 18495 10362
rect 18495 10310 18507 10362
rect 18507 10310 18537 10362
rect 18561 10310 18571 10362
rect 18571 10310 18617 10362
rect 18321 10308 18377 10310
rect 18401 10308 18457 10310
rect 18481 10308 18537 10310
rect 18561 10308 18617 10310
rect 18321 9274 18377 9276
rect 18401 9274 18457 9276
rect 18481 9274 18537 9276
rect 18561 9274 18617 9276
rect 18321 9222 18367 9274
rect 18367 9222 18377 9274
rect 18401 9222 18431 9274
rect 18431 9222 18443 9274
rect 18443 9222 18457 9274
rect 18481 9222 18495 9274
rect 18495 9222 18507 9274
rect 18507 9222 18537 9274
rect 18561 9222 18571 9274
rect 18571 9222 18617 9274
rect 18321 9220 18377 9222
rect 18401 9220 18457 9222
rect 18481 9220 18537 9222
rect 18561 9220 18617 9222
rect 18321 8186 18377 8188
rect 18401 8186 18457 8188
rect 18481 8186 18537 8188
rect 18561 8186 18617 8188
rect 18321 8134 18367 8186
rect 18367 8134 18377 8186
rect 18401 8134 18431 8186
rect 18431 8134 18443 8186
rect 18443 8134 18457 8186
rect 18481 8134 18495 8186
rect 18495 8134 18507 8186
rect 18507 8134 18537 8186
rect 18561 8134 18571 8186
rect 18571 8134 18617 8186
rect 18321 8132 18377 8134
rect 18401 8132 18457 8134
rect 18481 8132 18537 8134
rect 18561 8132 18617 8134
rect 21794 20698 21850 20700
rect 21874 20698 21930 20700
rect 21954 20698 22010 20700
rect 22034 20698 22090 20700
rect 21794 20646 21840 20698
rect 21840 20646 21850 20698
rect 21874 20646 21904 20698
rect 21904 20646 21916 20698
rect 21916 20646 21930 20698
rect 21954 20646 21968 20698
rect 21968 20646 21980 20698
rect 21980 20646 22010 20698
rect 22034 20646 22044 20698
rect 22044 20646 22090 20698
rect 21794 20644 21850 20646
rect 21874 20644 21930 20646
rect 21954 20644 22010 20646
rect 22034 20644 22090 20646
rect 21794 19610 21850 19612
rect 21874 19610 21930 19612
rect 21954 19610 22010 19612
rect 22034 19610 22090 19612
rect 21794 19558 21840 19610
rect 21840 19558 21850 19610
rect 21874 19558 21904 19610
rect 21904 19558 21916 19610
rect 21916 19558 21930 19610
rect 21954 19558 21968 19610
rect 21968 19558 21980 19610
rect 21980 19558 22010 19610
rect 22034 19558 22044 19610
rect 22044 19558 22090 19610
rect 21794 19556 21850 19558
rect 21874 19556 21930 19558
rect 21954 19556 22010 19558
rect 22034 19556 22090 19558
rect 21794 18522 21850 18524
rect 21874 18522 21930 18524
rect 21954 18522 22010 18524
rect 22034 18522 22090 18524
rect 21794 18470 21840 18522
rect 21840 18470 21850 18522
rect 21874 18470 21904 18522
rect 21904 18470 21916 18522
rect 21916 18470 21930 18522
rect 21954 18470 21968 18522
rect 21968 18470 21980 18522
rect 21980 18470 22010 18522
rect 22034 18470 22044 18522
rect 22044 18470 22090 18522
rect 21794 18468 21850 18470
rect 21874 18468 21930 18470
rect 21954 18468 22010 18470
rect 22034 18468 22090 18470
rect 21794 17434 21850 17436
rect 21874 17434 21930 17436
rect 21954 17434 22010 17436
rect 22034 17434 22090 17436
rect 21794 17382 21840 17434
rect 21840 17382 21850 17434
rect 21874 17382 21904 17434
rect 21904 17382 21916 17434
rect 21916 17382 21930 17434
rect 21954 17382 21968 17434
rect 21968 17382 21980 17434
rect 21980 17382 22010 17434
rect 22034 17382 22044 17434
rect 22044 17382 22090 17434
rect 21794 17380 21850 17382
rect 21874 17380 21930 17382
rect 21954 17380 22010 17382
rect 22034 17380 22090 17382
rect 21794 16346 21850 16348
rect 21874 16346 21930 16348
rect 21954 16346 22010 16348
rect 22034 16346 22090 16348
rect 21794 16294 21840 16346
rect 21840 16294 21850 16346
rect 21874 16294 21904 16346
rect 21904 16294 21916 16346
rect 21916 16294 21930 16346
rect 21954 16294 21968 16346
rect 21968 16294 21980 16346
rect 21980 16294 22010 16346
rect 22034 16294 22044 16346
rect 22044 16294 22090 16346
rect 21794 16292 21850 16294
rect 21874 16292 21930 16294
rect 21954 16292 22010 16294
rect 22034 16292 22090 16294
rect 21794 15258 21850 15260
rect 21874 15258 21930 15260
rect 21954 15258 22010 15260
rect 22034 15258 22090 15260
rect 21794 15206 21840 15258
rect 21840 15206 21850 15258
rect 21874 15206 21904 15258
rect 21904 15206 21916 15258
rect 21916 15206 21930 15258
rect 21954 15206 21968 15258
rect 21968 15206 21980 15258
rect 21980 15206 22010 15258
rect 22034 15206 22044 15258
rect 22044 15206 22090 15258
rect 21794 15204 21850 15206
rect 21874 15204 21930 15206
rect 21954 15204 22010 15206
rect 22034 15204 22090 15206
rect 21794 14170 21850 14172
rect 21874 14170 21930 14172
rect 21954 14170 22010 14172
rect 22034 14170 22090 14172
rect 21794 14118 21840 14170
rect 21840 14118 21850 14170
rect 21874 14118 21904 14170
rect 21904 14118 21916 14170
rect 21916 14118 21930 14170
rect 21954 14118 21968 14170
rect 21968 14118 21980 14170
rect 21980 14118 22010 14170
rect 22034 14118 22044 14170
rect 22044 14118 22090 14170
rect 21794 14116 21850 14118
rect 21874 14116 21930 14118
rect 21954 14116 22010 14118
rect 22034 14116 22090 14118
rect 21794 13082 21850 13084
rect 21874 13082 21930 13084
rect 21954 13082 22010 13084
rect 22034 13082 22090 13084
rect 21794 13030 21840 13082
rect 21840 13030 21850 13082
rect 21874 13030 21904 13082
rect 21904 13030 21916 13082
rect 21916 13030 21930 13082
rect 21954 13030 21968 13082
rect 21968 13030 21980 13082
rect 21980 13030 22010 13082
rect 22034 13030 22044 13082
rect 22044 13030 22090 13082
rect 21794 13028 21850 13030
rect 21874 13028 21930 13030
rect 21954 13028 22010 13030
rect 22034 13028 22090 13030
rect 21794 11994 21850 11996
rect 21874 11994 21930 11996
rect 21954 11994 22010 11996
rect 22034 11994 22090 11996
rect 21794 11942 21840 11994
rect 21840 11942 21850 11994
rect 21874 11942 21904 11994
rect 21904 11942 21916 11994
rect 21916 11942 21930 11994
rect 21954 11942 21968 11994
rect 21968 11942 21980 11994
rect 21980 11942 22010 11994
rect 22034 11942 22044 11994
rect 22044 11942 22090 11994
rect 21794 11940 21850 11942
rect 21874 11940 21930 11942
rect 21954 11940 22010 11942
rect 22034 11940 22090 11942
rect 21794 10906 21850 10908
rect 21874 10906 21930 10908
rect 21954 10906 22010 10908
rect 22034 10906 22090 10908
rect 21794 10854 21840 10906
rect 21840 10854 21850 10906
rect 21874 10854 21904 10906
rect 21904 10854 21916 10906
rect 21916 10854 21930 10906
rect 21954 10854 21968 10906
rect 21968 10854 21980 10906
rect 21980 10854 22010 10906
rect 22034 10854 22044 10906
rect 22044 10854 22090 10906
rect 21794 10852 21850 10854
rect 21874 10852 21930 10854
rect 21954 10852 22010 10854
rect 22034 10852 22090 10854
rect 21794 9818 21850 9820
rect 21874 9818 21930 9820
rect 21954 9818 22010 9820
rect 22034 9818 22090 9820
rect 21794 9766 21840 9818
rect 21840 9766 21850 9818
rect 21874 9766 21904 9818
rect 21904 9766 21916 9818
rect 21916 9766 21930 9818
rect 21954 9766 21968 9818
rect 21968 9766 21980 9818
rect 21980 9766 22010 9818
rect 22034 9766 22044 9818
rect 22044 9766 22090 9818
rect 21794 9764 21850 9766
rect 21874 9764 21930 9766
rect 21954 9764 22010 9766
rect 22034 9764 22090 9766
rect 25267 26682 25323 26684
rect 25347 26682 25403 26684
rect 25427 26682 25483 26684
rect 25507 26682 25563 26684
rect 25267 26630 25313 26682
rect 25313 26630 25323 26682
rect 25347 26630 25377 26682
rect 25377 26630 25389 26682
rect 25389 26630 25403 26682
rect 25427 26630 25441 26682
rect 25441 26630 25453 26682
rect 25453 26630 25483 26682
rect 25507 26630 25517 26682
rect 25517 26630 25563 26682
rect 25267 26628 25323 26630
rect 25347 26628 25403 26630
rect 25427 26628 25483 26630
rect 25507 26628 25563 26630
rect 25267 25594 25323 25596
rect 25347 25594 25403 25596
rect 25427 25594 25483 25596
rect 25507 25594 25563 25596
rect 25267 25542 25313 25594
rect 25313 25542 25323 25594
rect 25347 25542 25377 25594
rect 25377 25542 25389 25594
rect 25389 25542 25403 25594
rect 25427 25542 25441 25594
rect 25441 25542 25453 25594
rect 25453 25542 25483 25594
rect 25507 25542 25517 25594
rect 25517 25542 25563 25594
rect 25267 25540 25323 25542
rect 25347 25540 25403 25542
rect 25427 25540 25483 25542
rect 25507 25540 25563 25542
rect 25267 24506 25323 24508
rect 25347 24506 25403 24508
rect 25427 24506 25483 24508
rect 25507 24506 25563 24508
rect 25267 24454 25313 24506
rect 25313 24454 25323 24506
rect 25347 24454 25377 24506
rect 25377 24454 25389 24506
rect 25389 24454 25403 24506
rect 25427 24454 25441 24506
rect 25441 24454 25453 24506
rect 25453 24454 25483 24506
rect 25507 24454 25517 24506
rect 25517 24454 25563 24506
rect 25267 24452 25323 24454
rect 25347 24452 25403 24454
rect 25427 24452 25483 24454
rect 25507 24452 25563 24454
rect 28740 27226 28796 27228
rect 28820 27226 28876 27228
rect 28900 27226 28956 27228
rect 28980 27226 29036 27228
rect 28740 27174 28786 27226
rect 28786 27174 28796 27226
rect 28820 27174 28850 27226
rect 28850 27174 28862 27226
rect 28862 27174 28876 27226
rect 28900 27174 28914 27226
rect 28914 27174 28926 27226
rect 28926 27174 28956 27226
rect 28980 27174 28990 27226
rect 28990 27174 29036 27226
rect 28740 27172 28796 27174
rect 28820 27172 28876 27174
rect 28900 27172 28956 27174
rect 28980 27172 29036 27174
rect 28740 26138 28796 26140
rect 28820 26138 28876 26140
rect 28900 26138 28956 26140
rect 28980 26138 29036 26140
rect 28740 26086 28786 26138
rect 28786 26086 28796 26138
rect 28820 26086 28850 26138
rect 28850 26086 28862 26138
rect 28862 26086 28876 26138
rect 28900 26086 28914 26138
rect 28914 26086 28926 26138
rect 28926 26086 28956 26138
rect 28980 26086 28990 26138
rect 28990 26086 29036 26138
rect 28740 26084 28796 26086
rect 28820 26084 28876 26086
rect 28900 26084 28956 26086
rect 28980 26084 29036 26086
rect 28740 25050 28796 25052
rect 28820 25050 28876 25052
rect 28900 25050 28956 25052
rect 28980 25050 29036 25052
rect 28740 24998 28786 25050
rect 28786 24998 28796 25050
rect 28820 24998 28850 25050
rect 28850 24998 28862 25050
rect 28862 24998 28876 25050
rect 28900 24998 28914 25050
rect 28914 24998 28926 25050
rect 28926 24998 28956 25050
rect 28980 24998 28990 25050
rect 28990 24998 29036 25050
rect 28740 24996 28796 24998
rect 28820 24996 28876 24998
rect 28900 24996 28956 24998
rect 28980 24996 29036 24998
rect 25267 23418 25323 23420
rect 25347 23418 25403 23420
rect 25427 23418 25483 23420
rect 25507 23418 25563 23420
rect 25267 23366 25313 23418
rect 25313 23366 25323 23418
rect 25347 23366 25377 23418
rect 25377 23366 25389 23418
rect 25389 23366 25403 23418
rect 25427 23366 25441 23418
rect 25441 23366 25453 23418
rect 25453 23366 25483 23418
rect 25507 23366 25517 23418
rect 25517 23366 25563 23418
rect 25267 23364 25323 23366
rect 25347 23364 25403 23366
rect 25427 23364 25483 23366
rect 25507 23364 25563 23366
rect 25267 22330 25323 22332
rect 25347 22330 25403 22332
rect 25427 22330 25483 22332
rect 25507 22330 25563 22332
rect 25267 22278 25313 22330
rect 25313 22278 25323 22330
rect 25347 22278 25377 22330
rect 25377 22278 25389 22330
rect 25389 22278 25403 22330
rect 25427 22278 25441 22330
rect 25441 22278 25453 22330
rect 25453 22278 25483 22330
rect 25507 22278 25517 22330
rect 25517 22278 25563 22330
rect 25267 22276 25323 22278
rect 25347 22276 25403 22278
rect 25427 22276 25483 22278
rect 25507 22276 25563 22278
rect 25267 21242 25323 21244
rect 25347 21242 25403 21244
rect 25427 21242 25483 21244
rect 25507 21242 25563 21244
rect 25267 21190 25313 21242
rect 25313 21190 25323 21242
rect 25347 21190 25377 21242
rect 25377 21190 25389 21242
rect 25389 21190 25403 21242
rect 25427 21190 25441 21242
rect 25441 21190 25453 21242
rect 25453 21190 25483 21242
rect 25507 21190 25517 21242
rect 25517 21190 25563 21242
rect 25267 21188 25323 21190
rect 25347 21188 25403 21190
rect 25427 21188 25483 21190
rect 25507 21188 25563 21190
rect 25267 20154 25323 20156
rect 25347 20154 25403 20156
rect 25427 20154 25483 20156
rect 25507 20154 25563 20156
rect 25267 20102 25313 20154
rect 25313 20102 25323 20154
rect 25347 20102 25377 20154
rect 25377 20102 25389 20154
rect 25389 20102 25403 20154
rect 25427 20102 25441 20154
rect 25441 20102 25453 20154
rect 25453 20102 25483 20154
rect 25507 20102 25517 20154
rect 25517 20102 25563 20154
rect 25267 20100 25323 20102
rect 25347 20100 25403 20102
rect 25427 20100 25483 20102
rect 25507 20100 25563 20102
rect 28170 24132 28226 24168
rect 28170 24112 28172 24132
rect 28172 24112 28224 24132
rect 28224 24112 28226 24132
rect 28740 23962 28796 23964
rect 28820 23962 28876 23964
rect 28900 23962 28956 23964
rect 28980 23962 29036 23964
rect 28740 23910 28786 23962
rect 28786 23910 28796 23962
rect 28820 23910 28850 23962
rect 28850 23910 28862 23962
rect 28862 23910 28876 23962
rect 28900 23910 28914 23962
rect 28914 23910 28926 23962
rect 28926 23910 28956 23962
rect 28980 23910 28990 23962
rect 28990 23910 29036 23962
rect 28740 23908 28796 23910
rect 28820 23908 28876 23910
rect 28900 23908 28956 23910
rect 28980 23908 29036 23910
rect 28740 22874 28796 22876
rect 28820 22874 28876 22876
rect 28900 22874 28956 22876
rect 28980 22874 29036 22876
rect 28740 22822 28786 22874
rect 28786 22822 28796 22874
rect 28820 22822 28850 22874
rect 28850 22822 28862 22874
rect 28862 22822 28876 22874
rect 28900 22822 28914 22874
rect 28914 22822 28926 22874
rect 28926 22822 28956 22874
rect 28980 22822 28990 22874
rect 28990 22822 29036 22874
rect 28740 22820 28796 22822
rect 28820 22820 28876 22822
rect 28900 22820 28956 22822
rect 28980 22820 29036 22822
rect 28740 21786 28796 21788
rect 28820 21786 28876 21788
rect 28900 21786 28956 21788
rect 28980 21786 29036 21788
rect 28740 21734 28786 21786
rect 28786 21734 28796 21786
rect 28820 21734 28850 21786
rect 28850 21734 28862 21786
rect 28862 21734 28876 21786
rect 28900 21734 28914 21786
rect 28914 21734 28926 21786
rect 28926 21734 28956 21786
rect 28980 21734 28990 21786
rect 28990 21734 29036 21786
rect 28740 21732 28796 21734
rect 28820 21732 28876 21734
rect 28900 21732 28956 21734
rect 28980 21732 29036 21734
rect 25267 19066 25323 19068
rect 25347 19066 25403 19068
rect 25427 19066 25483 19068
rect 25507 19066 25563 19068
rect 25267 19014 25313 19066
rect 25313 19014 25323 19066
rect 25347 19014 25377 19066
rect 25377 19014 25389 19066
rect 25389 19014 25403 19066
rect 25427 19014 25441 19066
rect 25441 19014 25453 19066
rect 25453 19014 25483 19066
rect 25507 19014 25517 19066
rect 25517 19014 25563 19066
rect 25267 19012 25323 19014
rect 25347 19012 25403 19014
rect 25427 19012 25483 19014
rect 25507 19012 25563 19014
rect 25267 17978 25323 17980
rect 25347 17978 25403 17980
rect 25427 17978 25483 17980
rect 25507 17978 25563 17980
rect 25267 17926 25313 17978
rect 25313 17926 25323 17978
rect 25347 17926 25377 17978
rect 25377 17926 25389 17978
rect 25389 17926 25403 17978
rect 25427 17926 25441 17978
rect 25441 17926 25453 17978
rect 25453 17926 25483 17978
rect 25507 17926 25517 17978
rect 25517 17926 25563 17978
rect 25267 17924 25323 17926
rect 25347 17924 25403 17926
rect 25427 17924 25483 17926
rect 25507 17924 25563 17926
rect 25267 16890 25323 16892
rect 25347 16890 25403 16892
rect 25427 16890 25483 16892
rect 25507 16890 25563 16892
rect 25267 16838 25313 16890
rect 25313 16838 25323 16890
rect 25347 16838 25377 16890
rect 25377 16838 25389 16890
rect 25389 16838 25403 16890
rect 25427 16838 25441 16890
rect 25441 16838 25453 16890
rect 25453 16838 25483 16890
rect 25507 16838 25517 16890
rect 25517 16838 25563 16890
rect 25267 16836 25323 16838
rect 25347 16836 25403 16838
rect 25427 16836 25483 16838
rect 25507 16836 25563 16838
rect 21794 8730 21850 8732
rect 21874 8730 21930 8732
rect 21954 8730 22010 8732
rect 22034 8730 22090 8732
rect 21794 8678 21840 8730
rect 21840 8678 21850 8730
rect 21874 8678 21904 8730
rect 21904 8678 21916 8730
rect 21916 8678 21930 8730
rect 21954 8678 21968 8730
rect 21968 8678 21980 8730
rect 21980 8678 22010 8730
rect 22034 8678 22044 8730
rect 22044 8678 22090 8730
rect 21794 8676 21850 8678
rect 21874 8676 21930 8678
rect 21954 8676 22010 8678
rect 22034 8676 22090 8678
rect 18321 7098 18377 7100
rect 18401 7098 18457 7100
rect 18481 7098 18537 7100
rect 18561 7098 18617 7100
rect 18321 7046 18367 7098
rect 18367 7046 18377 7098
rect 18401 7046 18431 7098
rect 18431 7046 18443 7098
rect 18443 7046 18457 7098
rect 18481 7046 18495 7098
rect 18495 7046 18507 7098
rect 18507 7046 18537 7098
rect 18561 7046 18571 7098
rect 18571 7046 18617 7098
rect 18321 7044 18377 7046
rect 18401 7044 18457 7046
rect 18481 7044 18537 7046
rect 18561 7044 18617 7046
rect 21794 7642 21850 7644
rect 21874 7642 21930 7644
rect 21954 7642 22010 7644
rect 22034 7642 22090 7644
rect 21794 7590 21840 7642
rect 21840 7590 21850 7642
rect 21874 7590 21904 7642
rect 21904 7590 21916 7642
rect 21916 7590 21930 7642
rect 21954 7590 21968 7642
rect 21968 7590 21980 7642
rect 21980 7590 22010 7642
rect 22034 7590 22044 7642
rect 22044 7590 22090 7642
rect 21794 7588 21850 7590
rect 21874 7588 21930 7590
rect 21954 7588 22010 7590
rect 22034 7588 22090 7590
rect 25267 15802 25323 15804
rect 25347 15802 25403 15804
rect 25427 15802 25483 15804
rect 25507 15802 25563 15804
rect 25267 15750 25313 15802
rect 25313 15750 25323 15802
rect 25347 15750 25377 15802
rect 25377 15750 25389 15802
rect 25389 15750 25403 15802
rect 25427 15750 25441 15802
rect 25441 15750 25453 15802
rect 25453 15750 25483 15802
rect 25507 15750 25517 15802
rect 25517 15750 25563 15802
rect 25267 15748 25323 15750
rect 25347 15748 25403 15750
rect 25427 15748 25483 15750
rect 25507 15748 25563 15750
rect 25267 14714 25323 14716
rect 25347 14714 25403 14716
rect 25427 14714 25483 14716
rect 25507 14714 25563 14716
rect 25267 14662 25313 14714
rect 25313 14662 25323 14714
rect 25347 14662 25377 14714
rect 25377 14662 25389 14714
rect 25389 14662 25403 14714
rect 25427 14662 25441 14714
rect 25441 14662 25453 14714
rect 25453 14662 25483 14714
rect 25507 14662 25517 14714
rect 25517 14662 25563 14714
rect 25267 14660 25323 14662
rect 25347 14660 25403 14662
rect 25427 14660 25483 14662
rect 25507 14660 25563 14662
rect 25267 13626 25323 13628
rect 25347 13626 25403 13628
rect 25427 13626 25483 13628
rect 25507 13626 25563 13628
rect 25267 13574 25313 13626
rect 25313 13574 25323 13626
rect 25347 13574 25377 13626
rect 25377 13574 25389 13626
rect 25389 13574 25403 13626
rect 25427 13574 25441 13626
rect 25441 13574 25453 13626
rect 25453 13574 25483 13626
rect 25507 13574 25517 13626
rect 25517 13574 25563 13626
rect 25267 13572 25323 13574
rect 25347 13572 25403 13574
rect 25427 13572 25483 13574
rect 25507 13572 25563 13574
rect 25267 12538 25323 12540
rect 25347 12538 25403 12540
rect 25427 12538 25483 12540
rect 25507 12538 25563 12540
rect 25267 12486 25313 12538
rect 25313 12486 25323 12538
rect 25347 12486 25377 12538
rect 25377 12486 25389 12538
rect 25389 12486 25403 12538
rect 25427 12486 25441 12538
rect 25441 12486 25453 12538
rect 25453 12486 25483 12538
rect 25507 12486 25517 12538
rect 25517 12486 25563 12538
rect 25267 12484 25323 12486
rect 25347 12484 25403 12486
rect 25427 12484 25483 12486
rect 25507 12484 25563 12486
rect 25267 11450 25323 11452
rect 25347 11450 25403 11452
rect 25427 11450 25483 11452
rect 25507 11450 25563 11452
rect 25267 11398 25313 11450
rect 25313 11398 25323 11450
rect 25347 11398 25377 11450
rect 25377 11398 25389 11450
rect 25389 11398 25403 11450
rect 25427 11398 25441 11450
rect 25441 11398 25453 11450
rect 25453 11398 25483 11450
rect 25507 11398 25517 11450
rect 25517 11398 25563 11450
rect 25267 11396 25323 11398
rect 25347 11396 25403 11398
rect 25427 11396 25483 11398
rect 25507 11396 25563 11398
rect 25267 10362 25323 10364
rect 25347 10362 25403 10364
rect 25427 10362 25483 10364
rect 25507 10362 25563 10364
rect 25267 10310 25313 10362
rect 25313 10310 25323 10362
rect 25347 10310 25377 10362
rect 25377 10310 25389 10362
rect 25389 10310 25403 10362
rect 25427 10310 25441 10362
rect 25441 10310 25453 10362
rect 25453 10310 25483 10362
rect 25507 10310 25517 10362
rect 25517 10310 25563 10362
rect 25267 10308 25323 10310
rect 25347 10308 25403 10310
rect 25427 10308 25483 10310
rect 25507 10308 25563 10310
rect 25267 9274 25323 9276
rect 25347 9274 25403 9276
rect 25427 9274 25483 9276
rect 25507 9274 25563 9276
rect 25267 9222 25313 9274
rect 25313 9222 25323 9274
rect 25347 9222 25377 9274
rect 25377 9222 25389 9274
rect 25389 9222 25403 9274
rect 25427 9222 25441 9274
rect 25441 9222 25453 9274
rect 25453 9222 25483 9274
rect 25507 9222 25517 9274
rect 25517 9222 25563 9274
rect 25267 9220 25323 9222
rect 25347 9220 25403 9222
rect 25427 9220 25483 9222
rect 25507 9220 25563 9222
rect 28740 20698 28796 20700
rect 28820 20698 28876 20700
rect 28900 20698 28956 20700
rect 28980 20698 29036 20700
rect 28740 20646 28786 20698
rect 28786 20646 28796 20698
rect 28820 20646 28850 20698
rect 28850 20646 28862 20698
rect 28862 20646 28876 20698
rect 28900 20646 28914 20698
rect 28914 20646 28926 20698
rect 28926 20646 28956 20698
rect 28980 20646 28990 20698
rect 28990 20646 29036 20698
rect 28740 20644 28796 20646
rect 28820 20644 28876 20646
rect 28900 20644 28956 20646
rect 28980 20644 29036 20646
rect 28170 20440 28226 20496
rect 28740 19610 28796 19612
rect 28820 19610 28876 19612
rect 28900 19610 28956 19612
rect 28980 19610 29036 19612
rect 28740 19558 28786 19610
rect 28786 19558 28796 19610
rect 28820 19558 28850 19610
rect 28850 19558 28862 19610
rect 28862 19558 28876 19610
rect 28900 19558 28914 19610
rect 28914 19558 28926 19610
rect 28926 19558 28956 19610
rect 28980 19558 28990 19610
rect 28990 19558 29036 19610
rect 28740 19556 28796 19558
rect 28820 19556 28876 19558
rect 28900 19556 28956 19558
rect 28980 19556 29036 19558
rect 28740 18522 28796 18524
rect 28820 18522 28876 18524
rect 28900 18522 28956 18524
rect 28980 18522 29036 18524
rect 28740 18470 28786 18522
rect 28786 18470 28796 18522
rect 28820 18470 28850 18522
rect 28850 18470 28862 18522
rect 28862 18470 28876 18522
rect 28900 18470 28914 18522
rect 28914 18470 28926 18522
rect 28926 18470 28956 18522
rect 28980 18470 28990 18522
rect 28990 18470 29036 18522
rect 28740 18468 28796 18470
rect 28820 18468 28876 18470
rect 28900 18468 28956 18470
rect 28980 18468 29036 18470
rect 28740 17434 28796 17436
rect 28820 17434 28876 17436
rect 28900 17434 28956 17436
rect 28980 17434 29036 17436
rect 28740 17382 28786 17434
rect 28786 17382 28796 17434
rect 28820 17382 28850 17434
rect 28850 17382 28862 17434
rect 28862 17382 28876 17434
rect 28900 17382 28914 17434
rect 28914 17382 28926 17434
rect 28926 17382 28956 17434
rect 28980 17382 28990 17434
rect 28990 17382 29036 17434
rect 28740 17380 28796 17382
rect 28820 17380 28876 17382
rect 28900 17380 28956 17382
rect 28980 17380 29036 17382
rect 28170 16768 28226 16824
rect 28740 16346 28796 16348
rect 28820 16346 28876 16348
rect 28900 16346 28956 16348
rect 28980 16346 29036 16348
rect 28740 16294 28786 16346
rect 28786 16294 28796 16346
rect 28820 16294 28850 16346
rect 28850 16294 28862 16346
rect 28862 16294 28876 16346
rect 28900 16294 28914 16346
rect 28914 16294 28926 16346
rect 28926 16294 28956 16346
rect 28980 16294 28990 16346
rect 28990 16294 29036 16346
rect 28740 16292 28796 16294
rect 28820 16292 28876 16294
rect 28900 16292 28956 16294
rect 28980 16292 29036 16294
rect 28740 15258 28796 15260
rect 28820 15258 28876 15260
rect 28900 15258 28956 15260
rect 28980 15258 29036 15260
rect 28740 15206 28786 15258
rect 28786 15206 28796 15258
rect 28820 15206 28850 15258
rect 28850 15206 28862 15258
rect 28862 15206 28876 15258
rect 28900 15206 28914 15258
rect 28914 15206 28926 15258
rect 28926 15206 28956 15258
rect 28980 15206 28990 15258
rect 28990 15206 29036 15258
rect 28740 15204 28796 15206
rect 28820 15204 28876 15206
rect 28900 15204 28956 15206
rect 28980 15204 29036 15206
rect 28740 14170 28796 14172
rect 28820 14170 28876 14172
rect 28900 14170 28956 14172
rect 28980 14170 29036 14172
rect 28740 14118 28786 14170
rect 28786 14118 28796 14170
rect 28820 14118 28850 14170
rect 28850 14118 28862 14170
rect 28862 14118 28876 14170
rect 28900 14118 28914 14170
rect 28914 14118 28926 14170
rect 28926 14118 28956 14170
rect 28980 14118 28990 14170
rect 28990 14118 29036 14170
rect 28740 14116 28796 14118
rect 28820 14116 28876 14118
rect 28900 14116 28956 14118
rect 28980 14116 29036 14118
rect 28170 13232 28226 13288
rect 28740 13082 28796 13084
rect 28820 13082 28876 13084
rect 28900 13082 28956 13084
rect 28980 13082 29036 13084
rect 28740 13030 28786 13082
rect 28786 13030 28796 13082
rect 28820 13030 28850 13082
rect 28850 13030 28862 13082
rect 28862 13030 28876 13082
rect 28900 13030 28914 13082
rect 28914 13030 28926 13082
rect 28926 13030 28956 13082
rect 28980 13030 28990 13082
rect 28990 13030 29036 13082
rect 28740 13028 28796 13030
rect 28820 13028 28876 13030
rect 28900 13028 28956 13030
rect 28980 13028 29036 13030
rect 28740 11994 28796 11996
rect 28820 11994 28876 11996
rect 28900 11994 28956 11996
rect 28980 11994 29036 11996
rect 28740 11942 28786 11994
rect 28786 11942 28796 11994
rect 28820 11942 28850 11994
rect 28850 11942 28862 11994
rect 28862 11942 28876 11994
rect 28900 11942 28914 11994
rect 28914 11942 28926 11994
rect 28926 11942 28956 11994
rect 28980 11942 28990 11994
rect 28990 11942 29036 11994
rect 28740 11940 28796 11942
rect 28820 11940 28876 11942
rect 28900 11940 28956 11942
rect 28980 11940 29036 11942
rect 28740 10906 28796 10908
rect 28820 10906 28876 10908
rect 28900 10906 28956 10908
rect 28980 10906 29036 10908
rect 28740 10854 28786 10906
rect 28786 10854 28796 10906
rect 28820 10854 28850 10906
rect 28850 10854 28862 10906
rect 28862 10854 28876 10906
rect 28900 10854 28914 10906
rect 28914 10854 28926 10906
rect 28926 10854 28956 10906
rect 28980 10854 28990 10906
rect 28990 10854 29036 10906
rect 28740 10852 28796 10854
rect 28820 10852 28876 10854
rect 28900 10852 28956 10854
rect 28980 10852 29036 10854
rect 18321 6010 18377 6012
rect 18401 6010 18457 6012
rect 18481 6010 18537 6012
rect 18561 6010 18617 6012
rect 18321 5958 18367 6010
rect 18367 5958 18377 6010
rect 18401 5958 18431 6010
rect 18431 5958 18443 6010
rect 18443 5958 18457 6010
rect 18481 5958 18495 6010
rect 18495 5958 18507 6010
rect 18507 5958 18537 6010
rect 18561 5958 18571 6010
rect 18571 5958 18617 6010
rect 18321 5956 18377 5958
rect 18401 5956 18457 5958
rect 18481 5956 18537 5958
rect 18561 5956 18617 5958
rect 18321 4922 18377 4924
rect 18401 4922 18457 4924
rect 18481 4922 18537 4924
rect 18561 4922 18617 4924
rect 18321 4870 18367 4922
rect 18367 4870 18377 4922
rect 18401 4870 18431 4922
rect 18431 4870 18443 4922
rect 18443 4870 18457 4922
rect 18481 4870 18495 4922
rect 18495 4870 18507 4922
rect 18507 4870 18537 4922
rect 18561 4870 18571 4922
rect 18571 4870 18617 4922
rect 18321 4868 18377 4870
rect 18401 4868 18457 4870
rect 18481 4868 18537 4870
rect 18561 4868 18617 4870
rect 21794 6554 21850 6556
rect 21874 6554 21930 6556
rect 21954 6554 22010 6556
rect 22034 6554 22090 6556
rect 21794 6502 21840 6554
rect 21840 6502 21850 6554
rect 21874 6502 21904 6554
rect 21904 6502 21916 6554
rect 21916 6502 21930 6554
rect 21954 6502 21968 6554
rect 21968 6502 21980 6554
rect 21980 6502 22010 6554
rect 22034 6502 22044 6554
rect 22044 6502 22090 6554
rect 21794 6500 21850 6502
rect 21874 6500 21930 6502
rect 21954 6500 22010 6502
rect 22034 6500 22090 6502
rect 18321 3834 18377 3836
rect 18401 3834 18457 3836
rect 18481 3834 18537 3836
rect 18561 3834 18617 3836
rect 18321 3782 18367 3834
rect 18367 3782 18377 3834
rect 18401 3782 18431 3834
rect 18431 3782 18443 3834
rect 18443 3782 18457 3834
rect 18481 3782 18495 3834
rect 18495 3782 18507 3834
rect 18507 3782 18537 3834
rect 18561 3782 18571 3834
rect 18571 3782 18617 3834
rect 18321 3780 18377 3782
rect 18401 3780 18457 3782
rect 18481 3780 18537 3782
rect 18561 3780 18617 3782
rect 14848 3290 14904 3292
rect 14928 3290 14984 3292
rect 15008 3290 15064 3292
rect 15088 3290 15144 3292
rect 14848 3238 14894 3290
rect 14894 3238 14904 3290
rect 14928 3238 14958 3290
rect 14958 3238 14970 3290
rect 14970 3238 14984 3290
rect 15008 3238 15022 3290
rect 15022 3238 15034 3290
rect 15034 3238 15064 3290
rect 15088 3238 15098 3290
rect 15098 3238 15144 3290
rect 14848 3236 14904 3238
rect 14928 3236 14984 3238
rect 15008 3236 15064 3238
rect 15088 3236 15144 3238
rect 21794 5466 21850 5468
rect 21874 5466 21930 5468
rect 21954 5466 22010 5468
rect 22034 5466 22090 5468
rect 21794 5414 21840 5466
rect 21840 5414 21850 5466
rect 21874 5414 21904 5466
rect 21904 5414 21916 5466
rect 21916 5414 21930 5466
rect 21954 5414 21968 5466
rect 21968 5414 21980 5466
rect 21980 5414 22010 5466
rect 22034 5414 22044 5466
rect 22044 5414 22090 5466
rect 21794 5412 21850 5414
rect 21874 5412 21930 5414
rect 21954 5412 22010 5414
rect 22034 5412 22090 5414
rect 21794 4378 21850 4380
rect 21874 4378 21930 4380
rect 21954 4378 22010 4380
rect 22034 4378 22090 4380
rect 21794 4326 21840 4378
rect 21840 4326 21850 4378
rect 21874 4326 21904 4378
rect 21904 4326 21916 4378
rect 21916 4326 21930 4378
rect 21954 4326 21968 4378
rect 21968 4326 21980 4378
rect 21980 4326 22010 4378
rect 22034 4326 22044 4378
rect 22044 4326 22090 4378
rect 21794 4324 21850 4326
rect 21874 4324 21930 4326
rect 21954 4324 22010 4326
rect 22034 4324 22090 4326
rect 25267 8186 25323 8188
rect 25347 8186 25403 8188
rect 25427 8186 25483 8188
rect 25507 8186 25563 8188
rect 25267 8134 25313 8186
rect 25313 8134 25323 8186
rect 25347 8134 25377 8186
rect 25377 8134 25389 8186
rect 25389 8134 25403 8186
rect 25427 8134 25441 8186
rect 25441 8134 25453 8186
rect 25453 8134 25483 8186
rect 25507 8134 25517 8186
rect 25517 8134 25563 8186
rect 25267 8132 25323 8134
rect 25347 8132 25403 8134
rect 25427 8132 25483 8134
rect 25507 8132 25563 8134
rect 25267 7098 25323 7100
rect 25347 7098 25403 7100
rect 25427 7098 25483 7100
rect 25507 7098 25563 7100
rect 25267 7046 25313 7098
rect 25313 7046 25323 7098
rect 25347 7046 25377 7098
rect 25377 7046 25389 7098
rect 25389 7046 25403 7098
rect 25427 7046 25441 7098
rect 25441 7046 25453 7098
rect 25453 7046 25483 7098
rect 25507 7046 25517 7098
rect 25517 7046 25563 7098
rect 25267 7044 25323 7046
rect 25347 7044 25403 7046
rect 25427 7044 25483 7046
rect 25507 7044 25563 7046
rect 25267 6010 25323 6012
rect 25347 6010 25403 6012
rect 25427 6010 25483 6012
rect 25507 6010 25563 6012
rect 25267 5958 25313 6010
rect 25313 5958 25323 6010
rect 25347 5958 25377 6010
rect 25377 5958 25389 6010
rect 25389 5958 25403 6010
rect 25427 5958 25441 6010
rect 25441 5958 25453 6010
rect 25453 5958 25483 6010
rect 25507 5958 25517 6010
rect 25517 5958 25563 6010
rect 25267 5956 25323 5958
rect 25347 5956 25403 5958
rect 25427 5956 25483 5958
rect 25507 5956 25563 5958
rect 26422 7692 26424 7712
rect 26424 7692 26476 7712
rect 26476 7692 26478 7712
rect 26422 7656 26478 7692
rect 21794 3290 21850 3292
rect 21874 3290 21930 3292
rect 21954 3290 22010 3292
rect 22034 3290 22090 3292
rect 21794 3238 21840 3290
rect 21840 3238 21850 3290
rect 21874 3238 21904 3290
rect 21904 3238 21916 3290
rect 21916 3238 21930 3290
rect 21954 3238 21968 3290
rect 21968 3238 21980 3290
rect 21980 3238 22010 3290
rect 22034 3238 22044 3290
rect 22044 3238 22090 3290
rect 21794 3236 21850 3238
rect 21874 3236 21930 3238
rect 21954 3236 22010 3238
rect 22034 3236 22090 3238
rect 25267 4922 25323 4924
rect 25347 4922 25403 4924
rect 25427 4922 25483 4924
rect 25507 4922 25563 4924
rect 25267 4870 25313 4922
rect 25313 4870 25323 4922
rect 25347 4870 25377 4922
rect 25377 4870 25389 4922
rect 25389 4870 25403 4922
rect 25427 4870 25441 4922
rect 25441 4870 25453 4922
rect 25453 4870 25483 4922
rect 25507 4870 25517 4922
rect 25517 4870 25563 4922
rect 25267 4868 25323 4870
rect 25347 4868 25403 4870
rect 25427 4868 25483 4870
rect 25507 4868 25563 4870
rect 25267 3834 25323 3836
rect 25347 3834 25403 3836
rect 25427 3834 25483 3836
rect 25507 3834 25563 3836
rect 25267 3782 25313 3834
rect 25313 3782 25323 3834
rect 25347 3782 25377 3834
rect 25377 3782 25389 3834
rect 25389 3782 25403 3834
rect 25427 3782 25441 3834
rect 25441 3782 25453 3834
rect 25453 3782 25483 3834
rect 25507 3782 25517 3834
rect 25517 3782 25563 3834
rect 25267 3780 25323 3782
rect 25347 3780 25403 3782
rect 25427 3780 25483 3782
rect 25507 3780 25563 3782
rect 28740 9818 28796 9820
rect 28820 9818 28876 9820
rect 28900 9818 28956 9820
rect 28980 9818 29036 9820
rect 28740 9766 28786 9818
rect 28786 9766 28796 9818
rect 28820 9766 28850 9818
rect 28850 9766 28862 9818
rect 28862 9766 28876 9818
rect 28900 9766 28914 9818
rect 28914 9766 28926 9818
rect 28926 9766 28956 9818
rect 28980 9766 28990 9818
rect 28990 9766 29036 9818
rect 28740 9764 28796 9766
rect 28820 9764 28876 9766
rect 28900 9764 28956 9766
rect 28980 9764 29036 9766
rect 28170 9424 28226 9480
rect 28740 8730 28796 8732
rect 28820 8730 28876 8732
rect 28900 8730 28956 8732
rect 28980 8730 29036 8732
rect 28740 8678 28786 8730
rect 28786 8678 28796 8730
rect 28820 8678 28850 8730
rect 28850 8678 28862 8730
rect 28862 8678 28876 8730
rect 28900 8678 28914 8730
rect 28914 8678 28926 8730
rect 28926 8678 28956 8730
rect 28980 8678 28990 8730
rect 28990 8678 29036 8730
rect 28740 8676 28796 8678
rect 28820 8676 28876 8678
rect 28900 8676 28956 8678
rect 28980 8676 29036 8678
rect 27618 7692 27620 7712
rect 27620 7692 27672 7712
rect 27672 7692 27674 7712
rect 27618 7656 27674 7692
rect 28740 7642 28796 7644
rect 28820 7642 28876 7644
rect 28900 7642 28956 7644
rect 28980 7642 29036 7644
rect 28740 7590 28786 7642
rect 28786 7590 28796 7642
rect 28820 7590 28850 7642
rect 28850 7590 28862 7642
rect 28862 7590 28876 7642
rect 28900 7590 28914 7642
rect 28914 7590 28926 7642
rect 28926 7590 28956 7642
rect 28980 7590 28990 7642
rect 28990 7590 29036 7642
rect 28740 7588 28796 7590
rect 28820 7588 28876 7590
rect 28900 7588 28956 7590
rect 28980 7588 29036 7590
rect 28740 6554 28796 6556
rect 28820 6554 28876 6556
rect 28900 6554 28956 6556
rect 28980 6554 29036 6556
rect 28740 6502 28786 6554
rect 28786 6502 28796 6554
rect 28820 6502 28850 6554
rect 28850 6502 28862 6554
rect 28862 6502 28876 6554
rect 28900 6502 28914 6554
rect 28914 6502 28926 6554
rect 28926 6502 28956 6554
rect 28980 6502 28990 6554
rect 28990 6502 29036 6554
rect 28740 6500 28796 6502
rect 28820 6500 28876 6502
rect 28900 6500 28956 6502
rect 28980 6500 29036 6502
rect 28170 5752 28226 5808
rect 28740 5466 28796 5468
rect 28820 5466 28876 5468
rect 28900 5466 28956 5468
rect 28980 5466 29036 5468
rect 28740 5414 28786 5466
rect 28786 5414 28796 5466
rect 28820 5414 28850 5466
rect 28850 5414 28862 5466
rect 28862 5414 28876 5466
rect 28900 5414 28914 5466
rect 28914 5414 28926 5466
rect 28926 5414 28956 5466
rect 28980 5414 28990 5466
rect 28990 5414 29036 5466
rect 28740 5412 28796 5414
rect 28820 5412 28876 5414
rect 28900 5412 28956 5414
rect 28980 5412 29036 5414
rect 28740 4378 28796 4380
rect 28820 4378 28876 4380
rect 28900 4378 28956 4380
rect 28980 4378 29036 4380
rect 28740 4326 28786 4378
rect 28786 4326 28796 4378
rect 28820 4326 28850 4378
rect 28850 4326 28862 4378
rect 28862 4326 28876 4378
rect 28900 4326 28914 4378
rect 28914 4326 28926 4378
rect 28926 4326 28956 4378
rect 28980 4326 28990 4378
rect 28990 4326 29036 4378
rect 28740 4324 28796 4326
rect 28820 4324 28876 4326
rect 28900 4324 28956 4326
rect 28980 4324 29036 4326
rect 28740 3290 28796 3292
rect 28820 3290 28876 3292
rect 28900 3290 28956 3292
rect 28980 3290 29036 3292
rect 28740 3238 28786 3290
rect 28786 3238 28796 3290
rect 28820 3238 28850 3290
rect 28850 3238 28862 3290
rect 28862 3238 28876 3290
rect 28900 3238 28914 3290
rect 28914 3238 28926 3290
rect 28926 3238 28956 3290
rect 28980 3238 28990 3290
rect 28990 3238 29036 3290
rect 28740 3236 28796 3238
rect 28820 3236 28876 3238
rect 28900 3236 28956 3238
rect 28980 3236 29036 3238
rect 18321 2746 18377 2748
rect 18401 2746 18457 2748
rect 18481 2746 18537 2748
rect 18561 2746 18617 2748
rect 18321 2694 18367 2746
rect 18367 2694 18377 2746
rect 18401 2694 18431 2746
rect 18431 2694 18443 2746
rect 18443 2694 18457 2746
rect 18481 2694 18495 2746
rect 18495 2694 18507 2746
rect 18507 2694 18537 2746
rect 18561 2694 18571 2746
rect 18571 2694 18617 2746
rect 18321 2692 18377 2694
rect 18401 2692 18457 2694
rect 18481 2692 18537 2694
rect 18561 2692 18617 2694
rect 25267 2746 25323 2748
rect 25347 2746 25403 2748
rect 25427 2746 25483 2748
rect 25507 2746 25563 2748
rect 25267 2694 25313 2746
rect 25313 2694 25323 2746
rect 25347 2694 25377 2746
rect 25377 2694 25389 2746
rect 25389 2694 25403 2746
rect 25427 2694 25441 2746
rect 25441 2694 25453 2746
rect 25453 2694 25483 2746
rect 25507 2694 25517 2746
rect 25517 2694 25563 2746
rect 25267 2692 25323 2694
rect 25347 2692 25403 2694
rect 25427 2692 25483 2694
rect 25507 2692 25563 2694
rect 28170 2372 28226 2408
rect 28170 2352 28172 2372
rect 28172 2352 28224 2372
rect 28224 2352 28226 2372
rect 7902 2202 7958 2204
rect 7982 2202 8038 2204
rect 8062 2202 8118 2204
rect 8142 2202 8198 2204
rect 7902 2150 7948 2202
rect 7948 2150 7958 2202
rect 7982 2150 8012 2202
rect 8012 2150 8024 2202
rect 8024 2150 8038 2202
rect 8062 2150 8076 2202
rect 8076 2150 8088 2202
rect 8088 2150 8118 2202
rect 8142 2150 8152 2202
rect 8152 2150 8198 2202
rect 7902 2148 7958 2150
rect 7982 2148 8038 2150
rect 8062 2148 8118 2150
rect 8142 2148 8198 2150
rect 14848 2202 14904 2204
rect 14928 2202 14984 2204
rect 15008 2202 15064 2204
rect 15088 2202 15144 2204
rect 14848 2150 14894 2202
rect 14894 2150 14904 2202
rect 14928 2150 14958 2202
rect 14958 2150 14970 2202
rect 14970 2150 14984 2202
rect 15008 2150 15022 2202
rect 15022 2150 15034 2202
rect 15034 2150 15064 2202
rect 15088 2150 15098 2202
rect 15098 2150 15144 2202
rect 14848 2148 14904 2150
rect 14928 2148 14984 2150
rect 15008 2148 15064 2150
rect 15088 2148 15144 2150
rect 21794 2202 21850 2204
rect 21874 2202 21930 2204
rect 21954 2202 22010 2204
rect 22034 2202 22090 2204
rect 21794 2150 21840 2202
rect 21840 2150 21850 2202
rect 21874 2150 21904 2202
rect 21904 2150 21916 2202
rect 21916 2150 21930 2202
rect 21954 2150 21968 2202
rect 21968 2150 21980 2202
rect 21980 2150 22010 2202
rect 22034 2150 22044 2202
rect 22044 2150 22090 2202
rect 21794 2148 21850 2150
rect 21874 2148 21930 2150
rect 21954 2148 22010 2150
rect 22034 2148 22090 2150
rect 28740 2202 28796 2204
rect 28820 2202 28876 2204
rect 28900 2202 28956 2204
rect 28980 2202 29036 2204
rect 28740 2150 28786 2202
rect 28786 2150 28796 2202
rect 28820 2150 28850 2202
rect 28850 2150 28862 2202
rect 28862 2150 28876 2202
rect 28900 2150 28914 2202
rect 28914 2150 28926 2202
rect 28926 2150 28956 2202
rect 28980 2150 28990 2202
rect 28990 2150 29036 2202
rect 28740 2148 28796 2150
rect 28820 2148 28876 2150
rect 28900 2148 28956 2150
rect 28980 2148 29036 2150
<< metal3 >>
rect 27521 27842 27587 27845
rect 29200 27842 30000 27872
rect 27521 27840 30000 27842
rect 27521 27784 27526 27840
rect 27582 27784 30000 27840
rect 27521 27782 30000 27784
rect 27521 27779 27587 27782
rect 4419 27776 4735 27777
rect 4419 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4735 27776
rect 4419 27711 4735 27712
rect 11365 27776 11681 27777
rect 11365 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11681 27776
rect 11365 27711 11681 27712
rect 18311 27776 18627 27777
rect 18311 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18627 27776
rect 18311 27711 18627 27712
rect 25257 27776 25573 27777
rect 25257 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25573 27776
rect 29200 27752 30000 27782
rect 25257 27711 25573 27712
rect 7892 27232 8208 27233
rect 7892 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8208 27232
rect 7892 27167 8208 27168
rect 14838 27232 15154 27233
rect 14838 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15154 27232
rect 14838 27167 15154 27168
rect 21784 27232 22100 27233
rect 21784 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22100 27232
rect 21784 27167 22100 27168
rect 28730 27232 29046 27233
rect 28730 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29046 27232
rect 28730 27167 29046 27168
rect 4419 26688 4735 26689
rect 4419 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4735 26688
rect 4419 26623 4735 26624
rect 11365 26688 11681 26689
rect 11365 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11681 26688
rect 11365 26623 11681 26624
rect 18311 26688 18627 26689
rect 18311 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18627 26688
rect 18311 26623 18627 26624
rect 25257 26688 25573 26689
rect 25257 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25573 26688
rect 25257 26623 25573 26624
rect 7892 26144 8208 26145
rect 7892 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8208 26144
rect 7892 26079 8208 26080
rect 14838 26144 15154 26145
rect 14838 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15154 26144
rect 14838 26079 15154 26080
rect 21784 26144 22100 26145
rect 21784 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22100 26144
rect 21784 26079 22100 26080
rect 28730 26144 29046 26145
rect 28730 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29046 26144
rect 28730 26079 29046 26080
rect 4419 25600 4735 25601
rect 4419 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4735 25600
rect 4419 25535 4735 25536
rect 11365 25600 11681 25601
rect 11365 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11681 25600
rect 11365 25535 11681 25536
rect 18311 25600 18627 25601
rect 18311 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18627 25600
rect 18311 25535 18627 25536
rect 25257 25600 25573 25601
rect 25257 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25573 25600
rect 25257 25535 25573 25536
rect 7892 25056 8208 25057
rect 7892 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8208 25056
rect 7892 24991 8208 24992
rect 14838 25056 15154 25057
rect 14838 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15154 25056
rect 14838 24991 15154 24992
rect 21784 25056 22100 25057
rect 21784 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22100 25056
rect 21784 24991 22100 24992
rect 28730 25056 29046 25057
rect 28730 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29046 25056
rect 28730 24991 29046 24992
rect 4419 24512 4735 24513
rect 4419 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4735 24512
rect 4419 24447 4735 24448
rect 11365 24512 11681 24513
rect 11365 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11681 24512
rect 11365 24447 11681 24448
rect 18311 24512 18627 24513
rect 18311 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18627 24512
rect 18311 24447 18627 24448
rect 25257 24512 25573 24513
rect 25257 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25573 24512
rect 25257 24447 25573 24448
rect 28165 24170 28231 24173
rect 29200 24170 30000 24200
rect 28165 24168 30000 24170
rect 28165 24112 28170 24168
rect 28226 24112 30000 24168
rect 28165 24110 30000 24112
rect 28165 24107 28231 24110
rect 29200 24080 30000 24110
rect 7892 23968 8208 23969
rect 7892 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8208 23968
rect 7892 23903 8208 23904
rect 14838 23968 15154 23969
rect 14838 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15154 23968
rect 14838 23903 15154 23904
rect 21784 23968 22100 23969
rect 21784 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22100 23968
rect 21784 23903 22100 23904
rect 28730 23968 29046 23969
rect 28730 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29046 23968
rect 28730 23903 29046 23904
rect 4419 23424 4735 23425
rect 4419 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4735 23424
rect 4419 23359 4735 23360
rect 11365 23424 11681 23425
rect 11365 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11681 23424
rect 11365 23359 11681 23360
rect 18311 23424 18627 23425
rect 18311 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18627 23424
rect 18311 23359 18627 23360
rect 25257 23424 25573 23425
rect 25257 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25573 23424
rect 25257 23359 25573 23360
rect 7892 22880 8208 22881
rect 7892 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8208 22880
rect 7892 22815 8208 22816
rect 14838 22880 15154 22881
rect 14838 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15154 22880
rect 14838 22815 15154 22816
rect 21784 22880 22100 22881
rect 21784 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22100 22880
rect 21784 22815 22100 22816
rect 28730 22880 29046 22881
rect 28730 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29046 22880
rect 28730 22815 29046 22816
rect 4419 22336 4735 22337
rect 4419 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4735 22336
rect 4419 22271 4735 22272
rect 11365 22336 11681 22337
rect 11365 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11681 22336
rect 11365 22271 11681 22272
rect 18311 22336 18627 22337
rect 18311 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18627 22336
rect 18311 22271 18627 22272
rect 25257 22336 25573 22337
rect 25257 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25573 22336
rect 25257 22271 25573 22272
rect 7892 21792 8208 21793
rect 7892 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8208 21792
rect 7892 21727 8208 21728
rect 14838 21792 15154 21793
rect 14838 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15154 21792
rect 14838 21727 15154 21728
rect 21784 21792 22100 21793
rect 21784 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22100 21792
rect 21784 21727 22100 21728
rect 28730 21792 29046 21793
rect 28730 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29046 21792
rect 28730 21727 29046 21728
rect 4419 21248 4735 21249
rect 4419 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4735 21248
rect 4419 21183 4735 21184
rect 11365 21248 11681 21249
rect 11365 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11681 21248
rect 11365 21183 11681 21184
rect 18311 21248 18627 21249
rect 18311 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18627 21248
rect 18311 21183 18627 21184
rect 25257 21248 25573 21249
rect 25257 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25573 21248
rect 25257 21183 25573 21184
rect 7892 20704 8208 20705
rect 7892 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8208 20704
rect 7892 20639 8208 20640
rect 14838 20704 15154 20705
rect 14838 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15154 20704
rect 14838 20639 15154 20640
rect 21784 20704 22100 20705
rect 21784 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22100 20704
rect 21784 20639 22100 20640
rect 28730 20704 29046 20705
rect 28730 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29046 20704
rect 28730 20639 29046 20640
rect 28165 20498 28231 20501
rect 29200 20498 30000 20528
rect 28165 20496 30000 20498
rect 28165 20440 28170 20496
rect 28226 20440 30000 20496
rect 28165 20438 30000 20440
rect 28165 20435 28231 20438
rect 29200 20408 30000 20438
rect 4419 20160 4735 20161
rect 4419 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4735 20160
rect 4419 20095 4735 20096
rect 11365 20160 11681 20161
rect 11365 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11681 20160
rect 11365 20095 11681 20096
rect 18311 20160 18627 20161
rect 18311 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18627 20160
rect 18311 20095 18627 20096
rect 25257 20160 25573 20161
rect 25257 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25573 20160
rect 25257 20095 25573 20096
rect 7892 19616 8208 19617
rect 7892 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8208 19616
rect 7892 19551 8208 19552
rect 14838 19616 15154 19617
rect 14838 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15154 19616
rect 14838 19551 15154 19552
rect 21784 19616 22100 19617
rect 21784 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22100 19616
rect 21784 19551 22100 19552
rect 28730 19616 29046 19617
rect 28730 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29046 19616
rect 28730 19551 29046 19552
rect 4419 19072 4735 19073
rect 4419 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4735 19072
rect 4419 19007 4735 19008
rect 11365 19072 11681 19073
rect 11365 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11681 19072
rect 11365 19007 11681 19008
rect 18311 19072 18627 19073
rect 18311 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18627 19072
rect 18311 19007 18627 19008
rect 25257 19072 25573 19073
rect 25257 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25573 19072
rect 25257 19007 25573 19008
rect 7892 18528 8208 18529
rect 7892 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8208 18528
rect 7892 18463 8208 18464
rect 14838 18528 15154 18529
rect 14838 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15154 18528
rect 14838 18463 15154 18464
rect 21784 18528 22100 18529
rect 21784 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22100 18528
rect 21784 18463 22100 18464
rect 28730 18528 29046 18529
rect 28730 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29046 18528
rect 28730 18463 29046 18464
rect 4419 17984 4735 17985
rect 4419 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4735 17984
rect 4419 17919 4735 17920
rect 11365 17984 11681 17985
rect 11365 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11681 17984
rect 11365 17919 11681 17920
rect 18311 17984 18627 17985
rect 18311 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18627 17984
rect 18311 17919 18627 17920
rect 25257 17984 25573 17985
rect 25257 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25573 17984
rect 25257 17919 25573 17920
rect 7892 17440 8208 17441
rect 7892 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8208 17440
rect 7892 17375 8208 17376
rect 14838 17440 15154 17441
rect 14838 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15154 17440
rect 14838 17375 15154 17376
rect 21784 17440 22100 17441
rect 21784 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22100 17440
rect 21784 17375 22100 17376
rect 28730 17440 29046 17441
rect 28730 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29046 17440
rect 28730 17375 29046 17376
rect 4419 16896 4735 16897
rect 4419 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4735 16896
rect 4419 16831 4735 16832
rect 11365 16896 11681 16897
rect 11365 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11681 16896
rect 11365 16831 11681 16832
rect 18311 16896 18627 16897
rect 18311 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18627 16896
rect 18311 16831 18627 16832
rect 25257 16896 25573 16897
rect 25257 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25573 16896
rect 25257 16831 25573 16832
rect 28165 16826 28231 16829
rect 29200 16826 30000 16856
rect 28165 16824 30000 16826
rect 28165 16768 28170 16824
rect 28226 16768 30000 16824
rect 28165 16766 30000 16768
rect 28165 16763 28231 16766
rect 29200 16736 30000 16766
rect 7892 16352 8208 16353
rect 7892 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8208 16352
rect 7892 16287 8208 16288
rect 14838 16352 15154 16353
rect 14838 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15154 16352
rect 14838 16287 15154 16288
rect 21784 16352 22100 16353
rect 21784 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22100 16352
rect 21784 16287 22100 16288
rect 28730 16352 29046 16353
rect 28730 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29046 16352
rect 28730 16287 29046 16288
rect 4419 15808 4735 15809
rect 4419 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4735 15808
rect 4419 15743 4735 15744
rect 11365 15808 11681 15809
rect 11365 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11681 15808
rect 11365 15743 11681 15744
rect 18311 15808 18627 15809
rect 18311 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18627 15808
rect 18311 15743 18627 15744
rect 25257 15808 25573 15809
rect 25257 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25573 15808
rect 25257 15743 25573 15744
rect 7892 15264 8208 15265
rect 7892 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8208 15264
rect 7892 15199 8208 15200
rect 14838 15264 15154 15265
rect 14838 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15154 15264
rect 14838 15199 15154 15200
rect 21784 15264 22100 15265
rect 21784 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22100 15264
rect 21784 15199 22100 15200
rect 28730 15264 29046 15265
rect 28730 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29046 15264
rect 28730 15199 29046 15200
rect 4419 14720 4735 14721
rect 4419 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4735 14720
rect 4419 14655 4735 14656
rect 11365 14720 11681 14721
rect 11365 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11681 14720
rect 11365 14655 11681 14656
rect 18311 14720 18627 14721
rect 18311 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18627 14720
rect 18311 14655 18627 14656
rect 25257 14720 25573 14721
rect 25257 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25573 14720
rect 25257 14655 25573 14656
rect 7892 14176 8208 14177
rect 7892 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8208 14176
rect 7892 14111 8208 14112
rect 14838 14176 15154 14177
rect 14838 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15154 14176
rect 14838 14111 15154 14112
rect 21784 14176 22100 14177
rect 21784 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22100 14176
rect 21784 14111 22100 14112
rect 28730 14176 29046 14177
rect 28730 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29046 14176
rect 28730 14111 29046 14112
rect 4419 13632 4735 13633
rect 4419 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4735 13632
rect 4419 13567 4735 13568
rect 11365 13632 11681 13633
rect 11365 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11681 13632
rect 11365 13567 11681 13568
rect 18311 13632 18627 13633
rect 18311 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18627 13632
rect 18311 13567 18627 13568
rect 25257 13632 25573 13633
rect 25257 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25573 13632
rect 25257 13567 25573 13568
rect 28165 13290 28231 13293
rect 28165 13288 29194 13290
rect 28165 13232 28170 13288
rect 28226 13232 29194 13288
rect 28165 13230 29194 13232
rect 28165 13227 28231 13230
rect 29134 13188 29194 13230
rect 29134 13184 29378 13188
rect 29134 13128 30000 13184
rect 7892 13088 8208 13089
rect 7892 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8208 13088
rect 7892 13023 8208 13024
rect 14838 13088 15154 13089
rect 14838 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15154 13088
rect 14838 13023 15154 13024
rect 21784 13088 22100 13089
rect 21784 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22100 13088
rect 21784 13023 22100 13024
rect 28730 13088 29046 13089
rect 28730 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29046 13088
rect 29200 13064 30000 13128
rect 28730 13023 29046 13024
rect 4419 12544 4735 12545
rect 4419 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4735 12544
rect 4419 12479 4735 12480
rect 11365 12544 11681 12545
rect 11365 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11681 12544
rect 11365 12479 11681 12480
rect 18311 12544 18627 12545
rect 18311 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18627 12544
rect 18311 12479 18627 12480
rect 25257 12544 25573 12545
rect 25257 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25573 12544
rect 25257 12479 25573 12480
rect 7892 12000 8208 12001
rect 7892 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8208 12000
rect 7892 11935 8208 11936
rect 14838 12000 15154 12001
rect 14838 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15154 12000
rect 14838 11935 15154 11936
rect 21784 12000 22100 12001
rect 21784 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22100 12000
rect 21784 11935 22100 11936
rect 28730 12000 29046 12001
rect 28730 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29046 12000
rect 28730 11935 29046 11936
rect 4419 11456 4735 11457
rect 4419 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4735 11456
rect 4419 11391 4735 11392
rect 11365 11456 11681 11457
rect 11365 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11681 11456
rect 11365 11391 11681 11392
rect 18311 11456 18627 11457
rect 18311 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18627 11456
rect 18311 11391 18627 11392
rect 25257 11456 25573 11457
rect 25257 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25573 11456
rect 25257 11391 25573 11392
rect 7892 10912 8208 10913
rect 7892 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8208 10912
rect 7892 10847 8208 10848
rect 14838 10912 15154 10913
rect 14838 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15154 10912
rect 14838 10847 15154 10848
rect 21784 10912 22100 10913
rect 21784 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22100 10912
rect 21784 10847 22100 10848
rect 28730 10912 29046 10913
rect 28730 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29046 10912
rect 28730 10847 29046 10848
rect 4419 10368 4735 10369
rect 4419 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4735 10368
rect 4419 10303 4735 10304
rect 11365 10368 11681 10369
rect 11365 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11681 10368
rect 11365 10303 11681 10304
rect 18311 10368 18627 10369
rect 18311 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18627 10368
rect 18311 10303 18627 10304
rect 25257 10368 25573 10369
rect 25257 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25573 10368
rect 25257 10303 25573 10304
rect 7892 9824 8208 9825
rect 7892 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8208 9824
rect 7892 9759 8208 9760
rect 14838 9824 15154 9825
rect 14838 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15154 9824
rect 14838 9759 15154 9760
rect 21784 9824 22100 9825
rect 21784 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22100 9824
rect 21784 9759 22100 9760
rect 28730 9824 29046 9825
rect 28730 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29046 9824
rect 28730 9759 29046 9760
rect 28165 9482 28231 9485
rect 29200 9482 30000 9512
rect 28165 9480 30000 9482
rect 28165 9424 28170 9480
rect 28226 9424 30000 9480
rect 28165 9422 30000 9424
rect 28165 9419 28231 9422
rect 29200 9392 30000 9422
rect 4419 9280 4735 9281
rect 4419 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4735 9280
rect 4419 9215 4735 9216
rect 11365 9280 11681 9281
rect 11365 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11681 9280
rect 11365 9215 11681 9216
rect 18311 9280 18627 9281
rect 18311 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18627 9280
rect 18311 9215 18627 9216
rect 25257 9280 25573 9281
rect 25257 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25573 9280
rect 25257 9215 25573 9216
rect 7892 8736 8208 8737
rect 7892 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8208 8736
rect 7892 8671 8208 8672
rect 14838 8736 15154 8737
rect 14838 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15154 8736
rect 14838 8671 15154 8672
rect 21784 8736 22100 8737
rect 21784 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22100 8736
rect 21784 8671 22100 8672
rect 28730 8736 29046 8737
rect 28730 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29046 8736
rect 28730 8671 29046 8672
rect 4419 8192 4735 8193
rect 4419 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4735 8192
rect 4419 8127 4735 8128
rect 11365 8192 11681 8193
rect 11365 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11681 8192
rect 11365 8127 11681 8128
rect 18311 8192 18627 8193
rect 18311 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18627 8192
rect 18311 8127 18627 8128
rect 25257 8192 25573 8193
rect 25257 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25573 8192
rect 25257 8127 25573 8128
rect 26417 7714 26483 7717
rect 27613 7714 27679 7717
rect 26417 7712 27679 7714
rect 26417 7656 26422 7712
rect 26478 7656 27618 7712
rect 27674 7656 27679 7712
rect 26417 7654 27679 7656
rect 26417 7651 26483 7654
rect 27613 7651 27679 7654
rect 7892 7648 8208 7649
rect 7892 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8208 7648
rect 7892 7583 8208 7584
rect 14838 7648 15154 7649
rect 14838 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15154 7648
rect 14838 7583 15154 7584
rect 21784 7648 22100 7649
rect 21784 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22100 7648
rect 21784 7583 22100 7584
rect 28730 7648 29046 7649
rect 28730 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29046 7648
rect 28730 7583 29046 7584
rect 4419 7104 4735 7105
rect 4419 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4735 7104
rect 4419 7039 4735 7040
rect 11365 7104 11681 7105
rect 11365 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11681 7104
rect 11365 7039 11681 7040
rect 18311 7104 18627 7105
rect 18311 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18627 7104
rect 18311 7039 18627 7040
rect 25257 7104 25573 7105
rect 25257 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25573 7104
rect 25257 7039 25573 7040
rect 7892 6560 8208 6561
rect 7892 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8208 6560
rect 7892 6495 8208 6496
rect 14838 6560 15154 6561
rect 14838 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15154 6560
rect 14838 6495 15154 6496
rect 21784 6560 22100 6561
rect 21784 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22100 6560
rect 21784 6495 22100 6496
rect 28730 6560 29046 6561
rect 28730 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29046 6560
rect 28730 6495 29046 6496
rect 4419 6016 4735 6017
rect 4419 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4735 6016
rect 4419 5951 4735 5952
rect 11365 6016 11681 6017
rect 11365 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11681 6016
rect 11365 5951 11681 5952
rect 18311 6016 18627 6017
rect 18311 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18627 6016
rect 18311 5951 18627 5952
rect 25257 6016 25573 6017
rect 25257 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25573 6016
rect 25257 5951 25573 5952
rect 28165 5810 28231 5813
rect 29200 5810 30000 5840
rect 28165 5808 30000 5810
rect 28165 5752 28170 5808
rect 28226 5752 30000 5808
rect 28165 5750 30000 5752
rect 28165 5747 28231 5750
rect 29200 5720 30000 5750
rect 7892 5472 8208 5473
rect 7892 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8208 5472
rect 7892 5407 8208 5408
rect 14838 5472 15154 5473
rect 14838 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15154 5472
rect 14838 5407 15154 5408
rect 21784 5472 22100 5473
rect 21784 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22100 5472
rect 21784 5407 22100 5408
rect 28730 5472 29046 5473
rect 28730 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29046 5472
rect 28730 5407 29046 5408
rect 4419 4928 4735 4929
rect 4419 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4735 4928
rect 4419 4863 4735 4864
rect 11365 4928 11681 4929
rect 11365 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11681 4928
rect 11365 4863 11681 4864
rect 18311 4928 18627 4929
rect 18311 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18627 4928
rect 18311 4863 18627 4864
rect 25257 4928 25573 4929
rect 25257 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25573 4928
rect 25257 4863 25573 4864
rect 7892 4384 8208 4385
rect 7892 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8208 4384
rect 7892 4319 8208 4320
rect 14838 4384 15154 4385
rect 14838 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15154 4384
rect 14838 4319 15154 4320
rect 21784 4384 22100 4385
rect 21784 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22100 4384
rect 21784 4319 22100 4320
rect 28730 4384 29046 4385
rect 28730 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29046 4384
rect 28730 4319 29046 4320
rect 4419 3840 4735 3841
rect 4419 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4735 3840
rect 4419 3775 4735 3776
rect 11365 3840 11681 3841
rect 11365 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11681 3840
rect 11365 3775 11681 3776
rect 18311 3840 18627 3841
rect 18311 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18627 3840
rect 18311 3775 18627 3776
rect 25257 3840 25573 3841
rect 25257 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25573 3840
rect 25257 3775 25573 3776
rect 7892 3296 8208 3297
rect 7892 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8208 3296
rect 7892 3231 8208 3232
rect 14838 3296 15154 3297
rect 14838 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15154 3296
rect 14838 3231 15154 3232
rect 21784 3296 22100 3297
rect 21784 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22100 3296
rect 21784 3231 22100 3232
rect 28730 3296 29046 3297
rect 28730 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29046 3296
rect 28730 3231 29046 3232
rect 4419 2752 4735 2753
rect 4419 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4735 2752
rect 4419 2687 4735 2688
rect 11365 2752 11681 2753
rect 11365 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11681 2752
rect 11365 2687 11681 2688
rect 18311 2752 18627 2753
rect 18311 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18627 2752
rect 18311 2687 18627 2688
rect 25257 2752 25573 2753
rect 25257 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25573 2752
rect 25257 2687 25573 2688
rect 28165 2410 28231 2413
rect 28165 2408 29378 2410
rect 28165 2352 28170 2408
rect 28226 2352 29378 2408
rect 28165 2350 29378 2352
rect 28165 2347 28231 2350
rect 7892 2208 8208 2209
rect 7892 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8208 2208
rect 7892 2143 8208 2144
rect 14838 2208 15154 2209
rect 14838 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15154 2208
rect 14838 2143 15154 2144
rect 21784 2208 22100 2209
rect 21784 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22100 2208
rect 21784 2143 22100 2144
rect 28730 2208 29046 2209
rect 28730 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29046 2208
rect 29318 2168 29378 2350
rect 28730 2143 29046 2144
rect 29200 2048 30000 2168
<< via3 >>
rect 4425 27772 4489 27776
rect 4425 27716 4429 27772
rect 4429 27716 4485 27772
rect 4485 27716 4489 27772
rect 4425 27712 4489 27716
rect 4505 27772 4569 27776
rect 4505 27716 4509 27772
rect 4509 27716 4565 27772
rect 4565 27716 4569 27772
rect 4505 27712 4569 27716
rect 4585 27772 4649 27776
rect 4585 27716 4589 27772
rect 4589 27716 4645 27772
rect 4645 27716 4649 27772
rect 4585 27712 4649 27716
rect 4665 27772 4729 27776
rect 4665 27716 4669 27772
rect 4669 27716 4725 27772
rect 4725 27716 4729 27772
rect 4665 27712 4729 27716
rect 11371 27772 11435 27776
rect 11371 27716 11375 27772
rect 11375 27716 11431 27772
rect 11431 27716 11435 27772
rect 11371 27712 11435 27716
rect 11451 27772 11515 27776
rect 11451 27716 11455 27772
rect 11455 27716 11511 27772
rect 11511 27716 11515 27772
rect 11451 27712 11515 27716
rect 11531 27772 11595 27776
rect 11531 27716 11535 27772
rect 11535 27716 11591 27772
rect 11591 27716 11595 27772
rect 11531 27712 11595 27716
rect 11611 27772 11675 27776
rect 11611 27716 11615 27772
rect 11615 27716 11671 27772
rect 11671 27716 11675 27772
rect 11611 27712 11675 27716
rect 18317 27772 18381 27776
rect 18317 27716 18321 27772
rect 18321 27716 18377 27772
rect 18377 27716 18381 27772
rect 18317 27712 18381 27716
rect 18397 27772 18461 27776
rect 18397 27716 18401 27772
rect 18401 27716 18457 27772
rect 18457 27716 18461 27772
rect 18397 27712 18461 27716
rect 18477 27772 18541 27776
rect 18477 27716 18481 27772
rect 18481 27716 18537 27772
rect 18537 27716 18541 27772
rect 18477 27712 18541 27716
rect 18557 27772 18621 27776
rect 18557 27716 18561 27772
rect 18561 27716 18617 27772
rect 18617 27716 18621 27772
rect 18557 27712 18621 27716
rect 25263 27772 25327 27776
rect 25263 27716 25267 27772
rect 25267 27716 25323 27772
rect 25323 27716 25327 27772
rect 25263 27712 25327 27716
rect 25343 27772 25407 27776
rect 25343 27716 25347 27772
rect 25347 27716 25403 27772
rect 25403 27716 25407 27772
rect 25343 27712 25407 27716
rect 25423 27772 25487 27776
rect 25423 27716 25427 27772
rect 25427 27716 25483 27772
rect 25483 27716 25487 27772
rect 25423 27712 25487 27716
rect 25503 27772 25567 27776
rect 25503 27716 25507 27772
rect 25507 27716 25563 27772
rect 25563 27716 25567 27772
rect 25503 27712 25567 27716
rect 7898 27228 7962 27232
rect 7898 27172 7902 27228
rect 7902 27172 7958 27228
rect 7958 27172 7962 27228
rect 7898 27168 7962 27172
rect 7978 27228 8042 27232
rect 7978 27172 7982 27228
rect 7982 27172 8038 27228
rect 8038 27172 8042 27228
rect 7978 27168 8042 27172
rect 8058 27228 8122 27232
rect 8058 27172 8062 27228
rect 8062 27172 8118 27228
rect 8118 27172 8122 27228
rect 8058 27168 8122 27172
rect 8138 27228 8202 27232
rect 8138 27172 8142 27228
rect 8142 27172 8198 27228
rect 8198 27172 8202 27228
rect 8138 27168 8202 27172
rect 14844 27228 14908 27232
rect 14844 27172 14848 27228
rect 14848 27172 14904 27228
rect 14904 27172 14908 27228
rect 14844 27168 14908 27172
rect 14924 27228 14988 27232
rect 14924 27172 14928 27228
rect 14928 27172 14984 27228
rect 14984 27172 14988 27228
rect 14924 27168 14988 27172
rect 15004 27228 15068 27232
rect 15004 27172 15008 27228
rect 15008 27172 15064 27228
rect 15064 27172 15068 27228
rect 15004 27168 15068 27172
rect 15084 27228 15148 27232
rect 15084 27172 15088 27228
rect 15088 27172 15144 27228
rect 15144 27172 15148 27228
rect 15084 27168 15148 27172
rect 21790 27228 21854 27232
rect 21790 27172 21794 27228
rect 21794 27172 21850 27228
rect 21850 27172 21854 27228
rect 21790 27168 21854 27172
rect 21870 27228 21934 27232
rect 21870 27172 21874 27228
rect 21874 27172 21930 27228
rect 21930 27172 21934 27228
rect 21870 27168 21934 27172
rect 21950 27228 22014 27232
rect 21950 27172 21954 27228
rect 21954 27172 22010 27228
rect 22010 27172 22014 27228
rect 21950 27168 22014 27172
rect 22030 27228 22094 27232
rect 22030 27172 22034 27228
rect 22034 27172 22090 27228
rect 22090 27172 22094 27228
rect 22030 27168 22094 27172
rect 28736 27228 28800 27232
rect 28736 27172 28740 27228
rect 28740 27172 28796 27228
rect 28796 27172 28800 27228
rect 28736 27168 28800 27172
rect 28816 27228 28880 27232
rect 28816 27172 28820 27228
rect 28820 27172 28876 27228
rect 28876 27172 28880 27228
rect 28816 27168 28880 27172
rect 28896 27228 28960 27232
rect 28896 27172 28900 27228
rect 28900 27172 28956 27228
rect 28956 27172 28960 27228
rect 28896 27168 28960 27172
rect 28976 27228 29040 27232
rect 28976 27172 28980 27228
rect 28980 27172 29036 27228
rect 29036 27172 29040 27228
rect 28976 27168 29040 27172
rect 4425 26684 4489 26688
rect 4425 26628 4429 26684
rect 4429 26628 4485 26684
rect 4485 26628 4489 26684
rect 4425 26624 4489 26628
rect 4505 26684 4569 26688
rect 4505 26628 4509 26684
rect 4509 26628 4565 26684
rect 4565 26628 4569 26684
rect 4505 26624 4569 26628
rect 4585 26684 4649 26688
rect 4585 26628 4589 26684
rect 4589 26628 4645 26684
rect 4645 26628 4649 26684
rect 4585 26624 4649 26628
rect 4665 26684 4729 26688
rect 4665 26628 4669 26684
rect 4669 26628 4725 26684
rect 4725 26628 4729 26684
rect 4665 26624 4729 26628
rect 11371 26684 11435 26688
rect 11371 26628 11375 26684
rect 11375 26628 11431 26684
rect 11431 26628 11435 26684
rect 11371 26624 11435 26628
rect 11451 26684 11515 26688
rect 11451 26628 11455 26684
rect 11455 26628 11511 26684
rect 11511 26628 11515 26684
rect 11451 26624 11515 26628
rect 11531 26684 11595 26688
rect 11531 26628 11535 26684
rect 11535 26628 11591 26684
rect 11591 26628 11595 26684
rect 11531 26624 11595 26628
rect 11611 26684 11675 26688
rect 11611 26628 11615 26684
rect 11615 26628 11671 26684
rect 11671 26628 11675 26684
rect 11611 26624 11675 26628
rect 18317 26684 18381 26688
rect 18317 26628 18321 26684
rect 18321 26628 18377 26684
rect 18377 26628 18381 26684
rect 18317 26624 18381 26628
rect 18397 26684 18461 26688
rect 18397 26628 18401 26684
rect 18401 26628 18457 26684
rect 18457 26628 18461 26684
rect 18397 26624 18461 26628
rect 18477 26684 18541 26688
rect 18477 26628 18481 26684
rect 18481 26628 18537 26684
rect 18537 26628 18541 26684
rect 18477 26624 18541 26628
rect 18557 26684 18621 26688
rect 18557 26628 18561 26684
rect 18561 26628 18617 26684
rect 18617 26628 18621 26684
rect 18557 26624 18621 26628
rect 25263 26684 25327 26688
rect 25263 26628 25267 26684
rect 25267 26628 25323 26684
rect 25323 26628 25327 26684
rect 25263 26624 25327 26628
rect 25343 26684 25407 26688
rect 25343 26628 25347 26684
rect 25347 26628 25403 26684
rect 25403 26628 25407 26684
rect 25343 26624 25407 26628
rect 25423 26684 25487 26688
rect 25423 26628 25427 26684
rect 25427 26628 25483 26684
rect 25483 26628 25487 26684
rect 25423 26624 25487 26628
rect 25503 26684 25567 26688
rect 25503 26628 25507 26684
rect 25507 26628 25563 26684
rect 25563 26628 25567 26684
rect 25503 26624 25567 26628
rect 7898 26140 7962 26144
rect 7898 26084 7902 26140
rect 7902 26084 7958 26140
rect 7958 26084 7962 26140
rect 7898 26080 7962 26084
rect 7978 26140 8042 26144
rect 7978 26084 7982 26140
rect 7982 26084 8038 26140
rect 8038 26084 8042 26140
rect 7978 26080 8042 26084
rect 8058 26140 8122 26144
rect 8058 26084 8062 26140
rect 8062 26084 8118 26140
rect 8118 26084 8122 26140
rect 8058 26080 8122 26084
rect 8138 26140 8202 26144
rect 8138 26084 8142 26140
rect 8142 26084 8198 26140
rect 8198 26084 8202 26140
rect 8138 26080 8202 26084
rect 14844 26140 14908 26144
rect 14844 26084 14848 26140
rect 14848 26084 14904 26140
rect 14904 26084 14908 26140
rect 14844 26080 14908 26084
rect 14924 26140 14988 26144
rect 14924 26084 14928 26140
rect 14928 26084 14984 26140
rect 14984 26084 14988 26140
rect 14924 26080 14988 26084
rect 15004 26140 15068 26144
rect 15004 26084 15008 26140
rect 15008 26084 15064 26140
rect 15064 26084 15068 26140
rect 15004 26080 15068 26084
rect 15084 26140 15148 26144
rect 15084 26084 15088 26140
rect 15088 26084 15144 26140
rect 15144 26084 15148 26140
rect 15084 26080 15148 26084
rect 21790 26140 21854 26144
rect 21790 26084 21794 26140
rect 21794 26084 21850 26140
rect 21850 26084 21854 26140
rect 21790 26080 21854 26084
rect 21870 26140 21934 26144
rect 21870 26084 21874 26140
rect 21874 26084 21930 26140
rect 21930 26084 21934 26140
rect 21870 26080 21934 26084
rect 21950 26140 22014 26144
rect 21950 26084 21954 26140
rect 21954 26084 22010 26140
rect 22010 26084 22014 26140
rect 21950 26080 22014 26084
rect 22030 26140 22094 26144
rect 22030 26084 22034 26140
rect 22034 26084 22090 26140
rect 22090 26084 22094 26140
rect 22030 26080 22094 26084
rect 28736 26140 28800 26144
rect 28736 26084 28740 26140
rect 28740 26084 28796 26140
rect 28796 26084 28800 26140
rect 28736 26080 28800 26084
rect 28816 26140 28880 26144
rect 28816 26084 28820 26140
rect 28820 26084 28876 26140
rect 28876 26084 28880 26140
rect 28816 26080 28880 26084
rect 28896 26140 28960 26144
rect 28896 26084 28900 26140
rect 28900 26084 28956 26140
rect 28956 26084 28960 26140
rect 28896 26080 28960 26084
rect 28976 26140 29040 26144
rect 28976 26084 28980 26140
rect 28980 26084 29036 26140
rect 29036 26084 29040 26140
rect 28976 26080 29040 26084
rect 4425 25596 4489 25600
rect 4425 25540 4429 25596
rect 4429 25540 4485 25596
rect 4485 25540 4489 25596
rect 4425 25536 4489 25540
rect 4505 25596 4569 25600
rect 4505 25540 4509 25596
rect 4509 25540 4565 25596
rect 4565 25540 4569 25596
rect 4505 25536 4569 25540
rect 4585 25596 4649 25600
rect 4585 25540 4589 25596
rect 4589 25540 4645 25596
rect 4645 25540 4649 25596
rect 4585 25536 4649 25540
rect 4665 25596 4729 25600
rect 4665 25540 4669 25596
rect 4669 25540 4725 25596
rect 4725 25540 4729 25596
rect 4665 25536 4729 25540
rect 11371 25596 11435 25600
rect 11371 25540 11375 25596
rect 11375 25540 11431 25596
rect 11431 25540 11435 25596
rect 11371 25536 11435 25540
rect 11451 25596 11515 25600
rect 11451 25540 11455 25596
rect 11455 25540 11511 25596
rect 11511 25540 11515 25596
rect 11451 25536 11515 25540
rect 11531 25596 11595 25600
rect 11531 25540 11535 25596
rect 11535 25540 11591 25596
rect 11591 25540 11595 25596
rect 11531 25536 11595 25540
rect 11611 25596 11675 25600
rect 11611 25540 11615 25596
rect 11615 25540 11671 25596
rect 11671 25540 11675 25596
rect 11611 25536 11675 25540
rect 18317 25596 18381 25600
rect 18317 25540 18321 25596
rect 18321 25540 18377 25596
rect 18377 25540 18381 25596
rect 18317 25536 18381 25540
rect 18397 25596 18461 25600
rect 18397 25540 18401 25596
rect 18401 25540 18457 25596
rect 18457 25540 18461 25596
rect 18397 25536 18461 25540
rect 18477 25596 18541 25600
rect 18477 25540 18481 25596
rect 18481 25540 18537 25596
rect 18537 25540 18541 25596
rect 18477 25536 18541 25540
rect 18557 25596 18621 25600
rect 18557 25540 18561 25596
rect 18561 25540 18617 25596
rect 18617 25540 18621 25596
rect 18557 25536 18621 25540
rect 25263 25596 25327 25600
rect 25263 25540 25267 25596
rect 25267 25540 25323 25596
rect 25323 25540 25327 25596
rect 25263 25536 25327 25540
rect 25343 25596 25407 25600
rect 25343 25540 25347 25596
rect 25347 25540 25403 25596
rect 25403 25540 25407 25596
rect 25343 25536 25407 25540
rect 25423 25596 25487 25600
rect 25423 25540 25427 25596
rect 25427 25540 25483 25596
rect 25483 25540 25487 25596
rect 25423 25536 25487 25540
rect 25503 25596 25567 25600
rect 25503 25540 25507 25596
rect 25507 25540 25563 25596
rect 25563 25540 25567 25596
rect 25503 25536 25567 25540
rect 7898 25052 7962 25056
rect 7898 24996 7902 25052
rect 7902 24996 7958 25052
rect 7958 24996 7962 25052
rect 7898 24992 7962 24996
rect 7978 25052 8042 25056
rect 7978 24996 7982 25052
rect 7982 24996 8038 25052
rect 8038 24996 8042 25052
rect 7978 24992 8042 24996
rect 8058 25052 8122 25056
rect 8058 24996 8062 25052
rect 8062 24996 8118 25052
rect 8118 24996 8122 25052
rect 8058 24992 8122 24996
rect 8138 25052 8202 25056
rect 8138 24996 8142 25052
rect 8142 24996 8198 25052
rect 8198 24996 8202 25052
rect 8138 24992 8202 24996
rect 14844 25052 14908 25056
rect 14844 24996 14848 25052
rect 14848 24996 14904 25052
rect 14904 24996 14908 25052
rect 14844 24992 14908 24996
rect 14924 25052 14988 25056
rect 14924 24996 14928 25052
rect 14928 24996 14984 25052
rect 14984 24996 14988 25052
rect 14924 24992 14988 24996
rect 15004 25052 15068 25056
rect 15004 24996 15008 25052
rect 15008 24996 15064 25052
rect 15064 24996 15068 25052
rect 15004 24992 15068 24996
rect 15084 25052 15148 25056
rect 15084 24996 15088 25052
rect 15088 24996 15144 25052
rect 15144 24996 15148 25052
rect 15084 24992 15148 24996
rect 21790 25052 21854 25056
rect 21790 24996 21794 25052
rect 21794 24996 21850 25052
rect 21850 24996 21854 25052
rect 21790 24992 21854 24996
rect 21870 25052 21934 25056
rect 21870 24996 21874 25052
rect 21874 24996 21930 25052
rect 21930 24996 21934 25052
rect 21870 24992 21934 24996
rect 21950 25052 22014 25056
rect 21950 24996 21954 25052
rect 21954 24996 22010 25052
rect 22010 24996 22014 25052
rect 21950 24992 22014 24996
rect 22030 25052 22094 25056
rect 22030 24996 22034 25052
rect 22034 24996 22090 25052
rect 22090 24996 22094 25052
rect 22030 24992 22094 24996
rect 28736 25052 28800 25056
rect 28736 24996 28740 25052
rect 28740 24996 28796 25052
rect 28796 24996 28800 25052
rect 28736 24992 28800 24996
rect 28816 25052 28880 25056
rect 28816 24996 28820 25052
rect 28820 24996 28876 25052
rect 28876 24996 28880 25052
rect 28816 24992 28880 24996
rect 28896 25052 28960 25056
rect 28896 24996 28900 25052
rect 28900 24996 28956 25052
rect 28956 24996 28960 25052
rect 28896 24992 28960 24996
rect 28976 25052 29040 25056
rect 28976 24996 28980 25052
rect 28980 24996 29036 25052
rect 29036 24996 29040 25052
rect 28976 24992 29040 24996
rect 4425 24508 4489 24512
rect 4425 24452 4429 24508
rect 4429 24452 4485 24508
rect 4485 24452 4489 24508
rect 4425 24448 4489 24452
rect 4505 24508 4569 24512
rect 4505 24452 4509 24508
rect 4509 24452 4565 24508
rect 4565 24452 4569 24508
rect 4505 24448 4569 24452
rect 4585 24508 4649 24512
rect 4585 24452 4589 24508
rect 4589 24452 4645 24508
rect 4645 24452 4649 24508
rect 4585 24448 4649 24452
rect 4665 24508 4729 24512
rect 4665 24452 4669 24508
rect 4669 24452 4725 24508
rect 4725 24452 4729 24508
rect 4665 24448 4729 24452
rect 11371 24508 11435 24512
rect 11371 24452 11375 24508
rect 11375 24452 11431 24508
rect 11431 24452 11435 24508
rect 11371 24448 11435 24452
rect 11451 24508 11515 24512
rect 11451 24452 11455 24508
rect 11455 24452 11511 24508
rect 11511 24452 11515 24508
rect 11451 24448 11515 24452
rect 11531 24508 11595 24512
rect 11531 24452 11535 24508
rect 11535 24452 11591 24508
rect 11591 24452 11595 24508
rect 11531 24448 11595 24452
rect 11611 24508 11675 24512
rect 11611 24452 11615 24508
rect 11615 24452 11671 24508
rect 11671 24452 11675 24508
rect 11611 24448 11675 24452
rect 18317 24508 18381 24512
rect 18317 24452 18321 24508
rect 18321 24452 18377 24508
rect 18377 24452 18381 24508
rect 18317 24448 18381 24452
rect 18397 24508 18461 24512
rect 18397 24452 18401 24508
rect 18401 24452 18457 24508
rect 18457 24452 18461 24508
rect 18397 24448 18461 24452
rect 18477 24508 18541 24512
rect 18477 24452 18481 24508
rect 18481 24452 18537 24508
rect 18537 24452 18541 24508
rect 18477 24448 18541 24452
rect 18557 24508 18621 24512
rect 18557 24452 18561 24508
rect 18561 24452 18617 24508
rect 18617 24452 18621 24508
rect 18557 24448 18621 24452
rect 25263 24508 25327 24512
rect 25263 24452 25267 24508
rect 25267 24452 25323 24508
rect 25323 24452 25327 24508
rect 25263 24448 25327 24452
rect 25343 24508 25407 24512
rect 25343 24452 25347 24508
rect 25347 24452 25403 24508
rect 25403 24452 25407 24508
rect 25343 24448 25407 24452
rect 25423 24508 25487 24512
rect 25423 24452 25427 24508
rect 25427 24452 25483 24508
rect 25483 24452 25487 24508
rect 25423 24448 25487 24452
rect 25503 24508 25567 24512
rect 25503 24452 25507 24508
rect 25507 24452 25563 24508
rect 25563 24452 25567 24508
rect 25503 24448 25567 24452
rect 7898 23964 7962 23968
rect 7898 23908 7902 23964
rect 7902 23908 7958 23964
rect 7958 23908 7962 23964
rect 7898 23904 7962 23908
rect 7978 23964 8042 23968
rect 7978 23908 7982 23964
rect 7982 23908 8038 23964
rect 8038 23908 8042 23964
rect 7978 23904 8042 23908
rect 8058 23964 8122 23968
rect 8058 23908 8062 23964
rect 8062 23908 8118 23964
rect 8118 23908 8122 23964
rect 8058 23904 8122 23908
rect 8138 23964 8202 23968
rect 8138 23908 8142 23964
rect 8142 23908 8198 23964
rect 8198 23908 8202 23964
rect 8138 23904 8202 23908
rect 14844 23964 14908 23968
rect 14844 23908 14848 23964
rect 14848 23908 14904 23964
rect 14904 23908 14908 23964
rect 14844 23904 14908 23908
rect 14924 23964 14988 23968
rect 14924 23908 14928 23964
rect 14928 23908 14984 23964
rect 14984 23908 14988 23964
rect 14924 23904 14988 23908
rect 15004 23964 15068 23968
rect 15004 23908 15008 23964
rect 15008 23908 15064 23964
rect 15064 23908 15068 23964
rect 15004 23904 15068 23908
rect 15084 23964 15148 23968
rect 15084 23908 15088 23964
rect 15088 23908 15144 23964
rect 15144 23908 15148 23964
rect 15084 23904 15148 23908
rect 21790 23964 21854 23968
rect 21790 23908 21794 23964
rect 21794 23908 21850 23964
rect 21850 23908 21854 23964
rect 21790 23904 21854 23908
rect 21870 23964 21934 23968
rect 21870 23908 21874 23964
rect 21874 23908 21930 23964
rect 21930 23908 21934 23964
rect 21870 23904 21934 23908
rect 21950 23964 22014 23968
rect 21950 23908 21954 23964
rect 21954 23908 22010 23964
rect 22010 23908 22014 23964
rect 21950 23904 22014 23908
rect 22030 23964 22094 23968
rect 22030 23908 22034 23964
rect 22034 23908 22090 23964
rect 22090 23908 22094 23964
rect 22030 23904 22094 23908
rect 28736 23964 28800 23968
rect 28736 23908 28740 23964
rect 28740 23908 28796 23964
rect 28796 23908 28800 23964
rect 28736 23904 28800 23908
rect 28816 23964 28880 23968
rect 28816 23908 28820 23964
rect 28820 23908 28876 23964
rect 28876 23908 28880 23964
rect 28816 23904 28880 23908
rect 28896 23964 28960 23968
rect 28896 23908 28900 23964
rect 28900 23908 28956 23964
rect 28956 23908 28960 23964
rect 28896 23904 28960 23908
rect 28976 23964 29040 23968
rect 28976 23908 28980 23964
rect 28980 23908 29036 23964
rect 29036 23908 29040 23964
rect 28976 23904 29040 23908
rect 4425 23420 4489 23424
rect 4425 23364 4429 23420
rect 4429 23364 4485 23420
rect 4485 23364 4489 23420
rect 4425 23360 4489 23364
rect 4505 23420 4569 23424
rect 4505 23364 4509 23420
rect 4509 23364 4565 23420
rect 4565 23364 4569 23420
rect 4505 23360 4569 23364
rect 4585 23420 4649 23424
rect 4585 23364 4589 23420
rect 4589 23364 4645 23420
rect 4645 23364 4649 23420
rect 4585 23360 4649 23364
rect 4665 23420 4729 23424
rect 4665 23364 4669 23420
rect 4669 23364 4725 23420
rect 4725 23364 4729 23420
rect 4665 23360 4729 23364
rect 11371 23420 11435 23424
rect 11371 23364 11375 23420
rect 11375 23364 11431 23420
rect 11431 23364 11435 23420
rect 11371 23360 11435 23364
rect 11451 23420 11515 23424
rect 11451 23364 11455 23420
rect 11455 23364 11511 23420
rect 11511 23364 11515 23420
rect 11451 23360 11515 23364
rect 11531 23420 11595 23424
rect 11531 23364 11535 23420
rect 11535 23364 11591 23420
rect 11591 23364 11595 23420
rect 11531 23360 11595 23364
rect 11611 23420 11675 23424
rect 11611 23364 11615 23420
rect 11615 23364 11671 23420
rect 11671 23364 11675 23420
rect 11611 23360 11675 23364
rect 18317 23420 18381 23424
rect 18317 23364 18321 23420
rect 18321 23364 18377 23420
rect 18377 23364 18381 23420
rect 18317 23360 18381 23364
rect 18397 23420 18461 23424
rect 18397 23364 18401 23420
rect 18401 23364 18457 23420
rect 18457 23364 18461 23420
rect 18397 23360 18461 23364
rect 18477 23420 18541 23424
rect 18477 23364 18481 23420
rect 18481 23364 18537 23420
rect 18537 23364 18541 23420
rect 18477 23360 18541 23364
rect 18557 23420 18621 23424
rect 18557 23364 18561 23420
rect 18561 23364 18617 23420
rect 18617 23364 18621 23420
rect 18557 23360 18621 23364
rect 25263 23420 25327 23424
rect 25263 23364 25267 23420
rect 25267 23364 25323 23420
rect 25323 23364 25327 23420
rect 25263 23360 25327 23364
rect 25343 23420 25407 23424
rect 25343 23364 25347 23420
rect 25347 23364 25403 23420
rect 25403 23364 25407 23420
rect 25343 23360 25407 23364
rect 25423 23420 25487 23424
rect 25423 23364 25427 23420
rect 25427 23364 25483 23420
rect 25483 23364 25487 23420
rect 25423 23360 25487 23364
rect 25503 23420 25567 23424
rect 25503 23364 25507 23420
rect 25507 23364 25563 23420
rect 25563 23364 25567 23420
rect 25503 23360 25567 23364
rect 7898 22876 7962 22880
rect 7898 22820 7902 22876
rect 7902 22820 7958 22876
rect 7958 22820 7962 22876
rect 7898 22816 7962 22820
rect 7978 22876 8042 22880
rect 7978 22820 7982 22876
rect 7982 22820 8038 22876
rect 8038 22820 8042 22876
rect 7978 22816 8042 22820
rect 8058 22876 8122 22880
rect 8058 22820 8062 22876
rect 8062 22820 8118 22876
rect 8118 22820 8122 22876
rect 8058 22816 8122 22820
rect 8138 22876 8202 22880
rect 8138 22820 8142 22876
rect 8142 22820 8198 22876
rect 8198 22820 8202 22876
rect 8138 22816 8202 22820
rect 14844 22876 14908 22880
rect 14844 22820 14848 22876
rect 14848 22820 14904 22876
rect 14904 22820 14908 22876
rect 14844 22816 14908 22820
rect 14924 22876 14988 22880
rect 14924 22820 14928 22876
rect 14928 22820 14984 22876
rect 14984 22820 14988 22876
rect 14924 22816 14988 22820
rect 15004 22876 15068 22880
rect 15004 22820 15008 22876
rect 15008 22820 15064 22876
rect 15064 22820 15068 22876
rect 15004 22816 15068 22820
rect 15084 22876 15148 22880
rect 15084 22820 15088 22876
rect 15088 22820 15144 22876
rect 15144 22820 15148 22876
rect 15084 22816 15148 22820
rect 21790 22876 21854 22880
rect 21790 22820 21794 22876
rect 21794 22820 21850 22876
rect 21850 22820 21854 22876
rect 21790 22816 21854 22820
rect 21870 22876 21934 22880
rect 21870 22820 21874 22876
rect 21874 22820 21930 22876
rect 21930 22820 21934 22876
rect 21870 22816 21934 22820
rect 21950 22876 22014 22880
rect 21950 22820 21954 22876
rect 21954 22820 22010 22876
rect 22010 22820 22014 22876
rect 21950 22816 22014 22820
rect 22030 22876 22094 22880
rect 22030 22820 22034 22876
rect 22034 22820 22090 22876
rect 22090 22820 22094 22876
rect 22030 22816 22094 22820
rect 28736 22876 28800 22880
rect 28736 22820 28740 22876
rect 28740 22820 28796 22876
rect 28796 22820 28800 22876
rect 28736 22816 28800 22820
rect 28816 22876 28880 22880
rect 28816 22820 28820 22876
rect 28820 22820 28876 22876
rect 28876 22820 28880 22876
rect 28816 22816 28880 22820
rect 28896 22876 28960 22880
rect 28896 22820 28900 22876
rect 28900 22820 28956 22876
rect 28956 22820 28960 22876
rect 28896 22816 28960 22820
rect 28976 22876 29040 22880
rect 28976 22820 28980 22876
rect 28980 22820 29036 22876
rect 29036 22820 29040 22876
rect 28976 22816 29040 22820
rect 4425 22332 4489 22336
rect 4425 22276 4429 22332
rect 4429 22276 4485 22332
rect 4485 22276 4489 22332
rect 4425 22272 4489 22276
rect 4505 22332 4569 22336
rect 4505 22276 4509 22332
rect 4509 22276 4565 22332
rect 4565 22276 4569 22332
rect 4505 22272 4569 22276
rect 4585 22332 4649 22336
rect 4585 22276 4589 22332
rect 4589 22276 4645 22332
rect 4645 22276 4649 22332
rect 4585 22272 4649 22276
rect 4665 22332 4729 22336
rect 4665 22276 4669 22332
rect 4669 22276 4725 22332
rect 4725 22276 4729 22332
rect 4665 22272 4729 22276
rect 11371 22332 11435 22336
rect 11371 22276 11375 22332
rect 11375 22276 11431 22332
rect 11431 22276 11435 22332
rect 11371 22272 11435 22276
rect 11451 22332 11515 22336
rect 11451 22276 11455 22332
rect 11455 22276 11511 22332
rect 11511 22276 11515 22332
rect 11451 22272 11515 22276
rect 11531 22332 11595 22336
rect 11531 22276 11535 22332
rect 11535 22276 11591 22332
rect 11591 22276 11595 22332
rect 11531 22272 11595 22276
rect 11611 22332 11675 22336
rect 11611 22276 11615 22332
rect 11615 22276 11671 22332
rect 11671 22276 11675 22332
rect 11611 22272 11675 22276
rect 18317 22332 18381 22336
rect 18317 22276 18321 22332
rect 18321 22276 18377 22332
rect 18377 22276 18381 22332
rect 18317 22272 18381 22276
rect 18397 22332 18461 22336
rect 18397 22276 18401 22332
rect 18401 22276 18457 22332
rect 18457 22276 18461 22332
rect 18397 22272 18461 22276
rect 18477 22332 18541 22336
rect 18477 22276 18481 22332
rect 18481 22276 18537 22332
rect 18537 22276 18541 22332
rect 18477 22272 18541 22276
rect 18557 22332 18621 22336
rect 18557 22276 18561 22332
rect 18561 22276 18617 22332
rect 18617 22276 18621 22332
rect 18557 22272 18621 22276
rect 25263 22332 25327 22336
rect 25263 22276 25267 22332
rect 25267 22276 25323 22332
rect 25323 22276 25327 22332
rect 25263 22272 25327 22276
rect 25343 22332 25407 22336
rect 25343 22276 25347 22332
rect 25347 22276 25403 22332
rect 25403 22276 25407 22332
rect 25343 22272 25407 22276
rect 25423 22332 25487 22336
rect 25423 22276 25427 22332
rect 25427 22276 25483 22332
rect 25483 22276 25487 22332
rect 25423 22272 25487 22276
rect 25503 22332 25567 22336
rect 25503 22276 25507 22332
rect 25507 22276 25563 22332
rect 25563 22276 25567 22332
rect 25503 22272 25567 22276
rect 7898 21788 7962 21792
rect 7898 21732 7902 21788
rect 7902 21732 7958 21788
rect 7958 21732 7962 21788
rect 7898 21728 7962 21732
rect 7978 21788 8042 21792
rect 7978 21732 7982 21788
rect 7982 21732 8038 21788
rect 8038 21732 8042 21788
rect 7978 21728 8042 21732
rect 8058 21788 8122 21792
rect 8058 21732 8062 21788
rect 8062 21732 8118 21788
rect 8118 21732 8122 21788
rect 8058 21728 8122 21732
rect 8138 21788 8202 21792
rect 8138 21732 8142 21788
rect 8142 21732 8198 21788
rect 8198 21732 8202 21788
rect 8138 21728 8202 21732
rect 14844 21788 14908 21792
rect 14844 21732 14848 21788
rect 14848 21732 14904 21788
rect 14904 21732 14908 21788
rect 14844 21728 14908 21732
rect 14924 21788 14988 21792
rect 14924 21732 14928 21788
rect 14928 21732 14984 21788
rect 14984 21732 14988 21788
rect 14924 21728 14988 21732
rect 15004 21788 15068 21792
rect 15004 21732 15008 21788
rect 15008 21732 15064 21788
rect 15064 21732 15068 21788
rect 15004 21728 15068 21732
rect 15084 21788 15148 21792
rect 15084 21732 15088 21788
rect 15088 21732 15144 21788
rect 15144 21732 15148 21788
rect 15084 21728 15148 21732
rect 21790 21788 21854 21792
rect 21790 21732 21794 21788
rect 21794 21732 21850 21788
rect 21850 21732 21854 21788
rect 21790 21728 21854 21732
rect 21870 21788 21934 21792
rect 21870 21732 21874 21788
rect 21874 21732 21930 21788
rect 21930 21732 21934 21788
rect 21870 21728 21934 21732
rect 21950 21788 22014 21792
rect 21950 21732 21954 21788
rect 21954 21732 22010 21788
rect 22010 21732 22014 21788
rect 21950 21728 22014 21732
rect 22030 21788 22094 21792
rect 22030 21732 22034 21788
rect 22034 21732 22090 21788
rect 22090 21732 22094 21788
rect 22030 21728 22094 21732
rect 28736 21788 28800 21792
rect 28736 21732 28740 21788
rect 28740 21732 28796 21788
rect 28796 21732 28800 21788
rect 28736 21728 28800 21732
rect 28816 21788 28880 21792
rect 28816 21732 28820 21788
rect 28820 21732 28876 21788
rect 28876 21732 28880 21788
rect 28816 21728 28880 21732
rect 28896 21788 28960 21792
rect 28896 21732 28900 21788
rect 28900 21732 28956 21788
rect 28956 21732 28960 21788
rect 28896 21728 28960 21732
rect 28976 21788 29040 21792
rect 28976 21732 28980 21788
rect 28980 21732 29036 21788
rect 29036 21732 29040 21788
rect 28976 21728 29040 21732
rect 4425 21244 4489 21248
rect 4425 21188 4429 21244
rect 4429 21188 4485 21244
rect 4485 21188 4489 21244
rect 4425 21184 4489 21188
rect 4505 21244 4569 21248
rect 4505 21188 4509 21244
rect 4509 21188 4565 21244
rect 4565 21188 4569 21244
rect 4505 21184 4569 21188
rect 4585 21244 4649 21248
rect 4585 21188 4589 21244
rect 4589 21188 4645 21244
rect 4645 21188 4649 21244
rect 4585 21184 4649 21188
rect 4665 21244 4729 21248
rect 4665 21188 4669 21244
rect 4669 21188 4725 21244
rect 4725 21188 4729 21244
rect 4665 21184 4729 21188
rect 11371 21244 11435 21248
rect 11371 21188 11375 21244
rect 11375 21188 11431 21244
rect 11431 21188 11435 21244
rect 11371 21184 11435 21188
rect 11451 21244 11515 21248
rect 11451 21188 11455 21244
rect 11455 21188 11511 21244
rect 11511 21188 11515 21244
rect 11451 21184 11515 21188
rect 11531 21244 11595 21248
rect 11531 21188 11535 21244
rect 11535 21188 11591 21244
rect 11591 21188 11595 21244
rect 11531 21184 11595 21188
rect 11611 21244 11675 21248
rect 11611 21188 11615 21244
rect 11615 21188 11671 21244
rect 11671 21188 11675 21244
rect 11611 21184 11675 21188
rect 18317 21244 18381 21248
rect 18317 21188 18321 21244
rect 18321 21188 18377 21244
rect 18377 21188 18381 21244
rect 18317 21184 18381 21188
rect 18397 21244 18461 21248
rect 18397 21188 18401 21244
rect 18401 21188 18457 21244
rect 18457 21188 18461 21244
rect 18397 21184 18461 21188
rect 18477 21244 18541 21248
rect 18477 21188 18481 21244
rect 18481 21188 18537 21244
rect 18537 21188 18541 21244
rect 18477 21184 18541 21188
rect 18557 21244 18621 21248
rect 18557 21188 18561 21244
rect 18561 21188 18617 21244
rect 18617 21188 18621 21244
rect 18557 21184 18621 21188
rect 25263 21244 25327 21248
rect 25263 21188 25267 21244
rect 25267 21188 25323 21244
rect 25323 21188 25327 21244
rect 25263 21184 25327 21188
rect 25343 21244 25407 21248
rect 25343 21188 25347 21244
rect 25347 21188 25403 21244
rect 25403 21188 25407 21244
rect 25343 21184 25407 21188
rect 25423 21244 25487 21248
rect 25423 21188 25427 21244
rect 25427 21188 25483 21244
rect 25483 21188 25487 21244
rect 25423 21184 25487 21188
rect 25503 21244 25567 21248
rect 25503 21188 25507 21244
rect 25507 21188 25563 21244
rect 25563 21188 25567 21244
rect 25503 21184 25567 21188
rect 7898 20700 7962 20704
rect 7898 20644 7902 20700
rect 7902 20644 7958 20700
rect 7958 20644 7962 20700
rect 7898 20640 7962 20644
rect 7978 20700 8042 20704
rect 7978 20644 7982 20700
rect 7982 20644 8038 20700
rect 8038 20644 8042 20700
rect 7978 20640 8042 20644
rect 8058 20700 8122 20704
rect 8058 20644 8062 20700
rect 8062 20644 8118 20700
rect 8118 20644 8122 20700
rect 8058 20640 8122 20644
rect 8138 20700 8202 20704
rect 8138 20644 8142 20700
rect 8142 20644 8198 20700
rect 8198 20644 8202 20700
rect 8138 20640 8202 20644
rect 14844 20700 14908 20704
rect 14844 20644 14848 20700
rect 14848 20644 14904 20700
rect 14904 20644 14908 20700
rect 14844 20640 14908 20644
rect 14924 20700 14988 20704
rect 14924 20644 14928 20700
rect 14928 20644 14984 20700
rect 14984 20644 14988 20700
rect 14924 20640 14988 20644
rect 15004 20700 15068 20704
rect 15004 20644 15008 20700
rect 15008 20644 15064 20700
rect 15064 20644 15068 20700
rect 15004 20640 15068 20644
rect 15084 20700 15148 20704
rect 15084 20644 15088 20700
rect 15088 20644 15144 20700
rect 15144 20644 15148 20700
rect 15084 20640 15148 20644
rect 21790 20700 21854 20704
rect 21790 20644 21794 20700
rect 21794 20644 21850 20700
rect 21850 20644 21854 20700
rect 21790 20640 21854 20644
rect 21870 20700 21934 20704
rect 21870 20644 21874 20700
rect 21874 20644 21930 20700
rect 21930 20644 21934 20700
rect 21870 20640 21934 20644
rect 21950 20700 22014 20704
rect 21950 20644 21954 20700
rect 21954 20644 22010 20700
rect 22010 20644 22014 20700
rect 21950 20640 22014 20644
rect 22030 20700 22094 20704
rect 22030 20644 22034 20700
rect 22034 20644 22090 20700
rect 22090 20644 22094 20700
rect 22030 20640 22094 20644
rect 28736 20700 28800 20704
rect 28736 20644 28740 20700
rect 28740 20644 28796 20700
rect 28796 20644 28800 20700
rect 28736 20640 28800 20644
rect 28816 20700 28880 20704
rect 28816 20644 28820 20700
rect 28820 20644 28876 20700
rect 28876 20644 28880 20700
rect 28816 20640 28880 20644
rect 28896 20700 28960 20704
rect 28896 20644 28900 20700
rect 28900 20644 28956 20700
rect 28956 20644 28960 20700
rect 28896 20640 28960 20644
rect 28976 20700 29040 20704
rect 28976 20644 28980 20700
rect 28980 20644 29036 20700
rect 29036 20644 29040 20700
rect 28976 20640 29040 20644
rect 4425 20156 4489 20160
rect 4425 20100 4429 20156
rect 4429 20100 4485 20156
rect 4485 20100 4489 20156
rect 4425 20096 4489 20100
rect 4505 20156 4569 20160
rect 4505 20100 4509 20156
rect 4509 20100 4565 20156
rect 4565 20100 4569 20156
rect 4505 20096 4569 20100
rect 4585 20156 4649 20160
rect 4585 20100 4589 20156
rect 4589 20100 4645 20156
rect 4645 20100 4649 20156
rect 4585 20096 4649 20100
rect 4665 20156 4729 20160
rect 4665 20100 4669 20156
rect 4669 20100 4725 20156
rect 4725 20100 4729 20156
rect 4665 20096 4729 20100
rect 11371 20156 11435 20160
rect 11371 20100 11375 20156
rect 11375 20100 11431 20156
rect 11431 20100 11435 20156
rect 11371 20096 11435 20100
rect 11451 20156 11515 20160
rect 11451 20100 11455 20156
rect 11455 20100 11511 20156
rect 11511 20100 11515 20156
rect 11451 20096 11515 20100
rect 11531 20156 11595 20160
rect 11531 20100 11535 20156
rect 11535 20100 11591 20156
rect 11591 20100 11595 20156
rect 11531 20096 11595 20100
rect 11611 20156 11675 20160
rect 11611 20100 11615 20156
rect 11615 20100 11671 20156
rect 11671 20100 11675 20156
rect 11611 20096 11675 20100
rect 18317 20156 18381 20160
rect 18317 20100 18321 20156
rect 18321 20100 18377 20156
rect 18377 20100 18381 20156
rect 18317 20096 18381 20100
rect 18397 20156 18461 20160
rect 18397 20100 18401 20156
rect 18401 20100 18457 20156
rect 18457 20100 18461 20156
rect 18397 20096 18461 20100
rect 18477 20156 18541 20160
rect 18477 20100 18481 20156
rect 18481 20100 18537 20156
rect 18537 20100 18541 20156
rect 18477 20096 18541 20100
rect 18557 20156 18621 20160
rect 18557 20100 18561 20156
rect 18561 20100 18617 20156
rect 18617 20100 18621 20156
rect 18557 20096 18621 20100
rect 25263 20156 25327 20160
rect 25263 20100 25267 20156
rect 25267 20100 25323 20156
rect 25323 20100 25327 20156
rect 25263 20096 25327 20100
rect 25343 20156 25407 20160
rect 25343 20100 25347 20156
rect 25347 20100 25403 20156
rect 25403 20100 25407 20156
rect 25343 20096 25407 20100
rect 25423 20156 25487 20160
rect 25423 20100 25427 20156
rect 25427 20100 25483 20156
rect 25483 20100 25487 20156
rect 25423 20096 25487 20100
rect 25503 20156 25567 20160
rect 25503 20100 25507 20156
rect 25507 20100 25563 20156
rect 25563 20100 25567 20156
rect 25503 20096 25567 20100
rect 7898 19612 7962 19616
rect 7898 19556 7902 19612
rect 7902 19556 7958 19612
rect 7958 19556 7962 19612
rect 7898 19552 7962 19556
rect 7978 19612 8042 19616
rect 7978 19556 7982 19612
rect 7982 19556 8038 19612
rect 8038 19556 8042 19612
rect 7978 19552 8042 19556
rect 8058 19612 8122 19616
rect 8058 19556 8062 19612
rect 8062 19556 8118 19612
rect 8118 19556 8122 19612
rect 8058 19552 8122 19556
rect 8138 19612 8202 19616
rect 8138 19556 8142 19612
rect 8142 19556 8198 19612
rect 8198 19556 8202 19612
rect 8138 19552 8202 19556
rect 14844 19612 14908 19616
rect 14844 19556 14848 19612
rect 14848 19556 14904 19612
rect 14904 19556 14908 19612
rect 14844 19552 14908 19556
rect 14924 19612 14988 19616
rect 14924 19556 14928 19612
rect 14928 19556 14984 19612
rect 14984 19556 14988 19612
rect 14924 19552 14988 19556
rect 15004 19612 15068 19616
rect 15004 19556 15008 19612
rect 15008 19556 15064 19612
rect 15064 19556 15068 19612
rect 15004 19552 15068 19556
rect 15084 19612 15148 19616
rect 15084 19556 15088 19612
rect 15088 19556 15144 19612
rect 15144 19556 15148 19612
rect 15084 19552 15148 19556
rect 21790 19612 21854 19616
rect 21790 19556 21794 19612
rect 21794 19556 21850 19612
rect 21850 19556 21854 19612
rect 21790 19552 21854 19556
rect 21870 19612 21934 19616
rect 21870 19556 21874 19612
rect 21874 19556 21930 19612
rect 21930 19556 21934 19612
rect 21870 19552 21934 19556
rect 21950 19612 22014 19616
rect 21950 19556 21954 19612
rect 21954 19556 22010 19612
rect 22010 19556 22014 19612
rect 21950 19552 22014 19556
rect 22030 19612 22094 19616
rect 22030 19556 22034 19612
rect 22034 19556 22090 19612
rect 22090 19556 22094 19612
rect 22030 19552 22094 19556
rect 28736 19612 28800 19616
rect 28736 19556 28740 19612
rect 28740 19556 28796 19612
rect 28796 19556 28800 19612
rect 28736 19552 28800 19556
rect 28816 19612 28880 19616
rect 28816 19556 28820 19612
rect 28820 19556 28876 19612
rect 28876 19556 28880 19612
rect 28816 19552 28880 19556
rect 28896 19612 28960 19616
rect 28896 19556 28900 19612
rect 28900 19556 28956 19612
rect 28956 19556 28960 19612
rect 28896 19552 28960 19556
rect 28976 19612 29040 19616
rect 28976 19556 28980 19612
rect 28980 19556 29036 19612
rect 29036 19556 29040 19612
rect 28976 19552 29040 19556
rect 4425 19068 4489 19072
rect 4425 19012 4429 19068
rect 4429 19012 4485 19068
rect 4485 19012 4489 19068
rect 4425 19008 4489 19012
rect 4505 19068 4569 19072
rect 4505 19012 4509 19068
rect 4509 19012 4565 19068
rect 4565 19012 4569 19068
rect 4505 19008 4569 19012
rect 4585 19068 4649 19072
rect 4585 19012 4589 19068
rect 4589 19012 4645 19068
rect 4645 19012 4649 19068
rect 4585 19008 4649 19012
rect 4665 19068 4729 19072
rect 4665 19012 4669 19068
rect 4669 19012 4725 19068
rect 4725 19012 4729 19068
rect 4665 19008 4729 19012
rect 11371 19068 11435 19072
rect 11371 19012 11375 19068
rect 11375 19012 11431 19068
rect 11431 19012 11435 19068
rect 11371 19008 11435 19012
rect 11451 19068 11515 19072
rect 11451 19012 11455 19068
rect 11455 19012 11511 19068
rect 11511 19012 11515 19068
rect 11451 19008 11515 19012
rect 11531 19068 11595 19072
rect 11531 19012 11535 19068
rect 11535 19012 11591 19068
rect 11591 19012 11595 19068
rect 11531 19008 11595 19012
rect 11611 19068 11675 19072
rect 11611 19012 11615 19068
rect 11615 19012 11671 19068
rect 11671 19012 11675 19068
rect 11611 19008 11675 19012
rect 18317 19068 18381 19072
rect 18317 19012 18321 19068
rect 18321 19012 18377 19068
rect 18377 19012 18381 19068
rect 18317 19008 18381 19012
rect 18397 19068 18461 19072
rect 18397 19012 18401 19068
rect 18401 19012 18457 19068
rect 18457 19012 18461 19068
rect 18397 19008 18461 19012
rect 18477 19068 18541 19072
rect 18477 19012 18481 19068
rect 18481 19012 18537 19068
rect 18537 19012 18541 19068
rect 18477 19008 18541 19012
rect 18557 19068 18621 19072
rect 18557 19012 18561 19068
rect 18561 19012 18617 19068
rect 18617 19012 18621 19068
rect 18557 19008 18621 19012
rect 25263 19068 25327 19072
rect 25263 19012 25267 19068
rect 25267 19012 25323 19068
rect 25323 19012 25327 19068
rect 25263 19008 25327 19012
rect 25343 19068 25407 19072
rect 25343 19012 25347 19068
rect 25347 19012 25403 19068
rect 25403 19012 25407 19068
rect 25343 19008 25407 19012
rect 25423 19068 25487 19072
rect 25423 19012 25427 19068
rect 25427 19012 25483 19068
rect 25483 19012 25487 19068
rect 25423 19008 25487 19012
rect 25503 19068 25567 19072
rect 25503 19012 25507 19068
rect 25507 19012 25563 19068
rect 25563 19012 25567 19068
rect 25503 19008 25567 19012
rect 7898 18524 7962 18528
rect 7898 18468 7902 18524
rect 7902 18468 7958 18524
rect 7958 18468 7962 18524
rect 7898 18464 7962 18468
rect 7978 18524 8042 18528
rect 7978 18468 7982 18524
rect 7982 18468 8038 18524
rect 8038 18468 8042 18524
rect 7978 18464 8042 18468
rect 8058 18524 8122 18528
rect 8058 18468 8062 18524
rect 8062 18468 8118 18524
rect 8118 18468 8122 18524
rect 8058 18464 8122 18468
rect 8138 18524 8202 18528
rect 8138 18468 8142 18524
rect 8142 18468 8198 18524
rect 8198 18468 8202 18524
rect 8138 18464 8202 18468
rect 14844 18524 14908 18528
rect 14844 18468 14848 18524
rect 14848 18468 14904 18524
rect 14904 18468 14908 18524
rect 14844 18464 14908 18468
rect 14924 18524 14988 18528
rect 14924 18468 14928 18524
rect 14928 18468 14984 18524
rect 14984 18468 14988 18524
rect 14924 18464 14988 18468
rect 15004 18524 15068 18528
rect 15004 18468 15008 18524
rect 15008 18468 15064 18524
rect 15064 18468 15068 18524
rect 15004 18464 15068 18468
rect 15084 18524 15148 18528
rect 15084 18468 15088 18524
rect 15088 18468 15144 18524
rect 15144 18468 15148 18524
rect 15084 18464 15148 18468
rect 21790 18524 21854 18528
rect 21790 18468 21794 18524
rect 21794 18468 21850 18524
rect 21850 18468 21854 18524
rect 21790 18464 21854 18468
rect 21870 18524 21934 18528
rect 21870 18468 21874 18524
rect 21874 18468 21930 18524
rect 21930 18468 21934 18524
rect 21870 18464 21934 18468
rect 21950 18524 22014 18528
rect 21950 18468 21954 18524
rect 21954 18468 22010 18524
rect 22010 18468 22014 18524
rect 21950 18464 22014 18468
rect 22030 18524 22094 18528
rect 22030 18468 22034 18524
rect 22034 18468 22090 18524
rect 22090 18468 22094 18524
rect 22030 18464 22094 18468
rect 28736 18524 28800 18528
rect 28736 18468 28740 18524
rect 28740 18468 28796 18524
rect 28796 18468 28800 18524
rect 28736 18464 28800 18468
rect 28816 18524 28880 18528
rect 28816 18468 28820 18524
rect 28820 18468 28876 18524
rect 28876 18468 28880 18524
rect 28816 18464 28880 18468
rect 28896 18524 28960 18528
rect 28896 18468 28900 18524
rect 28900 18468 28956 18524
rect 28956 18468 28960 18524
rect 28896 18464 28960 18468
rect 28976 18524 29040 18528
rect 28976 18468 28980 18524
rect 28980 18468 29036 18524
rect 29036 18468 29040 18524
rect 28976 18464 29040 18468
rect 4425 17980 4489 17984
rect 4425 17924 4429 17980
rect 4429 17924 4485 17980
rect 4485 17924 4489 17980
rect 4425 17920 4489 17924
rect 4505 17980 4569 17984
rect 4505 17924 4509 17980
rect 4509 17924 4565 17980
rect 4565 17924 4569 17980
rect 4505 17920 4569 17924
rect 4585 17980 4649 17984
rect 4585 17924 4589 17980
rect 4589 17924 4645 17980
rect 4645 17924 4649 17980
rect 4585 17920 4649 17924
rect 4665 17980 4729 17984
rect 4665 17924 4669 17980
rect 4669 17924 4725 17980
rect 4725 17924 4729 17980
rect 4665 17920 4729 17924
rect 11371 17980 11435 17984
rect 11371 17924 11375 17980
rect 11375 17924 11431 17980
rect 11431 17924 11435 17980
rect 11371 17920 11435 17924
rect 11451 17980 11515 17984
rect 11451 17924 11455 17980
rect 11455 17924 11511 17980
rect 11511 17924 11515 17980
rect 11451 17920 11515 17924
rect 11531 17980 11595 17984
rect 11531 17924 11535 17980
rect 11535 17924 11591 17980
rect 11591 17924 11595 17980
rect 11531 17920 11595 17924
rect 11611 17980 11675 17984
rect 11611 17924 11615 17980
rect 11615 17924 11671 17980
rect 11671 17924 11675 17980
rect 11611 17920 11675 17924
rect 18317 17980 18381 17984
rect 18317 17924 18321 17980
rect 18321 17924 18377 17980
rect 18377 17924 18381 17980
rect 18317 17920 18381 17924
rect 18397 17980 18461 17984
rect 18397 17924 18401 17980
rect 18401 17924 18457 17980
rect 18457 17924 18461 17980
rect 18397 17920 18461 17924
rect 18477 17980 18541 17984
rect 18477 17924 18481 17980
rect 18481 17924 18537 17980
rect 18537 17924 18541 17980
rect 18477 17920 18541 17924
rect 18557 17980 18621 17984
rect 18557 17924 18561 17980
rect 18561 17924 18617 17980
rect 18617 17924 18621 17980
rect 18557 17920 18621 17924
rect 25263 17980 25327 17984
rect 25263 17924 25267 17980
rect 25267 17924 25323 17980
rect 25323 17924 25327 17980
rect 25263 17920 25327 17924
rect 25343 17980 25407 17984
rect 25343 17924 25347 17980
rect 25347 17924 25403 17980
rect 25403 17924 25407 17980
rect 25343 17920 25407 17924
rect 25423 17980 25487 17984
rect 25423 17924 25427 17980
rect 25427 17924 25483 17980
rect 25483 17924 25487 17980
rect 25423 17920 25487 17924
rect 25503 17980 25567 17984
rect 25503 17924 25507 17980
rect 25507 17924 25563 17980
rect 25563 17924 25567 17980
rect 25503 17920 25567 17924
rect 7898 17436 7962 17440
rect 7898 17380 7902 17436
rect 7902 17380 7958 17436
rect 7958 17380 7962 17436
rect 7898 17376 7962 17380
rect 7978 17436 8042 17440
rect 7978 17380 7982 17436
rect 7982 17380 8038 17436
rect 8038 17380 8042 17436
rect 7978 17376 8042 17380
rect 8058 17436 8122 17440
rect 8058 17380 8062 17436
rect 8062 17380 8118 17436
rect 8118 17380 8122 17436
rect 8058 17376 8122 17380
rect 8138 17436 8202 17440
rect 8138 17380 8142 17436
rect 8142 17380 8198 17436
rect 8198 17380 8202 17436
rect 8138 17376 8202 17380
rect 14844 17436 14908 17440
rect 14844 17380 14848 17436
rect 14848 17380 14904 17436
rect 14904 17380 14908 17436
rect 14844 17376 14908 17380
rect 14924 17436 14988 17440
rect 14924 17380 14928 17436
rect 14928 17380 14984 17436
rect 14984 17380 14988 17436
rect 14924 17376 14988 17380
rect 15004 17436 15068 17440
rect 15004 17380 15008 17436
rect 15008 17380 15064 17436
rect 15064 17380 15068 17436
rect 15004 17376 15068 17380
rect 15084 17436 15148 17440
rect 15084 17380 15088 17436
rect 15088 17380 15144 17436
rect 15144 17380 15148 17436
rect 15084 17376 15148 17380
rect 21790 17436 21854 17440
rect 21790 17380 21794 17436
rect 21794 17380 21850 17436
rect 21850 17380 21854 17436
rect 21790 17376 21854 17380
rect 21870 17436 21934 17440
rect 21870 17380 21874 17436
rect 21874 17380 21930 17436
rect 21930 17380 21934 17436
rect 21870 17376 21934 17380
rect 21950 17436 22014 17440
rect 21950 17380 21954 17436
rect 21954 17380 22010 17436
rect 22010 17380 22014 17436
rect 21950 17376 22014 17380
rect 22030 17436 22094 17440
rect 22030 17380 22034 17436
rect 22034 17380 22090 17436
rect 22090 17380 22094 17436
rect 22030 17376 22094 17380
rect 28736 17436 28800 17440
rect 28736 17380 28740 17436
rect 28740 17380 28796 17436
rect 28796 17380 28800 17436
rect 28736 17376 28800 17380
rect 28816 17436 28880 17440
rect 28816 17380 28820 17436
rect 28820 17380 28876 17436
rect 28876 17380 28880 17436
rect 28816 17376 28880 17380
rect 28896 17436 28960 17440
rect 28896 17380 28900 17436
rect 28900 17380 28956 17436
rect 28956 17380 28960 17436
rect 28896 17376 28960 17380
rect 28976 17436 29040 17440
rect 28976 17380 28980 17436
rect 28980 17380 29036 17436
rect 29036 17380 29040 17436
rect 28976 17376 29040 17380
rect 4425 16892 4489 16896
rect 4425 16836 4429 16892
rect 4429 16836 4485 16892
rect 4485 16836 4489 16892
rect 4425 16832 4489 16836
rect 4505 16892 4569 16896
rect 4505 16836 4509 16892
rect 4509 16836 4565 16892
rect 4565 16836 4569 16892
rect 4505 16832 4569 16836
rect 4585 16892 4649 16896
rect 4585 16836 4589 16892
rect 4589 16836 4645 16892
rect 4645 16836 4649 16892
rect 4585 16832 4649 16836
rect 4665 16892 4729 16896
rect 4665 16836 4669 16892
rect 4669 16836 4725 16892
rect 4725 16836 4729 16892
rect 4665 16832 4729 16836
rect 11371 16892 11435 16896
rect 11371 16836 11375 16892
rect 11375 16836 11431 16892
rect 11431 16836 11435 16892
rect 11371 16832 11435 16836
rect 11451 16892 11515 16896
rect 11451 16836 11455 16892
rect 11455 16836 11511 16892
rect 11511 16836 11515 16892
rect 11451 16832 11515 16836
rect 11531 16892 11595 16896
rect 11531 16836 11535 16892
rect 11535 16836 11591 16892
rect 11591 16836 11595 16892
rect 11531 16832 11595 16836
rect 11611 16892 11675 16896
rect 11611 16836 11615 16892
rect 11615 16836 11671 16892
rect 11671 16836 11675 16892
rect 11611 16832 11675 16836
rect 18317 16892 18381 16896
rect 18317 16836 18321 16892
rect 18321 16836 18377 16892
rect 18377 16836 18381 16892
rect 18317 16832 18381 16836
rect 18397 16892 18461 16896
rect 18397 16836 18401 16892
rect 18401 16836 18457 16892
rect 18457 16836 18461 16892
rect 18397 16832 18461 16836
rect 18477 16892 18541 16896
rect 18477 16836 18481 16892
rect 18481 16836 18537 16892
rect 18537 16836 18541 16892
rect 18477 16832 18541 16836
rect 18557 16892 18621 16896
rect 18557 16836 18561 16892
rect 18561 16836 18617 16892
rect 18617 16836 18621 16892
rect 18557 16832 18621 16836
rect 25263 16892 25327 16896
rect 25263 16836 25267 16892
rect 25267 16836 25323 16892
rect 25323 16836 25327 16892
rect 25263 16832 25327 16836
rect 25343 16892 25407 16896
rect 25343 16836 25347 16892
rect 25347 16836 25403 16892
rect 25403 16836 25407 16892
rect 25343 16832 25407 16836
rect 25423 16892 25487 16896
rect 25423 16836 25427 16892
rect 25427 16836 25483 16892
rect 25483 16836 25487 16892
rect 25423 16832 25487 16836
rect 25503 16892 25567 16896
rect 25503 16836 25507 16892
rect 25507 16836 25563 16892
rect 25563 16836 25567 16892
rect 25503 16832 25567 16836
rect 7898 16348 7962 16352
rect 7898 16292 7902 16348
rect 7902 16292 7958 16348
rect 7958 16292 7962 16348
rect 7898 16288 7962 16292
rect 7978 16348 8042 16352
rect 7978 16292 7982 16348
rect 7982 16292 8038 16348
rect 8038 16292 8042 16348
rect 7978 16288 8042 16292
rect 8058 16348 8122 16352
rect 8058 16292 8062 16348
rect 8062 16292 8118 16348
rect 8118 16292 8122 16348
rect 8058 16288 8122 16292
rect 8138 16348 8202 16352
rect 8138 16292 8142 16348
rect 8142 16292 8198 16348
rect 8198 16292 8202 16348
rect 8138 16288 8202 16292
rect 14844 16348 14908 16352
rect 14844 16292 14848 16348
rect 14848 16292 14904 16348
rect 14904 16292 14908 16348
rect 14844 16288 14908 16292
rect 14924 16348 14988 16352
rect 14924 16292 14928 16348
rect 14928 16292 14984 16348
rect 14984 16292 14988 16348
rect 14924 16288 14988 16292
rect 15004 16348 15068 16352
rect 15004 16292 15008 16348
rect 15008 16292 15064 16348
rect 15064 16292 15068 16348
rect 15004 16288 15068 16292
rect 15084 16348 15148 16352
rect 15084 16292 15088 16348
rect 15088 16292 15144 16348
rect 15144 16292 15148 16348
rect 15084 16288 15148 16292
rect 21790 16348 21854 16352
rect 21790 16292 21794 16348
rect 21794 16292 21850 16348
rect 21850 16292 21854 16348
rect 21790 16288 21854 16292
rect 21870 16348 21934 16352
rect 21870 16292 21874 16348
rect 21874 16292 21930 16348
rect 21930 16292 21934 16348
rect 21870 16288 21934 16292
rect 21950 16348 22014 16352
rect 21950 16292 21954 16348
rect 21954 16292 22010 16348
rect 22010 16292 22014 16348
rect 21950 16288 22014 16292
rect 22030 16348 22094 16352
rect 22030 16292 22034 16348
rect 22034 16292 22090 16348
rect 22090 16292 22094 16348
rect 22030 16288 22094 16292
rect 28736 16348 28800 16352
rect 28736 16292 28740 16348
rect 28740 16292 28796 16348
rect 28796 16292 28800 16348
rect 28736 16288 28800 16292
rect 28816 16348 28880 16352
rect 28816 16292 28820 16348
rect 28820 16292 28876 16348
rect 28876 16292 28880 16348
rect 28816 16288 28880 16292
rect 28896 16348 28960 16352
rect 28896 16292 28900 16348
rect 28900 16292 28956 16348
rect 28956 16292 28960 16348
rect 28896 16288 28960 16292
rect 28976 16348 29040 16352
rect 28976 16292 28980 16348
rect 28980 16292 29036 16348
rect 29036 16292 29040 16348
rect 28976 16288 29040 16292
rect 4425 15804 4489 15808
rect 4425 15748 4429 15804
rect 4429 15748 4485 15804
rect 4485 15748 4489 15804
rect 4425 15744 4489 15748
rect 4505 15804 4569 15808
rect 4505 15748 4509 15804
rect 4509 15748 4565 15804
rect 4565 15748 4569 15804
rect 4505 15744 4569 15748
rect 4585 15804 4649 15808
rect 4585 15748 4589 15804
rect 4589 15748 4645 15804
rect 4645 15748 4649 15804
rect 4585 15744 4649 15748
rect 4665 15804 4729 15808
rect 4665 15748 4669 15804
rect 4669 15748 4725 15804
rect 4725 15748 4729 15804
rect 4665 15744 4729 15748
rect 11371 15804 11435 15808
rect 11371 15748 11375 15804
rect 11375 15748 11431 15804
rect 11431 15748 11435 15804
rect 11371 15744 11435 15748
rect 11451 15804 11515 15808
rect 11451 15748 11455 15804
rect 11455 15748 11511 15804
rect 11511 15748 11515 15804
rect 11451 15744 11515 15748
rect 11531 15804 11595 15808
rect 11531 15748 11535 15804
rect 11535 15748 11591 15804
rect 11591 15748 11595 15804
rect 11531 15744 11595 15748
rect 11611 15804 11675 15808
rect 11611 15748 11615 15804
rect 11615 15748 11671 15804
rect 11671 15748 11675 15804
rect 11611 15744 11675 15748
rect 18317 15804 18381 15808
rect 18317 15748 18321 15804
rect 18321 15748 18377 15804
rect 18377 15748 18381 15804
rect 18317 15744 18381 15748
rect 18397 15804 18461 15808
rect 18397 15748 18401 15804
rect 18401 15748 18457 15804
rect 18457 15748 18461 15804
rect 18397 15744 18461 15748
rect 18477 15804 18541 15808
rect 18477 15748 18481 15804
rect 18481 15748 18537 15804
rect 18537 15748 18541 15804
rect 18477 15744 18541 15748
rect 18557 15804 18621 15808
rect 18557 15748 18561 15804
rect 18561 15748 18617 15804
rect 18617 15748 18621 15804
rect 18557 15744 18621 15748
rect 25263 15804 25327 15808
rect 25263 15748 25267 15804
rect 25267 15748 25323 15804
rect 25323 15748 25327 15804
rect 25263 15744 25327 15748
rect 25343 15804 25407 15808
rect 25343 15748 25347 15804
rect 25347 15748 25403 15804
rect 25403 15748 25407 15804
rect 25343 15744 25407 15748
rect 25423 15804 25487 15808
rect 25423 15748 25427 15804
rect 25427 15748 25483 15804
rect 25483 15748 25487 15804
rect 25423 15744 25487 15748
rect 25503 15804 25567 15808
rect 25503 15748 25507 15804
rect 25507 15748 25563 15804
rect 25563 15748 25567 15804
rect 25503 15744 25567 15748
rect 7898 15260 7962 15264
rect 7898 15204 7902 15260
rect 7902 15204 7958 15260
rect 7958 15204 7962 15260
rect 7898 15200 7962 15204
rect 7978 15260 8042 15264
rect 7978 15204 7982 15260
rect 7982 15204 8038 15260
rect 8038 15204 8042 15260
rect 7978 15200 8042 15204
rect 8058 15260 8122 15264
rect 8058 15204 8062 15260
rect 8062 15204 8118 15260
rect 8118 15204 8122 15260
rect 8058 15200 8122 15204
rect 8138 15260 8202 15264
rect 8138 15204 8142 15260
rect 8142 15204 8198 15260
rect 8198 15204 8202 15260
rect 8138 15200 8202 15204
rect 14844 15260 14908 15264
rect 14844 15204 14848 15260
rect 14848 15204 14904 15260
rect 14904 15204 14908 15260
rect 14844 15200 14908 15204
rect 14924 15260 14988 15264
rect 14924 15204 14928 15260
rect 14928 15204 14984 15260
rect 14984 15204 14988 15260
rect 14924 15200 14988 15204
rect 15004 15260 15068 15264
rect 15004 15204 15008 15260
rect 15008 15204 15064 15260
rect 15064 15204 15068 15260
rect 15004 15200 15068 15204
rect 15084 15260 15148 15264
rect 15084 15204 15088 15260
rect 15088 15204 15144 15260
rect 15144 15204 15148 15260
rect 15084 15200 15148 15204
rect 21790 15260 21854 15264
rect 21790 15204 21794 15260
rect 21794 15204 21850 15260
rect 21850 15204 21854 15260
rect 21790 15200 21854 15204
rect 21870 15260 21934 15264
rect 21870 15204 21874 15260
rect 21874 15204 21930 15260
rect 21930 15204 21934 15260
rect 21870 15200 21934 15204
rect 21950 15260 22014 15264
rect 21950 15204 21954 15260
rect 21954 15204 22010 15260
rect 22010 15204 22014 15260
rect 21950 15200 22014 15204
rect 22030 15260 22094 15264
rect 22030 15204 22034 15260
rect 22034 15204 22090 15260
rect 22090 15204 22094 15260
rect 22030 15200 22094 15204
rect 28736 15260 28800 15264
rect 28736 15204 28740 15260
rect 28740 15204 28796 15260
rect 28796 15204 28800 15260
rect 28736 15200 28800 15204
rect 28816 15260 28880 15264
rect 28816 15204 28820 15260
rect 28820 15204 28876 15260
rect 28876 15204 28880 15260
rect 28816 15200 28880 15204
rect 28896 15260 28960 15264
rect 28896 15204 28900 15260
rect 28900 15204 28956 15260
rect 28956 15204 28960 15260
rect 28896 15200 28960 15204
rect 28976 15260 29040 15264
rect 28976 15204 28980 15260
rect 28980 15204 29036 15260
rect 29036 15204 29040 15260
rect 28976 15200 29040 15204
rect 4425 14716 4489 14720
rect 4425 14660 4429 14716
rect 4429 14660 4485 14716
rect 4485 14660 4489 14716
rect 4425 14656 4489 14660
rect 4505 14716 4569 14720
rect 4505 14660 4509 14716
rect 4509 14660 4565 14716
rect 4565 14660 4569 14716
rect 4505 14656 4569 14660
rect 4585 14716 4649 14720
rect 4585 14660 4589 14716
rect 4589 14660 4645 14716
rect 4645 14660 4649 14716
rect 4585 14656 4649 14660
rect 4665 14716 4729 14720
rect 4665 14660 4669 14716
rect 4669 14660 4725 14716
rect 4725 14660 4729 14716
rect 4665 14656 4729 14660
rect 11371 14716 11435 14720
rect 11371 14660 11375 14716
rect 11375 14660 11431 14716
rect 11431 14660 11435 14716
rect 11371 14656 11435 14660
rect 11451 14716 11515 14720
rect 11451 14660 11455 14716
rect 11455 14660 11511 14716
rect 11511 14660 11515 14716
rect 11451 14656 11515 14660
rect 11531 14716 11595 14720
rect 11531 14660 11535 14716
rect 11535 14660 11591 14716
rect 11591 14660 11595 14716
rect 11531 14656 11595 14660
rect 11611 14716 11675 14720
rect 11611 14660 11615 14716
rect 11615 14660 11671 14716
rect 11671 14660 11675 14716
rect 11611 14656 11675 14660
rect 18317 14716 18381 14720
rect 18317 14660 18321 14716
rect 18321 14660 18377 14716
rect 18377 14660 18381 14716
rect 18317 14656 18381 14660
rect 18397 14716 18461 14720
rect 18397 14660 18401 14716
rect 18401 14660 18457 14716
rect 18457 14660 18461 14716
rect 18397 14656 18461 14660
rect 18477 14716 18541 14720
rect 18477 14660 18481 14716
rect 18481 14660 18537 14716
rect 18537 14660 18541 14716
rect 18477 14656 18541 14660
rect 18557 14716 18621 14720
rect 18557 14660 18561 14716
rect 18561 14660 18617 14716
rect 18617 14660 18621 14716
rect 18557 14656 18621 14660
rect 25263 14716 25327 14720
rect 25263 14660 25267 14716
rect 25267 14660 25323 14716
rect 25323 14660 25327 14716
rect 25263 14656 25327 14660
rect 25343 14716 25407 14720
rect 25343 14660 25347 14716
rect 25347 14660 25403 14716
rect 25403 14660 25407 14716
rect 25343 14656 25407 14660
rect 25423 14716 25487 14720
rect 25423 14660 25427 14716
rect 25427 14660 25483 14716
rect 25483 14660 25487 14716
rect 25423 14656 25487 14660
rect 25503 14716 25567 14720
rect 25503 14660 25507 14716
rect 25507 14660 25563 14716
rect 25563 14660 25567 14716
rect 25503 14656 25567 14660
rect 7898 14172 7962 14176
rect 7898 14116 7902 14172
rect 7902 14116 7958 14172
rect 7958 14116 7962 14172
rect 7898 14112 7962 14116
rect 7978 14172 8042 14176
rect 7978 14116 7982 14172
rect 7982 14116 8038 14172
rect 8038 14116 8042 14172
rect 7978 14112 8042 14116
rect 8058 14172 8122 14176
rect 8058 14116 8062 14172
rect 8062 14116 8118 14172
rect 8118 14116 8122 14172
rect 8058 14112 8122 14116
rect 8138 14172 8202 14176
rect 8138 14116 8142 14172
rect 8142 14116 8198 14172
rect 8198 14116 8202 14172
rect 8138 14112 8202 14116
rect 14844 14172 14908 14176
rect 14844 14116 14848 14172
rect 14848 14116 14904 14172
rect 14904 14116 14908 14172
rect 14844 14112 14908 14116
rect 14924 14172 14988 14176
rect 14924 14116 14928 14172
rect 14928 14116 14984 14172
rect 14984 14116 14988 14172
rect 14924 14112 14988 14116
rect 15004 14172 15068 14176
rect 15004 14116 15008 14172
rect 15008 14116 15064 14172
rect 15064 14116 15068 14172
rect 15004 14112 15068 14116
rect 15084 14172 15148 14176
rect 15084 14116 15088 14172
rect 15088 14116 15144 14172
rect 15144 14116 15148 14172
rect 15084 14112 15148 14116
rect 21790 14172 21854 14176
rect 21790 14116 21794 14172
rect 21794 14116 21850 14172
rect 21850 14116 21854 14172
rect 21790 14112 21854 14116
rect 21870 14172 21934 14176
rect 21870 14116 21874 14172
rect 21874 14116 21930 14172
rect 21930 14116 21934 14172
rect 21870 14112 21934 14116
rect 21950 14172 22014 14176
rect 21950 14116 21954 14172
rect 21954 14116 22010 14172
rect 22010 14116 22014 14172
rect 21950 14112 22014 14116
rect 22030 14172 22094 14176
rect 22030 14116 22034 14172
rect 22034 14116 22090 14172
rect 22090 14116 22094 14172
rect 22030 14112 22094 14116
rect 28736 14172 28800 14176
rect 28736 14116 28740 14172
rect 28740 14116 28796 14172
rect 28796 14116 28800 14172
rect 28736 14112 28800 14116
rect 28816 14172 28880 14176
rect 28816 14116 28820 14172
rect 28820 14116 28876 14172
rect 28876 14116 28880 14172
rect 28816 14112 28880 14116
rect 28896 14172 28960 14176
rect 28896 14116 28900 14172
rect 28900 14116 28956 14172
rect 28956 14116 28960 14172
rect 28896 14112 28960 14116
rect 28976 14172 29040 14176
rect 28976 14116 28980 14172
rect 28980 14116 29036 14172
rect 29036 14116 29040 14172
rect 28976 14112 29040 14116
rect 4425 13628 4489 13632
rect 4425 13572 4429 13628
rect 4429 13572 4485 13628
rect 4485 13572 4489 13628
rect 4425 13568 4489 13572
rect 4505 13628 4569 13632
rect 4505 13572 4509 13628
rect 4509 13572 4565 13628
rect 4565 13572 4569 13628
rect 4505 13568 4569 13572
rect 4585 13628 4649 13632
rect 4585 13572 4589 13628
rect 4589 13572 4645 13628
rect 4645 13572 4649 13628
rect 4585 13568 4649 13572
rect 4665 13628 4729 13632
rect 4665 13572 4669 13628
rect 4669 13572 4725 13628
rect 4725 13572 4729 13628
rect 4665 13568 4729 13572
rect 11371 13628 11435 13632
rect 11371 13572 11375 13628
rect 11375 13572 11431 13628
rect 11431 13572 11435 13628
rect 11371 13568 11435 13572
rect 11451 13628 11515 13632
rect 11451 13572 11455 13628
rect 11455 13572 11511 13628
rect 11511 13572 11515 13628
rect 11451 13568 11515 13572
rect 11531 13628 11595 13632
rect 11531 13572 11535 13628
rect 11535 13572 11591 13628
rect 11591 13572 11595 13628
rect 11531 13568 11595 13572
rect 11611 13628 11675 13632
rect 11611 13572 11615 13628
rect 11615 13572 11671 13628
rect 11671 13572 11675 13628
rect 11611 13568 11675 13572
rect 18317 13628 18381 13632
rect 18317 13572 18321 13628
rect 18321 13572 18377 13628
rect 18377 13572 18381 13628
rect 18317 13568 18381 13572
rect 18397 13628 18461 13632
rect 18397 13572 18401 13628
rect 18401 13572 18457 13628
rect 18457 13572 18461 13628
rect 18397 13568 18461 13572
rect 18477 13628 18541 13632
rect 18477 13572 18481 13628
rect 18481 13572 18537 13628
rect 18537 13572 18541 13628
rect 18477 13568 18541 13572
rect 18557 13628 18621 13632
rect 18557 13572 18561 13628
rect 18561 13572 18617 13628
rect 18617 13572 18621 13628
rect 18557 13568 18621 13572
rect 25263 13628 25327 13632
rect 25263 13572 25267 13628
rect 25267 13572 25323 13628
rect 25323 13572 25327 13628
rect 25263 13568 25327 13572
rect 25343 13628 25407 13632
rect 25343 13572 25347 13628
rect 25347 13572 25403 13628
rect 25403 13572 25407 13628
rect 25343 13568 25407 13572
rect 25423 13628 25487 13632
rect 25423 13572 25427 13628
rect 25427 13572 25483 13628
rect 25483 13572 25487 13628
rect 25423 13568 25487 13572
rect 25503 13628 25567 13632
rect 25503 13572 25507 13628
rect 25507 13572 25563 13628
rect 25563 13572 25567 13628
rect 25503 13568 25567 13572
rect 7898 13084 7962 13088
rect 7898 13028 7902 13084
rect 7902 13028 7958 13084
rect 7958 13028 7962 13084
rect 7898 13024 7962 13028
rect 7978 13084 8042 13088
rect 7978 13028 7982 13084
rect 7982 13028 8038 13084
rect 8038 13028 8042 13084
rect 7978 13024 8042 13028
rect 8058 13084 8122 13088
rect 8058 13028 8062 13084
rect 8062 13028 8118 13084
rect 8118 13028 8122 13084
rect 8058 13024 8122 13028
rect 8138 13084 8202 13088
rect 8138 13028 8142 13084
rect 8142 13028 8198 13084
rect 8198 13028 8202 13084
rect 8138 13024 8202 13028
rect 14844 13084 14908 13088
rect 14844 13028 14848 13084
rect 14848 13028 14904 13084
rect 14904 13028 14908 13084
rect 14844 13024 14908 13028
rect 14924 13084 14988 13088
rect 14924 13028 14928 13084
rect 14928 13028 14984 13084
rect 14984 13028 14988 13084
rect 14924 13024 14988 13028
rect 15004 13084 15068 13088
rect 15004 13028 15008 13084
rect 15008 13028 15064 13084
rect 15064 13028 15068 13084
rect 15004 13024 15068 13028
rect 15084 13084 15148 13088
rect 15084 13028 15088 13084
rect 15088 13028 15144 13084
rect 15144 13028 15148 13084
rect 15084 13024 15148 13028
rect 21790 13084 21854 13088
rect 21790 13028 21794 13084
rect 21794 13028 21850 13084
rect 21850 13028 21854 13084
rect 21790 13024 21854 13028
rect 21870 13084 21934 13088
rect 21870 13028 21874 13084
rect 21874 13028 21930 13084
rect 21930 13028 21934 13084
rect 21870 13024 21934 13028
rect 21950 13084 22014 13088
rect 21950 13028 21954 13084
rect 21954 13028 22010 13084
rect 22010 13028 22014 13084
rect 21950 13024 22014 13028
rect 22030 13084 22094 13088
rect 22030 13028 22034 13084
rect 22034 13028 22090 13084
rect 22090 13028 22094 13084
rect 22030 13024 22094 13028
rect 28736 13084 28800 13088
rect 28736 13028 28740 13084
rect 28740 13028 28796 13084
rect 28796 13028 28800 13084
rect 28736 13024 28800 13028
rect 28816 13084 28880 13088
rect 28816 13028 28820 13084
rect 28820 13028 28876 13084
rect 28876 13028 28880 13084
rect 28816 13024 28880 13028
rect 28896 13084 28960 13088
rect 28896 13028 28900 13084
rect 28900 13028 28956 13084
rect 28956 13028 28960 13084
rect 28896 13024 28960 13028
rect 28976 13084 29040 13088
rect 28976 13028 28980 13084
rect 28980 13028 29036 13084
rect 29036 13028 29040 13084
rect 28976 13024 29040 13028
rect 4425 12540 4489 12544
rect 4425 12484 4429 12540
rect 4429 12484 4485 12540
rect 4485 12484 4489 12540
rect 4425 12480 4489 12484
rect 4505 12540 4569 12544
rect 4505 12484 4509 12540
rect 4509 12484 4565 12540
rect 4565 12484 4569 12540
rect 4505 12480 4569 12484
rect 4585 12540 4649 12544
rect 4585 12484 4589 12540
rect 4589 12484 4645 12540
rect 4645 12484 4649 12540
rect 4585 12480 4649 12484
rect 4665 12540 4729 12544
rect 4665 12484 4669 12540
rect 4669 12484 4725 12540
rect 4725 12484 4729 12540
rect 4665 12480 4729 12484
rect 11371 12540 11435 12544
rect 11371 12484 11375 12540
rect 11375 12484 11431 12540
rect 11431 12484 11435 12540
rect 11371 12480 11435 12484
rect 11451 12540 11515 12544
rect 11451 12484 11455 12540
rect 11455 12484 11511 12540
rect 11511 12484 11515 12540
rect 11451 12480 11515 12484
rect 11531 12540 11595 12544
rect 11531 12484 11535 12540
rect 11535 12484 11591 12540
rect 11591 12484 11595 12540
rect 11531 12480 11595 12484
rect 11611 12540 11675 12544
rect 11611 12484 11615 12540
rect 11615 12484 11671 12540
rect 11671 12484 11675 12540
rect 11611 12480 11675 12484
rect 18317 12540 18381 12544
rect 18317 12484 18321 12540
rect 18321 12484 18377 12540
rect 18377 12484 18381 12540
rect 18317 12480 18381 12484
rect 18397 12540 18461 12544
rect 18397 12484 18401 12540
rect 18401 12484 18457 12540
rect 18457 12484 18461 12540
rect 18397 12480 18461 12484
rect 18477 12540 18541 12544
rect 18477 12484 18481 12540
rect 18481 12484 18537 12540
rect 18537 12484 18541 12540
rect 18477 12480 18541 12484
rect 18557 12540 18621 12544
rect 18557 12484 18561 12540
rect 18561 12484 18617 12540
rect 18617 12484 18621 12540
rect 18557 12480 18621 12484
rect 25263 12540 25327 12544
rect 25263 12484 25267 12540
rect 25267 12484 25323 12540
rect 25323 12484 25327 12540
rect 25263 12480 25327 12484
rect 25343 12540 25407 12544
rect 25343 12484 25347 12540
rect 25347 12484 25403 12540
rect 25403 12484 25407 12540
rect 25343 12480 25407 12484
rect 25423 12540 25487 12544
rect 25423 12484 25427 12540
rect 25427 12484 25483 12540
rect 25483 12484 25487 12540
rect 25423 12480 25487 12484
rect 25503 12540 25567 12544
rect 25503 12484 25507 12540
rect 25507 12484 25563 12540
rect 25563 12484 25567 12540
rect 25503 12480 25567 12484
rect 7898 11996 7962 12000
rect 7898 11940 7902 11996
rect 7902 11940 7958 11996
rect 7958 11940 7962 11996
rect 7898 11936 7962 11940
rect 7978 11996 8042 12000
rect 7978 11940 7982 11996
rect 7982 11940 8038 11996
rect 8038 11940 8042 11996
rect 7978 11936 8042 11940
rect 8058 11996 8122 12000
rect 8058 11940 8062 11996
rect 8062 11940 8118 11996
rect 8118 11940 8122 11996
rect 8058 11936 8122 11940
rect 8138 11996 8202 12000
rect 8138 11940 8142 11996
rect 8142 11940 8198 11996
rect 8198 11940 8202 11996
rect 8138 11936 8202 11940
rect 14844 11996 14908 12000
rect 14844 11940 14848 11996
rect 14848 11940 14904 11996
rect 14904 11940 14908 11996
rect 14844 11936 14908 11940
rect 14924 11996 14988 12000
rect 14924 11940 14928 11996
rect 14928 11940 14984 11996
rect 14984 11940 14988 11996
rect 14924 11936 14988 11940
rect 15004 11996 15068 12000
rect 15004 11940 15008 11996
rect 15008 11940 15064 11996
rect 15064 11940 15068 11996
rect 15004 11936 15068 11940
rect 15084 11996 15148 12000
rect 15084 11940 15088 11996
rect 15088 11940 15144 11996
rect 15144 11940 15148 11996
rect 15084 11936 15148 11940
rect 21790 11996 21854 12000
rect 21790 11940 21794 11996
rect 21794 11940 21850 11996
rect 21850 11940 21854 11996
rect 21790 11936 21854 11940
rect 21870 11996 21934 12000
rect 21870 11940 21874 11996
rect 21874 11940 21930 11996
rect 21930 11940 21934 11996
rect 21870 11936 21934 11940
rect 21950 11996 22014 12000
rect 21950 11940 21954 11996
rect 21954 11940 22010 11996
rect 22010 11940 22014 11996
rect 21950 11936 22014 11940
rect 22030 11996 22094 12000
rect 22030 11940 22034 11996
rect 22034 11940 22090 11996
rect 22090 11940 22094 11996
rect 22030 11936 22094 11940
rect 28736 11996 28800 12000
rect 28736 11940 28740 11996
rect 28740 11940 28796 11996
rect 28796 11940 28800 11996
rect 28736 11936 28800 11940
rect 28816 11996 28880 12000
rect 28816 11940 28820 11996
rect 28820 11940 28876 11996
rect 28876 11940 28880 11996
rect 28816 11936 28880 11940
rect 28896 11996 28960 12000
rect 28896 11940 28900 11996
rect 28900 11940 28956 11996
rect 28956 11940 28960 11996
rect 28896 11936 28960 11940
rect 28976 11996 29040 12000
rect 28976 11940 28980 11996
rect 28980 11940 29036 11996
rect 29036 11940 29040 11996
rect 28976 11936 29040 11940
rect 4425 11452 4489 11456
rect 4425 11396 4429 11452
rect 4429 11396 4485 11452
rect 4485 11396 4489 11452
rect 4425 11392 4489 11396
rect 4505 11452 4569 11456
rect 4505 11396 4509 11452
rect 4509 11396 4565 11452
rect 4565 11396 4569 11452
rect 4505 11392 4569 11396
rect 4585 11452 4649 11456
rect 4585 11396 4589 11452
rect 4589 11396 4645 11452
rect 4645 11396 4649 11452
rect 4585 11392 4649 11396
rect 4665 11452 4729 11456
rect 4665 11396 4669 11452
rect 4669 11396 4725 11452
rect 4725 11396 4729 11452
rect 4665 11392 4729 11396
rect 11371 11452 11435 11456
rect 11371 11396 11375 11452
rect 11375 11396 11431 11452
rect 11431 11396 11435 11452
rect 11371 11392 11435 11396
rect 11451 11452 11515 11456
rect 11451 11396 11455 11452
rect 11455 11396 11511 11452
rect 11511 11396 11515 11452
rect 11451 11392 11515 11396
rect 11531 11452 11595 11456
rect 11531 11396 11535 11452
rect 11535 11396 11591 11452
rect 11591 11396 11595 11452
rect 11531 11392 11595 11396
rect 11611 11452 11675 11456
rect 11611 11396 11615 11452
rect 11615 11396 11671 11452
rect 11671 11396 11675 11452
rect 11611 11392 11675 11396
rect 18317 11452 18381 11456
rect 18317 11396 18321 11452
rect 18321 11396 18377 11452
rect 18377 11396 18381 11452
rect 18317 11392 18381 11396
rect 18397 11452 18461 11456
rect 18397 11396 18401 11452
rect 18401 11396 18457 11452
rect 18457 11396 18461 11452
rect 18397 11392 18461 11396
rect 18477 11452 18541 11456
rect 18477 11396 18481 11452
rect 18481 11396 18537 11452
rect 18537 11396 18541 11452
rect 18477 11392 18541 11396
rect 18557 11452 18621 11456
rect 18557 11396 18561 11452
rect 18561 11396 18617 11452
rect 18617 11396 18621 11452
rect 18557 11392 18621 11396
rect 25263 11452 25327 11456
rect 25263 11396 25267 11452
rect 25267 11396 25323 11452
rect 25323 11396 25327 11452
rect 25263 11392 25327 11396
rect 25343 11452 25407 11456
rect 25343 11396 25347 11452
rect 25347 11396 25403 11452
rect 25403 11396 25407 11452
rect 25343 11392 25407 11396
rect 25423 11452 25487 11456
rect 25423 11396 25427 11452
rect 25427 11396 25483 11452
rect 25483 11396 25487 11452
rect 25423 11392 25487 11396
rect 25503 11452 25567 11456
rect 25503 11396 25507 11452
rect 25507 11396 25563 11452
rect 25563 11396 25567 11452
rect 25503 11392 25567 11396
rect 7898 10908 7962 10912
rect 7898 10852 7902 10908
rect 7902 10852 7958 10908
rect 7958 10852 7962 10908
rect 7898 10848 7962 10852
rect 7978 10908 8042 10912
rect 7978 10852 7982 10908
rect 7982 10852 8038 10908
rect 8038 10852 8042 10908
rect 7978 10848 8042 10852
rect 8058 10908 8122 10912
rect 8058 10852 8062 10908
rect 8062 10852 8118 10908
rect 8118 10852 8122 10908
rect 8058 10848 8122 10852
rect 8138 10908 8202 10912
rect 8138 10852 8142 10908
rect 8142 10852 8198 10908
rect 8198 10852 8202 10908
rect 8138 10848 8202 10852
rect 14844 10908 14908 10912
rect 14844 10852 14848 10908
rect 14848 10852 14904 10908
rect 14904 10852 14908 10908
rect 14844 10848 14908 10852
rect 14924 10908 14988 10912
rect 14924 10852 14928 10908
rect 14928 10852 14984 10908
rect 14984 10852 14988 10908
rect 14924 10848 14988 10852
rect 15004 10908 15068 10912
rect 15004 10852 15008 10908
rect 15008 10852 15064 10908
rect 15064 10852 15068 10908
rect 15004 10848 15068 10852
rect 15084 10908 15148 10912
rect 15084 10852 15088 10908
rect 15088 10852 15144 10908
rect 15144 10852 15148 10908
rect 15084 10848 15148 10852
rect 21790 10908 21854 10912
rect 21790 10852 21794 10908
rect 21794 10852 21850 10908
rect 21850 10852 21854 10908
rect 21790 10848 21854 10852
rect 21870 10908 21934 10912
rect 21870 10852 21874 10908
rect 21874 10852 21930 10908
rect 21930 10852 21934 10908
rect 21870 10848 21934 10852
rect 21950 10908 22014 10912
rect 21950 10852 21954 10908
rect 21954 10852 22010 10908
rect 22010 10852 22014 10908
rect 21950 10848 22014 10852
rect 22030 10908 22094 10912
rect 22030 10852 22034 10908
rect 22034 10852 22090 10908
rect 22090 10852 22094 10908
rect 22030 10848 22094 10852
rect 28736 10908 28800 10912
rect 28736 10852 28740 10908
rect 28740 10852 28796 10908
rect 28796 10852 28800 10908
rect 28736 10848 28800 10852
rect 28816 10908 28880 10912
rect 28816 10852 28820 10908
rect 28820 10852 28876 10908
rect 28876 10852 28880 10908
rect 28816 10848 28880 10852
rect 28896 10908 28960 10912
rect 28896 10852 28900 10908
rect 28900 10852 28956 10908
rect 28956 10852 28960 10908
rect 28896 10848 28960 10852
rect 28976 10908 29040 10912
rect 28976 10852 28980 10908
rect 28980 10852 29036 10908
rect 29036 10852 29040 10908
rect 28976 10848 29040 10852
rect 4425 10364 4489 10368
rect 4425 10308 4429 10364
rect 4429 10308 4485 10364
rect 4485 10308 4489 10364
rect 4425 10304 4489 10308
rect 4505 10364 4569 10368
rect 4505 10308 4509 10364
rect 4509 10308 4565 10364
rect 4565 10308 4569 10364
rect 4505 10304 4569 10308
rect 4585 10364 4649 10368
rect 4585 10308 4589 10364
rect 4589 10308 4645 10364
rect 4645 10308 4649 10364
rect 4585 10304 4649 10308
rect 4665 10364 4729 10368
rect 4665 10308 4669 10364
rect 4669 10308 4725 10364
rect 4725 10308 4729 10364
rect 4665 10304 4729 10308
rect 11371 10364 11435 10368
rect 11371 10308 11375 10364
rect 11375 10308 11431 10364
rect 11431 10308 11435 10364
rect 11371 10304 11435 10308
rect 11451 10364 11515 10368
rect 11451 10308 11455 10364
rect 11455 10308 11511 10364
rect 11511 10308 11515 10364
rect 11451 10304 11515 10308
rect 11531 10364 11595 10368
rect 11531 10308 11535 10364
rect 11535 10308 11591 10364
rect 11591 10308 11595 10364
rect 11531 10304 11595 10308
rect 11611 10364 11675 10368
rect 11611 10308 11615 10364
rect 11615 10308 11671 10364
rect 11671 10308 11675 10364
rect 11611 10304 11675 10308
rect 18317 10364 18381 10368
rect 18317 10308 18321 10364
rect 18321 10308 18377 10364
rect 18377 10308 18381 10364
rect 18317 10304 18381 10308
rect 18397 10364 18461 10368
rect 18397 10308 18401 10364
rect 18401 10308 18457 10364
rect 18457 10308 18461 10364
rect 18397 10304 18461 10308
rect 18477 10364 18541 10368
rect 18477 10308 18481 10364
rect 18481 10308 18537 10364
rect 18537 10308 18541 10364
rect 18477 10304 18541 10308
rect 18557 10364 18621 10368
rect 18557 10308 18561 10364
rect 18561 10308 18617 10364
rect 18617 10308 18621 10364
rect 18557 10304 18621 10308
rect 25263 10364 25327 10368
rect 25263 10308 25267 10364
rect 25267 10308 25323 10364
rect 25323 10308 25327 10364
rect 25263 10304 25327 10308
rect 25343 10364 25407 10368
rect 25343 10308 25347 10364
rect 25347 10308 25403 10364
rect 25403 10308 25407 10364
rect 25343 10304 25407 10308
rect 25423 10364 25487 10368
rect 25423 10308 25427 10364
rect 25427 10308 25483 10364
rect 25483 10308 25487 10364
rect 25423 10304 25487 10308
rect 25503 10364 25567 10368
rect 25503 10308 25507 10364
rect 25507 10308 25563 10364
rect 25563 10308 25567 10364
rect 25503 10304 25567 10308
rect 7898 9820 7962 9824
rect 7898 9764 7902 9820
rect 7902 9764 7958 9820
rect 7958 9764 7962 9820
rect 7898 9760 7962 9764
rect 7978 9820 8042 9824
rect 7978 9764 7982 9820
rect 7982 9764 8038 9820
rect 8038 9764 8042 9820
rect 7978 9760 8042 9764
rect 8058 9820 8122 9824
rect 8058 9764 8062 9820
rect 8062 9764 8118 9820
rect 8118 9764 8122 9820
rect 8058 9760 8122 9764
rect 8138 9820 8202 9824
rect 8138 9764 8142 9820
rect 8142 9764 8198 9820
rect 8198 9764 8202 9820
rect 8138 9760 8202 9764
rect 14844 9820 14908 9824
rect 14844 9764 14848 9820
rect 14848 9764 14904 9820
rect 14904 9764 14908 9820
rect 14844 9760 14908 9764
rect 14924 9820 14988 9824
rect 14924 9764 14928 9820
rect 14928 9764 14984 9820
rect 14984 9764 14988 9820
rect 14924 9760 14988 9764
rect 15004 9820 15068 9824
rect 15004 9764 15008 9820
rect 15008 9764 15064 9820
rect 15064 9764 15068 9820
rect 15004 9760 15068 9764
rect 15084 9820 15148 9824
rect 15084 9764 15088 9820
rect 15088 9764 15144 9820
rect 15144 9764 15148 9820
rect 15084 9760 15148 9764
rect 21790 9820 21854 9824
rect 21790 9764 21794 9820
rect 21794 9764 21850 9820
rect 21850 9764 21854 9820
rect 21790 9760 21854 9764
rect 21870 9820 21934 9824
rect 21870 9764 21874 9820
rect 21874 9764 21930 9820
rect 21930 9764 21934 9820
rect 21870 9760 21934 9764
rect 21950 9820 22014 9824
rect 21950 9764 21954 9820
rect 21954 9764 22010 9820
rect 22010 9764 22014 9820
rect 21950 9760 22014 9764
rect 22030 9820 22094 9824
rect 22030 9764 22034 9820
rect 22034 9764 22090 9820
rect 22090 9764 22094 9820
rect 22030 9760 22094 9764
rect 28736 9820 28800 9824
rect 28736 9764 28740 9820
rect 28740 9764 28796 9820
rect 28796 9764 28800 9820
rect 28736 9760 28800 9764
rect 28816 9820 28880 9824
rect 28816 9764 28820 9820
rect 28820 9764 28876 9820
rect 28876 9764 28880 9820
rect 28816 9760 28880 9764
rect 28896 9820 28960 9824
rect 28896 9764 28900 9820
rect 28900 9764 28956 9820
rect 28956 9764 28960 9820
rect 28896 9760 28960 9764
rect 28976 9820 29040 9824
rect 28976 9764 28980 9820
rect 28980 9764 29036 9820
rect 29036 9764 29040 9820
rect 28976 9760 29040 9764
rect 4425 9276 4489 9280
rect 4425 9220 4429 9276
rect 4429 9220 4485 9276
rect 4485 9220 4489 9276
rect 4425 9216 4489 9220
rect 4505 9276 4569 9280
rect 4505 9220 4509 9276
rect 4509 9220 4565 9276
rect 4565 9220 4569 9276
rect 4505 9216 4569 9220
rect 4585 9276 4649 9280
rect 4585 9220 4589 9276
rect 4589 9220 4645 9276
rect 4645 9220 4649 9276
rect 4585 9216 4649 9220
rect 4665 9276 4729 9280
rect 4665 9220 4669 9276
rect 4669 9220 4725 9276
rect 4725 9220 4729 9276
rect 4665 9216 4729 9220
rect 11371 9276 11435 9280
rect 11371 9220 11375 9276
rect 11375 9220 11431 9276
rect 11431 9220 11435 9276
rect 11371 9216 11435 9220
rect 11451 9276 11515 9280
rect 11451 9220 11455 9276
rect 11455 9220 11511 9276
rect 11511 9220 11515 9276
rect 11451 9216 11515 9220
rect 11531 9276 11595 9280
rect 11531 9220 11535 9276
rect 11535 9220 11591 9276
rect 11591 9220 11595 9276
rect 11531 9216 11595 9220
rect 11611 9276 11675 9280
rect 11611 9220 11615 9276
rect 11615 9220 11671 9276
rect 11671 9220 11675 9276
rect 11611 9216 11675 9220
rect 18317 9276 18381 9280
rect 18317 9220 18321 9276
rect 18321 9220 18377 9276
rect 18377 9220 18381 9276
rect 18317 9216 18381 9220
rect 18397 9276 18461 9280
rect 18397 9220 18401 9276
rect 18401 9220 18457 9276
rect 18457 9220 18461 9276
rect 18397 9216 18461 9220
rect 18477 9276 18541 9280
rect 18477 9220 18481 9276
rect 18481 9220 18537 9276
rect 18537 9220 18541 9276
rect 18477 9216 18541 9220
rect 18557 9276 18621 9280
rect 18557 9220 18561 9276
rect 18561 9220 18617 9276
rect 18617 9220 18621 9276
rect 18557 9216 18621 9220
rect 25263 9276 25327 9280
rect 25263 9220 25267 9276
rect 25267 9220 25323 9276
rect 25323 9220 25327 9276
rect 25263 9216 25327 9220
rect 25343 9276 25407 9280
rect 25343 9220 25347 9276
rect 25347 9220 25403 9276
rect 25403 9220 25407 9276
rect 25343 9216 25407 9220
rect 25423 9276 25487 9280
rect 25423 9220 25427 9276
rect 25427 9220 25483 9276
rect 25483 9220 25487 9276
rect 25423 9216 25487 9220
rect 25503 9276 25567 9280
rect 25503 9220 25507 9276
rect 25507 9220 25563 9276
rect 25563 9220 25567 9276
rect 25503 9216 25567 9220
rect 7898 8732 7962 8736
rect 7898 8676 7902 8732
rect 7902 8676 7958 8732
rect 7958 8676 7962 8732
rect 7898 8672 7962 8676
rect 7978 8732 8042 8736
rect 7978 8676 7982 8732
rect 7982 8676 8038 8732
rect 8038 8676 8042 8732
rect 7978 8672 8042 8676
rect 8058 8732 8122 8736
rect 8058 8676 8062 8732
rect 8062 8676 8118 8732
rect 8118 8676 8122 8732
rect 8058 8672 8122 8676
rect 8138 8732 8202 8736
rect 8138 8676 8142 8732
rect 8142 8676 8198 8732
rect 8198 8676 8202 8732
rect 8138 8672 8202 8676
rect 14844 8732 14908 8736
rect 14844 8676 14848 8732
rect 14848 8676 14904 8732
rect 14904 8676 14908 8732
rect 14844 8672 14908 8676
rect 14924 8732 14988 8736
rect 14924 8676 14928 8732
rect 14928 8676 14984 8732
rect 14984 8676 14988 8732
rect 14924 8672 14988 8676
rect 15004 8732 15068 8736
rect 15004 8676 15008 8732
rect 15008 8676 15064 8732
rect 15064 8676 15068 8732
rect 15004 8672 15068 8676
rect 15084 8732 15148 8736
rect 15084 8676 15088 8732
rect 15088 8676 15144 8732
rect 15144 8676 15148 8732
rect 15084 8672 15148 8676
rect 21790 8732 21854 8736
rect 21790 8676 21794 8732
rect 21794 8676 21850 8732
rect 21850 8676 21854 8732
rect 21790 8672 21854 8676
rect 21870 8732 21934 8736
rect 21870 8676 21874 8732
rect 21874 8676 21930 8732
rect 21930 8676 21934 8732
rect 21870 8672 21934 8676
rect 21950 8732 22014 8736
rect 21950 8676 21954 8732
rect 21954 8676 22010 8732
rect 22010 8676 22014 8732
rect 21950 8672 22014 8676
rect 22030 8732 22094 8736
rect 22030 8676 22034 8732
rect 22034 8676 22090 8732
rect 22090 8676 22094 8732
rect 22030 8672 22094 8676
rect 28736 8732 28800 8736
rect 28736 8676 28740 8732
rect 28740 8676 28796 8732
rect 28796 8676 28800 8732
rect 28736 8672 28800 8676
rect 28816 8732 28880 8736
rect 28816 8676 28820 8732
rect 28820 8676 28876 8732
rect 28876 8676 28880 8732
rect 28816 8672 28880 8676
rect 28896 8732 28960 8736
rect 28896 8676 28900 8732
rect 28900 8676 28956 8732
rect 28956 8676 28960 8732
rect 28896 8672 28960 8676
rect 28976 8732 29040 8736
rect 28976 8676 28980 8732
rect 28980 8676 29036 8732
rect 29036 8676 29040 8732
rect 28976 8672 29040 8676
rect 4425 8188 4489 8192
rect 4425 8132 4429 8188
rect 4429 8132 4485 8188
rect 4485 8132 4489 8188
rect 4425 8128 4489 8132
rect 4505 8188 4569 8192
rect 4505 8132 4509 8188
rect 4509 8132 4565 8188
rect 4565 8132 4569 8188
rect 4505 8128 4569 8132
rect 4585 8188 4649 8192
rect 4585 8132 4589 8188
rect 4589 8132 4645 8188
rect 4645 8132 4649 8188
rect 4585 8128 4649 8132
rect 4665 8188 4729 8192
rect 4665 8132 4669 8188
rect 4669 8132 4725 8188
rect 4725 8132 4729 8188
rect 4665 8128 4729 8132
rect 11371 8188 11435 8192
rect 11371 8132 11375 8188
rect 11375 8132 11431 8188
rect 11431 8132 11435 8188
rect 11371 8128 11435 8132
rect 11451 8188 11515 8192
rect 11451 8132 11455 8188
rect 11455 8132 11511 8188
rect 11511 8132 11515 8188
rect 11451 8128 11515 8132
rect 11531 8188 11595 8192
rect 11531 8132 11535 8188
rect 11535 8132 11591 8188
rect 11591 8132 11595 8188
rect 11531 8128 11595 8132
rect 11611 8188 11675 8192
rect 11611 8132 11615 8188
rect 11615 8132 11671 8188
rect 11671 8132 11675 8188
rect 11611 8128 11675 8132
rect 18317 8188 18381 8192
rect 18317 8132 18321 8188
rect 18321 8132 18377 8188
rect 18377 8132 18381 8188
rect 18317 8128 18381 8132
rect 18397 8188 18461 8192
rect 18397 8132 18401 8188
rect 18401 8132 18457 8188
rect 18457 8132 18461 8188
rect 18397 8128 18461 8132
rect 18477 8188 18541 8192
rect 18477 8132 18481 8188
rect 18481 8132 18537 8188
rect 18537 8132 18541 8188
rect 18477 8128 18541 8132
rect 18557 8188 18621 8192
rect 18557 8132 18561 8188
rect 18561 8132 18617 8188
rect 18617 8132 18621 8188
rect 18557 8128 18621 8132
rect 25263 8188 25327 8192
rect 25263 8132 25267 8188
rect 25267 8132 25323 8188
rect 25323 8132 25327 8188
rect 25263 8128 25327 8132
rect 25343 8188 25407 8192
rect 25343 8132 25347 8188
rect 25347 8132 25403 8188
rect 25403 8132 25407 8188
rect 25343 8128 25407 8132
rect 25423 8188 25487 8192
rect 25423 8132 25427 8188
rect 25427 8132 25483 8188
rect 25483 8132 25487 8188
rect 25423 8128 25487 8132
rect 25503 8188 25567 8192
rect 25503 8132 25507 8188
rect 25507 8132 25563 8188
rect 25563 8132 25567 8188
rect 25503 8128 25567 8132
rect 7898 7644 7962 7648
rect 7898 7588 7902 7644
rect 7902 7588 7958 7644
rect 7958 7588 7962 7644
rect 7898 7584 7962 7588
rect 7978 7644 8042 7648
rect 7978 7588 7982 7644
rect 7982 7588 8038 7644
rect 8038 7588 8042 7644
rect 7978 7584 8042 7588
rect 8058 7644 8122 7648
rect 8058 7588 8062 7644
rect 8062 7588 8118 7644
rect 8118 7588 8122 7644
rect 8058 7584 8122 7588
rect 8138 7644 8202 7648
rect 8138 7588 8142 7644
rect 8142 7588 8198 7644
rect 8198 7588 8202 7644
rect 8138 7584 8202 7588
rect 14844 7644 14908 7648
rect 14844 7588 14848 7644
rect 14848 7588 14904 7644
rect 14904 7588 14908 7644
rect 14844 7584 14908 7588
rect 14924 7644 14988 7648
rect 14924 7588 14928 7644
rect 14928 7588 14984 7644
rect 14984 7588 14988 7644
rect 14924 7584 14988 7588
rect 15004 7644 15068 7648
rect 15004 7588 15008 7644
rect 15008 7588 15064 7644
rect 15064 7588 15068 7644
rect 15004 7584 15068 7588
rect 15084 7644 15148 7648
rect 15084 7588 15088 7644
rect 15088 7588 15144 7644
rect 15144 7588 15148 7644
rect 15084 7584 15148 7588
rect 21790 7644 21854 7648
rect 21790 7588 21794 7644
rect 21794 7588 21850 7644
rect 21850 7588 21854 7644
rect 21790 7584 21854 7588
rect 21870 7644 21934 7648
rect 21870 7588 21874 7644
rect 21874 7588 21930 7644
rect 21930 7588 21934 7644
rect 21870 7584 21934 7588
rect 21950 7644 22014 7648
rect 21950 7588 21954 7644
rect 21954 7588 22010 7644
rect 22010 7588 22014 7644
rect 21950 7584 22014 7588
rect 22030 7644 22094 7648
rect 22030 7588 22034 7644
rect 22034 7588 22090 7644
rect 22090 7588 22094 7644
rect 22030 7584 22094 7588
rect 28736 7644 28800 7648
rect 28736 7588 28740 7644
rect 28740 7588 28796 7644
rect 28796 7588 28800 7644
rect 28736 7584 28800 7588
rect 28816 7644 28880 7648
rect 28816 7588 28820 7644
rect 28820 7588 28876 7644
rect 28876 7588 28880 7644
rect 28816 7584 28880 7588
rect 28896 7644 28960 7648
rect 28896 7588 28900 7644
rect 28900 7588 28956 7644
rect 28956 7588 28960 7644
rect 28896 7584 28960 7588
rect 28976 7644 29040 7648
rect 28976 7588 28980 7644
rect 28980 7588 29036 7644
rect 29036 7588 29040 7644
rect 28976 7584 29040 7588
rect 4425 7100 4489 7104
rect 4425 7044 4429 7100
rect 4429 7044 4485 7100
rect 4485 7044 4489 7100
rect 4425 7040 4489 7044
rect 4505 7100 4569 7104
rect 4505 7044 4509 7100
rect 4509 7044 4565 7100
rect 4565 7044 4569 7100
rect 4505 7040 4569 7044
rect 4585 7100 4649 7104
rect 4585 7044 4589 7100
rect 4589 7044 4645 7100
rect 4645 7044 4649 7100
rect 4585 7040 4649 7044
rect 4665 7100 4729 7104
rect 4665 7044 4669 7100
rect 4669 7044 4725 7100
rect 4725 7044 4729 7100
rect 4665 7040 4729 7044
rect 11371 7100 11435 7104
rect 11371 7044 11375 7100
rect 11375 7044 11431 7100
rect 11431 7044 11435 7100
rect 11371 7040 11435 7044
rect 11451 7100 11515 7104
rect 11451 7044 11455 7100
rect 11455 7044 11511 7100
rect 11511 7044 11515 7100
rect 11451 7040 11515 7044
rect 11531 7100 11595 7104
rect 11531 7044 11535 7100
rect 11535 7044 11591 7100
rect 11591 7044 11595 7100
rect 11531 7040 11595 7044
rect 11611 7100 11675 7104
rect 11611 7044 11615 7100
rect 11615 7044 11671 7100
rect 11671 7044 11675 7100
rect 11611 7040 11675 7044
rect 18317 7100 18381 7104
rect 18317 7044 18321 7100
rect 18321 7044 18377 7100
rect 18377 7044 18381 7100
rect 18317 7040 18381 7044
rect 18397 7100 18461 7104
rect 18397 7044 18401 7100
rect 18401 7044 18457 7100
rect 18457 7044 18461 7100
rect 18397 7040 18461 7044
rect 18477 7100 18541 7104
rect 18477 7044 18481 7100
rect 18481 7044 18537 7100
rect 18537 7044 18541 7100
rect 18477 7040 18541 7044
rect 18557 7100 18621 7104
rect 18557 7044 18561 7100
rect 18561 7044 18617 7100
rect 18617 7044 18621 7100
rect 18557 7040 18621 7044
rect 25263 7100 25327 7104
rect 25263 7044 25267 7100
rect 25267 7044 25323 7100
rect 25323 7044 25327 7100
rect 25263 7040 25327 7044
rect 25343 7100 25407 7104
rect 25343 7044 25347 7100
rect 25347 7044 25403 7100
rect 25403 7044 25407 7100
rect 25343 7040 25407 7044
rect 25423 7100 25487 7104
rect 25423 7044 25427 7100
rect 25427 7044 25483 7100
rect 25483 7044 25487 7100
rect 25423 7040 25487 7044
rect 25503 7100 25567 7104
rect 25503 7044 25507 7100
rect 25507 7044 25563 7100
rect 25563 7044 25567 7100
rect 25503 7040 25567 7044
rect 7898 6556 7962 6560
rect 7898 6500 7902 6556
rect 7902 6500 7958 6556
rect 7958 6500 7962 6556
rect 7898 6496 7962 6500
rect 7978 6556 8042 6560
rect 7978 6500 7982 6556
rect 7982 6500 8038 6556
rect 8038 6500 8042 6556
rect 7978 6496 8042 6500
rect 8058 6556 8122 6560
rect 8058 6500 8062 6556
rect 8062 6500 8118 6556
rect 8118 6500 8122 6556
rect 8058 6496 8122 6500
rect 8138 6556 8202 6560
rect 8138 6500 8142 6556
rect 8142 6500 8198 6556
rect 8198 6500 8202 6556
rect 8138 6496 8202 6500
rect 14844 6556 14908 6560
rect 14844 6500 14848 6556
rect 14848 6500 14904 6556
rect 14904 6500 14908 6556
rect 14844 6496 14908 6500
rect 14924 6556 14988 6560
rect 14924 6500 14928 6556
rect 14928 6500 14984 6556
rect 14984 6500 14988 6556
rect 14924 6496 14988 6500
rect 15004 6556 15068 6560
rect 15004 6500 15008 6556
rect 15008 6500 15064 6556
rect 15064 6500 15068 6556
rect 15004 6496 15068 6500
rect 15084 6556 15148 6560
rect 15084 6500 15088 6556
rect 15088 6500 15144 6556
rect 15144 6500 15148 6556
rect 15084 6496 15148 6500
rect 21790 6556 21854 6560
rect 21790 6500 21794 6556
rect 21794 6500 21850 6556
rect 21850 6500 21854 6556
rect 21790 6496 21854 6500
rect 21870 6556 21934 6560
rect 21870 6500 21874 6556
rect 21874 6500 21930 6556
rect 21930 6500 21934 6556
rect 21870 6496 21934 6500
rect 21950 6556 22014 6560
rect 21950 6500 21954 6556
rect 21954 6500 22010 6556
rect 22010 6500 22014 6556
rect 21950 6496 22014 6500
rect 22030 6556 22094 6560
rect 22030 6500 22034 6556
rect 22034 6500 22090 6556
rect 22090 6500 22094 6556
rect 22030 6496 22094 6500
rect 28736 6556 28800 6560
rect 28736 6500 28740 6556
rect 28740 6500 28796 6556
rect 28796 6500 28800 6556
rect 28736 6496 28800 6500
rect 28816 6556 28880 6560
rect 28816 6500 28820 6556
rect 28820 6500 28876 6556
rect 28876 6500 28880 6556
rect 28816 6496 28880 6500
rect 28896 6556 28960 6560
rect 28896 6500 28900 6556
rect 28900 6500 28956 6556
rect 28956 6500 28960 6556
rect 28896 6496 28960 6500
rect 28976 6556 29040 6560
rect 28976 6500 28980 6556
rect 28980 6500 29036 6556
rect 29036 6500 29040 6556
rect 28976 6496 29040 6500
rect 4425 6012 4489 6016
rect 4425 5956 4429 6012
rect 4429 5956 4485 6012
rect 4485 5956 4489 6012
rect 4425 5952 4489 5956
rect 4505 6012 4569 6016
rect 4505 5956 4509 6012
rect 4509 5956 4565 6012
rect 4565 5956 4569 6012
rect 4505 5952 4569 5956
rect 4585 6012 4649 6016
rect 4585 5956 4589 6012
rect 4589 5956 4645 6012
rect 4645 5956 4649 6012
rect 4585 5952 4649 5956
rect 4665 6012 4729 6016
rect 4665 5956 4669 6012
rect 4669 5956 4725 6012
rect 4725 5956 4729 6012
rect 4665 5952 4729 5956
rect 11371 6012 11435 6016
rect 11371 5956 11375 6012
rect 11375 5956 11431 6012
rect 11431 5956 11435 6012
rect 11371 5952 11435 5956
rect 11451 6012 11515 6016
rect 11451 5956 11455 6012
rect 11455 5956 11511 6012
rect 11511 5956 11515 6012
rect 11451 5952 11515 5956
rect 11531 6012 11595 6016
rect 11531 5956 11535 6012
rect 11535 5956 11591 6012
rect 11591 5956 11595 6012
rect 11531 5952 11595 5956
rect 11611 6012 11675 6016
rect 11611 5956 11615 6012
rect 11615 5956 11671 6012
rect 11671 5956 11675 6012
rect 11611 5952 11675 5956
rect 18317 6012 18381 6016
rect 18317 5956 18321 6012
rect 18321 5956 18377 6012
rect 18377 5956 18381 6012
rect 18317 5952 18381 5956
rect 18397 6012 18461 6016
rect 18397 5956 18401 6012
rect 18401 5956 18457 6012
rect 18457 5956 18461 6012
rect 18397 5952 18461 5956
rect 18477 6012 18541 6016
rect 18477 5956 18481 6012
rect 18481 5956 18537 6012
rect 18537 5956 18541 6012
rect 18477 5952 18541 5956
rect 18557 6012 18621 6016
rect 18557 5956 18561 6012
rect 18561 5956 18617 6012
rect 18617 5956 18621 6012
rect 18557 5952 18621 5956
rect 25263 6012 25327 6016
rect 25263 5956 25267 6012
rect 25267 5956 25323 6012
rect 25323 5956 25327 6012
rect 25263 5952 25327 5956
rect 25343 6012 25407 6016
rect 25343 5956 25347 6012
rect 25347 5956 25403 6012
rect 25403 5956 25407 6012
rect 25343 5952 25407 5956
rect 25423 6012 25487 6016
rect 25423 5956 25427 6012
rect 25427 5956 25483 6012
rect 25483 5956 25487 6012
rect 25423 5952 25487 5956
rect 25503 6012 25567 6016
rect 25503 5956 25507 6012
rect 25507 5956 25563 6012
rect 25563 5956 25567 6012
rect 25503 5952 25567 5956
rect 7898 5468 7962 5472
rect 7898 5412 7902 5468
rect 7902 5412 7958 5468
rect 7958 5412 7962 5468
rect 7898 5408 7962 5412
rect 7978 5468 8042 5472
rect 7978 5412 7982 5468
rect 7982 5412 8038 5468
rect 8038 5412 8042 5468
rect 7978 5408 8042 5412
rect 8058 5468 8122 5472
rect 8058 5412 8062 5468
rect 8062 5412 8118 5468
rect 8118 5412 8122 5468
rect 8058 5408 8122 5412
rect 8138 5468 8202 5472
rect 8138 5412 8142 5468
rect 8142 5412 8198 5468
rect 8198 5412 8202 5468
rect 8138 5408 8202 5412
rect 14844 5468 14908 5472
rect 14844 5412 14848 5468
rect 14848 5412 14904 5468
rect 14904 5412 14908 5468
rect 14844 5408 14908 5412
rect 14924 5468 14988 5472
rect 14924 5412 14928 5468
rect 14928 5412 14984 5468
rect 14984 5412 14988 5468
rect 14924 5408 14988 5412
rect 15004 5468 15068 5472
rect 15004 5412 15008 5468
rect 15008 5412 15064 5468
rect 15064 5412 15068 5468
rect 15004 5408 15068 5412
rect 15084 5468 15148 5472
rect 15084 5412 15088 5468
rect 15088 5412 15144 5468
rect 15144 5412 15148 5468
rect 15084 5408 15148 5412
rect 21790 5468 21854 5472
rect 21790 5412 21794 5468
rect 21794 5412 21850 5468
rect 21850 5412 21854 5468
rect 21790 5408 21854 5412
rect 21870 5468 21934 5472
rect 21870 5412 21874 5468
rect 21874 5412 21930 5468
rect 21930 5412 21934 5468
rect 21870 5408 21934 5412
rect 21950 5468 22014 5472
rect 21950 5412 21954 5468
rect 21954 5412 22010 5468
rect 22010 5412 22014 5468
rect 21950 5408 22014 5412
rect 22030 5468 22094 5472
rect 22030 5412 22034 5468
rect 22034 5412 22090 5468
rect 22090 5412 22094 5468
rect 22030 5408 22094 5412
rect 28736 5468 28800 5472
rect 28736 5412 28740 5468
rect 28740 5412 28796 5468
rect 28796 5412 28800 5468
rect 28736 5408 28800 5412
rect 28816 5468 28880 5472
rect 28816 5412 28820 5468
rect 28820 5412 28876 5468
rect 28876 5412 28880 5468
rect 28816 5408 28880 5412
rect 28896 5468 28960 5472
rect 28896 5412 28900 5468
rect 28900 5412 28956 5468
rect 28956 5412 28960 5468
rect 28896 5408 28960 5412
rect 28976 5468 29040 5472
rect 28976 5412 28980 5468
rect 28980 5412 29036 5468
rect 29036 5412 29040 5468
rect 28976 5408 29040 5412
rect 4425 4924 4489 4928
rect 4425 4868 4429 4924
rect 4429 4868 4485 4924
rect 4485 4868 4489 4924
rect 4425 4864 4489 4868
rect 4505 4924 4569 4928
rect 4505 4868 4509 4924
rect 4509 4868 4565 4924
rect 4565 4868 4569 4924
rect 4505 4864 4569 4868
rect 4585 4924 4649 4928
rect 4585 4868 4589 4924
rect 4589 4868 4645 4924
rect 4645 4868 4649 4924
rect 4585 4864 4649 4868
rect 4665 4924 4729 4928
rect 4665 4868 4669 4924
rect 4669 4868 4725 4924
rect 4725 4868 4729 4924
rect 4665 4864 4729 4868
rect 11371 4924 11435 4928
rect 11371 4868 11375 4924
rect 11375 4868 11431 4924
rect 11431 4868 11435 4924
rect 11371 4864 11435 4868
rect 11451 4924 11515 4928
rect 11451 4868 11455 4924
rect 11455 4868 11511 4924
rect 11511 4868 11515 4924
rect 11451 4864 11515 4868
rect 11531 4924 11595 4928
rect 11531 4868 11535 4924
rect 11535 4868 11591 4924
rect 11591 4868 11595 4924
rect 11531 4864 11595 4868
rect 11611 4924 11675 4928
rect 11611 4868 11615 4924
rect 11615 4868 11671 4924
rect 11671 4868 11675 4924
rect 11611 4864 11675 4868
rect 18317 4924 18381 4928
rect 18317 4868 18321 4924
rect 18321 4868 18377 4924
rect 18377 4868 18381 4924
rect 18317 4864 18381 4868
rect 18397 4924 18461 4928
rect 18397 4868 18401 4924
rect 18401 4868 18457 4924
rect 18457 4868 18461 4924
rect 18397 4864 18461 4868
rect 18477 4924 18541 4928
rect 18477 4868 18481 4924
rect 18481 4868 18537 4924
rect 18537 4868 18541 4924
rect 18477 4864 18541 4868
rect 18557 4924 18621 4928
rect 18557 4868 18561 4924
rect 18561 4868 18617 4924
rect 18617 4868 18621 4924
rect 18557 4864 18621 4868
rect 25263 4924 25327 4928
rect 25263 4868 25267 4924
rect 25267 4868 25323 4924
rect 25323 4868 25327 4924
rect 25263 4864 25327 4868
rect 25343 4924 25407 4928
rect 25343 4868 25347 4924
rect 25347 4868 25403 4924
rect 25403 4868 25407 4924
rect 25343 4864 25407 4868
rect 25423 4924 25487 4928
rect 25423 4868 25427 4924
rect 25427 4868 25483 4924
rect 25483 4868 25487 4924
rect 25423 4864 25487 4868
rect 25503 4924 25567 4928
rect 25503 4868 25507 4924
rect 25507 4868 25563 4924
rect 25563 4868 25567 4924
rect 25503 4864 25567 4868
rect 7898 4380 7962 4384
rect 7898 4324 7902 4380
rect 7902 4324 7958 4380
rect 7958 4324 7962 4380
rect 7898 4320 7962 4324
rect 7978 4380 8042 4384
rect 7978 4324 7982 4380
rect 7982 4324 8038 4380
rect 8038 4324 8042 4380
rect 7978 4320 8042 4324
rect 8058 4380 8122 4384
rect 8058 4324 8062 4380
rect 8062 4324 8118 4380
rect 8118 4324 8122 4380
rect 8058 4320 8122 4324
rect 8138 4380 8202 4384
rect 8138 4324 8142 4380
rect 8142 4324 8198 4380
rect 8198 4324 8202 4380
rect 8138 4320 8202 4324
rect 14844 4380 14908 4384
rect 14844 4324 14848 4380
rect 14848 4324 14904 4380
rect 14904 4324 14908 4380
rect 14844 4320 14908 4324
rect 14924 4380 14988 4384
rect 14924 4324 14928 4380
rect 14928 4324 14984 4380
rect 14984 4324 14988 4380
rect 14924 4320 14988 4324
rect 15004 4380 15068 4384
rect 15004 4324 15008 4380
rect 15008 4324 15064 4380
rect 15064 4324 15068 4380
rect 15004 4320 15068 4324
rect 15084 4380 15148 4384
rect 15084 4324 15088 4380
rect 15088 4324 15144 4380
rect 15144 4324 15148 4380
rect 15084 4320 15148 4324
rect 21790 4380 21854 4384
rect 21790 4324 21794 4380
rect 21794 4324 21850 4380
rect 21850 4324 21854 4380
rect 21790 4320 21854 4324
rect 21870 4380 21934 4384
rect 21870 4324 21874 4380
rect 21874 4324 21930 4380
rect 21930 4324 21934 4380
rect 21870 4320 21934 4324
rect 21950 4380 22014 4384
rect 21950 4324 21954 4380
rect 21954 4324 22010 4380
rect 22010 4324 22014 4380
rect 21950 4320 22014 4324
rect 22030 4380 22094 4384
rect 22030 4324 22034 4380
rect 22034 4324 22090 4380
rect 22090 4324 22094 4380
rect 22030 4320 22094 4324
rect 28736 4380 28800 4384
rect 28736 4324 28740 4380
rect 28740 4324 28796 4380
rect 28796 4324 28800 4380
rect 28736 4320 28800 4324
rect 28816 4380 28880 4384
rect 28816 4324 28820 4380
rect 28820 4324 28876 4380
rect 28876 4324 28880 4380
rect 28816 4320 28880 4324
rect 28896 4380 28960 4384
rect 28896 4324 28900 4380
rect 28900 4324 28956 4380
rect 28956 4324 28960 4380
rect 28896 4320 28960 4324
rect 28976 4380 29040 4384
rect 28976 4324 28980 4380
rect 28980 4324 29036 4380
rect 29036 4324 29040 4380
rect 28976 4320 29040 4324
rect 4425 3836 4489 3840
rect 4425 3780 4429 3836
rect 4429 3780 4485 3836
rect 4485 3780 4489 3836
rect 4425 3776 4489 3780
rect 4505 3836 4569 3840
rect 4505 3780 4509 3836
rect 4509 3780 4565 3836
rect 4565 3780 4569 3836
rect 4505 3776 4569 3780
rect 4585 3836 4649 3840
rect 4585 3780 4589 3836
rect 4589 3780 4645 3836
rect 4645 3780 4649 3836
rect 4585 3776 4649 3780
rect 4665 3836 4729 3840
rect 4665 3780 4669 3836
rect 4669 3780 4725 3836
rect 4725 3780 4729 3836
rect 4665 3776 4729 3780
rect 11371 3836 11435 3840
rect 11371 3780 11375 3836
rect 11375 3780 11431 3836
rect 11431 3780 11435 3836
rect 11371 3776 11435 3780
rect 11451 3836 11515 3840
rect 11451 3780 11455 3836
rect 11455 3780 11511 3836
rect 11511 3780 11515 3836
rect 11451 3776 11515 3780
rect 11531 3836 11595 3840
rect 11531 3780 11535 3836
rect 11535 3780 11591 3836
rect 11591 3780 11595 3836
rect 11531 3776 11595 3780
rect 11611 3836 11675 3840
rect 11611 3780 11615 3836
rect 11615 3780 11671 3836
rect 11671 3780 11675 3836
rect 11611 3776 11675 3780
rect 18317 3836 18381 3840
rect 18317 3780 18321 3836
rect 18321 3780 18377 3836
rect 18377 3780 18381 3836
rect 18317 3776 18381 3780
rect 18397 3836 18461 3840
rect 18397 3780 18401 3836
rect 18401 3780 18457 3836
rect 18457 3780 18461 3836
rect 18397 3776 18461 3780
rect 18477 3836 18541 3840
rect 18477 3780 18481 3836
rect 18481 3780 18537 3836
rect 18537 3780 18541 3836
rect 18477 3776 18541 3780
rect 18557 3836 18621 3840
rect 18557 3780 18561 3836
rect 18561 3780 18617 3836
rect 18617 3780 18621 3836
rect 18557 3776 18621 3780
rect 25263 3836 25327 3840
rect 25263 3780 25267 3836
rect 25267 3780 25323 3836
rect 25323 3780 25327 3836
rect 25263 3776 25327 3780
rect 25343 3836 25407 3840
rect 25343 3780 25347 3836
rect 25347 3780 25403 3836
rect 25403 3780 25407 3836
rect 25343 3776 25407 3780
rect 25423 3836 25487 3840
rect 25423 3780 25427 3836
rect 25427 3780 25483 3836
rect 25483 3780 25487 3836
rect 25423 3776 25487 3780
rect 25503 3836 25567 3840
rect 25503 3780 25507 3836
rect 25507 3780 25563 3836
rect 25563 3780 25567 3836
rect 25503 3776 25567 3780
rect 7898 3292 7962 3296
rect 7898 3236 7902 3292
rect 7902 3236 7958 3292
rect 7958 3236 7962 3292
rect 7898 3232 7962 3236
rect 7978 3292 8042 3296
rect 7978 3236 7982 3292
rect 7982 3236 8038 3292
rect 8038 3236 8042 3292
rect 7978 3232 8042 3236
rect 8058 3292 8122 3296
rect 8058 3236 8062 3292
rect 8062 3236 8118 3292
rect 8118 3236 8122 3292
rect 8058 3232 8122 3236
rect 8138 3292 8202 3296
rect 8138 3236 8142 3292
rect 8142 3236 8198 3292
rect 8198 3236 8202 3292
rect 8138 3232 8202 3236
rect 14844 3292 14908 3296
rect 14844 3236 14848 3292
rect 14848 3236 14904 3292
rect 14904 3236 14908 3292
rect 14844 3232 14908 3236
rect 14924 3292 14988 3296
rect 14924 3236 14928 3292
rect 14928 3236 14984 3292
rect 14984 3236 14988 3292
rect 14924 3232 14988 3236
rect 15004 3292 15068 3296
rect 15004 3236 15008 3292
rect 15008 3236 15064 3292
rect 15064 3236 15068 3292
rect 15004 3232 15068 3236
rect 15084 3292 15148 3296
rect 15084 3236 15088 3292
rect 15088 3236 15144 3292
rect 15144 3236 15148 3292
rect 15084 3232 15148 3236
rect 21790 3292 21854 3296
rect 21790 3236 21794 3292
rect 21794 3236 21850 3292
rect 21850 3236 21854 3292
rect 21790 3232 21854 3236
rect 21870 3292 21934 3296
rect 21870 3236 21874 3292
rect 21874 3236 21930 3292
rect 21930 3236 21934 3292
rect 21870 3232 21934 3236
rect 21950 3292 22014 3296
rect 21950 3236 21954 3292
rect 21954 3236 22010 3292
rect 22010 3236 22014 3292
rect 21950 3232 22014 3236
rect 22030 3292 22094 3296
rect 22030 3236 22034 3292
rect 22034 3236 22090 3292
rect 22090 3236 22094 3292
rect 22030 3232 22094 3236
rect 28736 3292 28800 3296
rect 28736 3236 28740 3292
rect 28740 3236 28796 3292
rect 28796 3236 28800 3292
rect 28736 3232 28800 3236
rect 28816 3292 28880 3296
rect 28816 3236 28820 3292
rect 28820 3236 28876 3292
rect 28876 3236 28880 3292
rect 28816 3232 28880 3236
rect 28896 3292 28960 3296
rect 28896 3236 28900 3292
rect 28900 3236 28956 3292
rect 28956 3236 28960 3292
rect 28896 3232 28960 3236
rect 28976 3292 29040 3296
rect 28976 3236 28980 3292
rect 28980 3236 29036 3292
rect 29036 3236 29040 3292
rect 28976 3232 29040 3236
rect 4425 2748 4489 2752
rect 4425 2692 4429 2748
rect 4429 2692 4485 2748
rect 4485 2692 4489 2748
rect 4425 2688 4489 2692
rect 4505 2748 4569 2752
rect 4505 2692 4509 2748
rect 4509 2692 4565 2748
rect 4565 2692 4569 2748
rect 4505 2688 4569 2692
rect 4585 2748 4649 2752
rect 4585 2692 4589 2748
rect 4589 2692 4645 2748
rect 4645 2692 4649 2748
rect 4585 2688 4649 2692
rect 4665 2748 4729 2752
rect 4665 2692 4669 2748
rect 4669 2692 4725 2748
rect 4725 2692 4729 2748
rect 4665 2688 4729 2692
rect 11371 2748 11435 2752
rect 11371 2692 11375 2748
rect 11375 2692 11431 2748
rect 11431 2692 11435 2748
rect 11371 2688 11435 2692
rect 11451 2748 11515 2752
rect 11451 2692 11455 2748
rect 11455 2692 11511 2748
rect 11511 2692 11515 2748
rect 11451 2688 11515 2692
rect 11531 2748 11595 2752
rect 11531 2692 11535 2748
rect 11535 2692 11591 2748
rect 11591 2692 11595 2748
rect 11531 2688 11595 2692
rect 11611 2748 11675 2752
rect 11611 2692 11615 2748
rect 11615 2692 11671 2748
rect 11671 2692 11675 2748
rect 11611 2688 11675 2692
rect 18317 2748 18381 2752
rect 18317 2692 18321 2748
rect 18321 2692 18377 2748
rect 18377 2692 18381 2748
rect 18317 2688 18381 2692
rect 18397 2748 18461 2752
rect 18397 2692 18401 2748
rect 18401 2692 18457 2748
rect 18457 2692 18461 2748
rect 18397 2688 18461 2692
rect 18477 2748 18541 2752
rect 18477 2692 18481 2748
rect 18481 2692 18537 2748
rect 18537 2692 18541 2748
rect 18477 2688 18541 2692
rect 18557 2748 18621 2752
rect 18557 2692 18561 2748
rect 18561 2692 18617 2748
rect 18617 2692 18621 2748
rect 18557 2688 18621 2692
rect 25263 2748 25327 2752
rect 25263 2692 25267 2748
rect 25267 2692 25323 2748
rect 25323 2692 25327 2748
rect 25263 2688 25327 2692
rect 25343 2748 25407 2752
rect 25343 2692 25347 2748
rect 25347 2692 25403 2748
rect 25403 2692 25407 2748
rect 25343 2688 25407 2692
rect 25423 2748 25487 2752
rect 25423 2692 25427 2748
rect 25427 2692 25483 2748
rect 25483 2692 25487 2748
rect 25423 2688 25487 2692
rect 25503 2748 25567 2752
rect 25503 2692 25507 2748
rect 25507 2692 25563 2748
rect 25563 2692 25567 2748
rect 25503 2688 25567 2692
rect 7898 2204 7962 2208
rect 7898 2148 7902 2204
rect 7902 2148 7958 2204
rect 7958 2148 7962 2204
rect 7898 2144 7962 2148
rect 7978 2204 8042 2208
rect 7978 2148 7982 2204
rect 7982 2148 8038 2204
rect 8038 2148 8042 2204
rect 7978 2144 8042 2148
rect 8058 2204 8122 2208
rect 8058 2148 8062 2204
rect 8062 2148 8118 2204
rect 8118 2148 8122 2204
rect 8058 2144 8122 2148
rect 8138 2204 8202 2208
rect 8138 2148 8142 2204
rect 8142 2148 8198 2204
rect 8198 2148 8202 2204
rect 8138 2144 8202 2148
rect 14844 2204 14908 2208
rect 14844 2148 14848 2204
rect 14848 2148 14904 2204
rect 14904 2148 14908 2204
rect 14844 2144 14908 2148
rect 14924 2204 14988 2208
rect 14924 2148 14928 2204
rect 14928 2148 14984 2204
rect 14984 2148 14988 2204
rect 14924 2144 14988 2148
rect 15004 2204 15068 2208
rect 15004 2148 15008 2204
rect 15008 2148 15064 2204
rect 15064 2148 15068 2204
rect 15004 2144 15068 2148
rect 15084 2204 15148 2208
rect 15084 2148 15088 2204
rect 15088 2148 15144 2204
rect 15144 2148 15148 2204
rect 15084 2144 15148 2148
rect 21790 2204 21854 2208
rect 21790 2148 21794 2204
rect 21794 2148 21850 2204
rect 21850 2148 21854 2204
rect 21790 2144 21854 2148
rect 21870 2204 21934 2208
rect 21870 2148 21874 2204
rect 21874 2148 21930 2204
rect 21930 2148 21934 2204
rect 21870 2144 21934 2148
rect 21950 2204 22014 2208
rect 21950 2148 21954 2204
rect 21954 2148 22010 2204
rect 22010 2148 22014 2204
rect 21950 2144 22014 2148
rect 22030 2204 22094 2208
rect 22030 2148 22034 2204
rect 22034 2148 22090 2204
rect 22090 2148 22094 2204
rect 22030 2144 22094 2148
rect 28736 2204 28800 2208
rect 28736 2148 28740 2204
rect 28740 2148 28796 2204
rect 28796 2148 28800 2204
rect 28736 2144 28800 2148
rect 28816 2204 28880 2208
rect 28816 2148 28820 2204
rect 28820 2148 28876 2204
rect 28876 2148 28880 2204
rect 28816 2144 28880 2148
rect 28896 2204 28960 2208
rect 28896 2148 28900 2204
rect 28900 2148 28956 2204
rect 28956 2148 28960 2204
rect 28896 2144 28960 2148
rect 28976 2204 29040 2208
rect 28976 2148 28980 2204
rect 28980 2148 29036 2204
rect 29036 2148 29040 2204
rect 28976 2144 29040 2148
<< metal4 >>
rect 4417 27776 4737 27792
rect 4417 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4737 27776
rect 4417 26688 4737 27712
rect 4417 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4737 26688
rect 4417 25600 4737 26624
rect 4417 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4737 25600
rect 4417 24512 4737 25536
rect 4417 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4737 24512
rect 4417 23424 4737 24448
rect 4417 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4737 23424
rect 4417 22336 4737 23360
rect 4417 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4737 22336
rect 4417 21248 4737 22272
rect 4417 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4737 21248
rect 4417 20160 4737 21184
rect 4417 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4737 20160
rect 4417 19072 4737 20096
rect 4417 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4737 19072
rect 4417 17984 4737 19008
rect 4417 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4737 17984
rect 4417 16896 4737 17920
rect 4417 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4737 16896
rect 4417 15808 4737 16832
rect 4417 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4737 15808
rect 4417 14720 4737 15744
rect 4417 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4737 14720
rect 4417 13632 4737 14656
rect 4417 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4737 13632
rect 4417 12544 4737 13568
rect 4417 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4737 12544
rect 4417 11456 4737 12480
rect 4417 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4737 11456
rect 4417 10368 4737 11392
rect 4417 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4737 10368
rect 4417 9280 4737 10304
rect 4417 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4737 9280
rect 4417 8192 4737 9216
rect 4417 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4737 8192
rect 4417 7104 4737 8128
rect 4417 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4737 7104
rect 4417 6016 4737 7040
rect 4417 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4737 6016
rect 4417 4928 4737 5952
rect 4417 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4737 4928
rect 4417 3840 4737 4864
rect 4417 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4737 3840
rect 4417 2752 4737 3776
rect 4417 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4737 2752
rect 4417 2128 4737 2688
rect 7890 27232 8210 27792
rect 7890 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8210 27232
rect 7890 26144 8210 27168
rect 7890 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8210 26144
rect 7890 25056 8210 26080
rect 7890 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8210 25056
rect 7890 23968 8210 24992
rect 7890 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8210 23968
rect 7890 22880 8210 23904
rect 7890 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8210 22880
rect 7890 21792 8210 22816
rect 7890 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8210 21792
rect 7890 20704 8210 21728
rect 7890 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8210 20704
rect 7890 19616 8210 20640
rect 7890 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8210 19616
rect 7890 18528 8210 19552
rect 7890 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8210 18528
rect 7890 17440 8210 18464
rect 7890 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8210 17440
rect 7890 16352 8210 17376
rect 7890 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8210 16352
rect 7890 15264 8210 16288
rect 7890 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8210 15264
rect 7890 14176 8210 15200
rect 7890 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8210 14176
rect 7890 13088 8210 14112
rect 7890 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8210 13088
rect 7890 12000 8210 13024
rect 7890 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8210 12000
rect 7890 10912 8210 11936
rect 7890 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8210 10912
rect 7890 9824 8210 10848
rect 7890 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8210 9824
rect 7890 8736 8210 9760
rect 7890 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8210 8736
rect 7890 7648 8210 8672
rect 7890 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8210 7648
rect 7890 6560 8210 7584
rect 7890 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8210 6560
rect 7890 5472 8210 6496
rect 7890 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8210 5472
rect 7890 4384 8210 5408
rect 7890 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8210 4384
rect 7890 3296 8210 4320
rect 7890 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8210 3296
rect 7890 2208 8210 3232
rect 7890 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8210 2208
rect 7890 2128 8210 2144
rect 11363 27776 11683 27792
rect 11363 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11683 27776
rect 11363 26688 11683 27712
rect 11363 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11683 26688
rect 11363 25600 11683 26624
rect 11363 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11683 25600
rect 11363 24512 11683 25536
rect 11363 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11683 24512
rect 11363 23424 11683 24448
rect 11363 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11683 23424
rect 11363 22336 11683 23360
rect 11363 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11683 22336
rect 11363 21248 11683 22272
rect 11363 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11683 21248
rect 11363 20160 11683 21184
rect 11363 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11683 20160
rect 11363 19072 11683 20096
rect 11363 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11683 19072
rect 11363 17984 11683 19008
rect 11363 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11683 17984
rect 11363 16896 11683 17920
rect 11363 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11683 16896
rect 11363 15808 11683 16832
rect 11363 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11683 15808
rect 11363 14720 11683 15744
rect 11363 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11683 14720
rect 11363 13632 11683 14656
rect 11363 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11683 13632
rect 11363 12544 11683 13568
rect 11363 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11683 12544
rect 11363 11456 11683 12480
rect 11363 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11683 11456
rect 11363 10368 11683 11392
rect 11363 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11683 10368
rect 11363 9280 11683 10304
rect 11363 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11683 9280
rect 11363 8192 11683 9216
rect 11363 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11683 8192
rect 11363 7104 11683 8128
rect 11363 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11683 7104
rect 11363 6016 11683 7040
rect 11363 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11683 6016
rect 11363 4928 11683 5952
rect 11363 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11683 4928
rect 11363 3840 11683 4864
rect 11363 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11683 3840
rect 11363 2752 11683 3776
rect 11363 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11683 2752
rect 11363 2128 11683 2688
rect 14836 27232 15156 27792
rect 14836 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15156 27232
rect 14836 26144 15156 27168
rect 14836 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15156 26144
rect 14836 25056 15156 26080
rect 14836 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15156 25056
rect 14836 23968 15156 24992
rect 14836 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15156 23968
rect 14836 22880 15156 23904
rect 14836 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15156 22880
rect 14836 21792 15156 22816
rect 14836 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15156 21792
rect 14836 20704 15156 21728
rect 14836 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15156 20704
rect 14836 19616 15156 20640
rect 14836 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15156 19616
rect 14836 18528 15156 19552
rect 14836 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15156 18528
rect 14836 17440 15156 18464
rect 14836 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15156 17440
rect 14836 16352 15156 17376
rect 14836 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15156 16352
rect 14836 15264 15156 16288
rect 14836 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15156 15264
rect 14836 14176 15156 15200
rect 14836 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15156 14176
rect 14836 13088 15156 14112
rect 14836 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15156 13088
rect 14836 12000 15156 13024
rect 14836 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15156 12000
rect 14836 10912 15156 11936
rect 14836 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15156 10912
rect 14836 9824 15156 10848
rect 14836 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15156 9824
rect 14836 8736 15156 9760
rect 14836 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15156 8736
rect 14836 7648 15156 8672
rect 14836 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15156 7648
rect 14836 6560 15156 7584
rect 14836 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15156 6560
rect 14836 5472 15156 6496
rect 14836 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15156 5472
rect 14836 4384 15156 5408
rect 14836 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15156 4384
rect 14836 3296 15156 4320
rect 14836 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15156 3296
rect 14836 2208 15156 3232
rect 14836 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15156 2208
rect 14836 2128 15156 2144
rect 18309 27776 18629 27792
rect 18309 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18629 27776
rect 18309 26688 18629 27712
rect 18309 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18629 26688
rect 18309 25600 18629 26624
rect 18309 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18629 25600
rect 18309 24512 18629 25536
rect 18309 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18629 24512
rect 18309 23424 18629 24448
rect 18309 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18629 23424
rect 18309 22336 18629 23360
rect 18309 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18629 22336
rect 18309 21248 18629 22272
rect 18309 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18629 21248
rect 18309 20160 18629 21184
rect 18309 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18629 20160
rect 18309 19072 18629 20096
rect 18309 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18629 19072
rect 18309 17984 18629 19008
rect 18309 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18629 17984
rect 18309 16896 18629 17920
rect 18309 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18629 16896
rect 18309 15808 18629 16832
rect 18309 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18629 15808
rect 18309 14720 18629 15744
rect 18309 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18629 14720
rect 18309 13632 18629 14656
rect 18309 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18629 13632
rect 18309 12544 18629 13568
rect 18309 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18629 12544
rect 18309 11456 18629 12480
rect 18309 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18629 11456
rect 18309 10368 18629 11392
rect 18309 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18629 10368
rect 18309 9280 18629 10304
rect 18309 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18629 9280
rect 18309 8192 18629 9216
rect 18309 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18629 8192
rect 18309 7104 18629 8128
rect 18309 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18629 7104
rect 18309 6016 18629 7040
rect 18309 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18629 6016
rect 18309 4928 18629 5952
rect 18309 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18629 4928
rect 18309 3840 18629 4864
rect 18309 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18629 3840
rect 18309 2752 18629 3776
rect 18309 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18629 2752
rect 18309 2128 18629 2688
rect 21782 27232 22102 27792
rect 21782 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22102 27232
rect 21782 26144 22102 27168
rect 21782 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22102 26144
rect 21782 25056 22102 26080
rect 21782 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22102 25056
rect 21782 23968 22102 24992
rect 21782 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22102 23968
rect 21782 22880 22102 23904
rect 21782 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22102 22880
rect 21782 21792 22102 22816
rect 21782 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22102 21792
rect 21782 20704 22102 21728
rect 21782 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22102 20704
rect 21782 19616 22102 20640
rect 21782 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22102 19616
rect 21782 18528 22102 19552
rect 21782 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22102 18528
rect 21782 17440 22102 18464
rect 21782 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22102 17440
rect 21782 16352 22102 17376
rect 21782 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22102 16352
rect 21782 15264 22102 16288
rect 21782 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22102 15264
rect 21782 14176 22102 15200
rect 21782 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22102 14176
rect 21782 13088 22102 14112
rect 21782 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22102 13088
rect 21782 12000 22102 13024
rect 21782 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22102 12000
rect 21782 10912 22102 11936
rect 21782 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22102 10912
rect 21782 9824 22102 10848
rect 21782 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22102 9824
rect 21782 8736 22102 9760
rect 21782 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22102 8736
rect 21782 7648 22102 8672
rect 21782 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22102 7648
rect 21782 6560 22102 7584
rect 21782 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22102 6560
rect 21782 5472 22102 6496
rect 21782 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22102 5472
rect 21782 4384 22102 5408
rect 21782 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22102 4384
rect 21782 3296 22102 4320
rect 21782 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22102 3296
rect 21782 2208 22102 3232
rect 21782 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22102 2208
rect 21782 2128 22102 2144
rect 25255 27776 25575 27792
rect 25255 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25575 27776
rect 25255 26688 25575 27712
rect 25255 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25575 26688
rect 25255 25600 25575 26624
rect 25255 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25575 25600
rect 25255 24512 25575 25536
rect 25255 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25575 24512
rect 25255 23424 25575 24448
rect 25255 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25575 23424
rect 25255 22336 25575 23360
rect 25255 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25575 22336
rect 25255 21248 25575 22272
rect 25255 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25575 21248
rect 25255 20160 25575 21184
rect 25255 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25575 20160
rect 25255 19072 25575 20096
rect 25255 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25575 19072
rect 25255 17984 25575 19008
rect 25255 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25575 17984
rect 25255 16896 25575 17920
rect 25255 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25575 16896
rect 25255 15808 25575 16832
rect 25255 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25575 15808
rect 25255 14720 25575 15744
rect 25255 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25575 14720
rect 25255 13632 25575 14656
rect 25255 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25575 13632
rect 25255 12544 25575 13568
rect 25255 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25575 12544
rect 25255 11456 25575 12480
rect 25255 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25575 11456
rect 25255 10368 25575 11392
rect 25255 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25575 10368
rect 25255 9280 25575 10304
rect 25255 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25575 9280
rect 25255 8192 25575 9216
rect 25255 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25575 8192
rect 25255 7104 25575 8128
rect 25255 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25575 7104
rect 25255 6016 25575 7040
rect 25255 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25575 6016
rect 25255 4928 25575 5952
rect 25255 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25575 4928
rect 25255 3840 25575 4864
rect 25255 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25575 3840
rect 25255 2752 25575 3776
rect 25255 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25575 2752
rect 25255 2128 25575 2688
rect 28728 27232 29048 27792
rect 28728 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29048 27232
rect 28728 26144 29048 27168
rect 28728 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29048 26144
rect 28728 25056 29048 26080
rect 28728 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29048 25056
rect 28728 23968 29048 24992
rect 28728 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29048 23968
rect 28728 22880 29048 23904
rect 28728 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29048 22880
rect 28728 21792 29048 22816
rect 28728 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29048 21792
rect 28728 20704 29048 21728
rect 28728 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29048 20704
rect 28728 19616 29048 20640
rect 28728 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29048 19616
rect 28728 18528 29048 19552
rect 28728 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29048 18528
rect 28728 17440 29048 18464
rect 28728 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29048 17440
rect 28728 16352 29048 17376
rect 28728 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29048 16352
rect 28728 15264 29048 16288
rect 28728 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29048 15264
rect 28728 14176 29048 15200
rect 28728 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29048 14176
rect 28728 13088 29048 14112
rect 28728 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29048 13088
rect 28728 12000 29048 13024
rect 28728 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29048 12000
rect 28728 10912 29048 11936
rect 28728 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29048 10912
rect 28728 9824 29048 10848
rect 28728 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29048 9824
rect 28728 8736 29048 9760
rect 28728 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29048 8736
rect 28728 7648 29048 8672
rect 28728 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29048 7648
rect 28728 6560 29048 7584
rect 28728 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29048 6560
rect 28728 5472 29048 6496
rect 28728 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29048 5472
rect 28728 4384 29048 5408
rect 28728 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29048 4384
rect 28728 3296 29048 4320
rect 28728 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29048 3296
rect 28728 2208 29048 3232
rect 28728 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29048 2208
rect 28728 2128 29048 2144
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121
timestamp 1676037725
transform 1 0 12236 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1676037725
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1676037725
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1676037725
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1676037725
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_289
timestamp 1676037725
transform 1 0 27692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_297
timestamp 1676037725
transform 1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_33
timestamp 1676037725
transform 1 0 4140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_80
timestamp 1676037725
transform 1 0 8464 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_92
timestamp 1676037725
transform 1 0 9568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_141
timestamp 1676037725
transform 1 0 14076 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_177
timestamp 1676037725
transform 1 0 17388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1676037725
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_206
timestamp 1676037725
transform 1 0 20056 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1676037725
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1676037725
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_268
timestamp 1676037725
transform 1 0 25760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_275
timestamp 1676037725
transform 1 0 26404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_286
timestamp 1676037725
transform 1 0 27416 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_298
timestamp 1676037725
transform 1 0 28520 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_44
timestamp 1676037725
transform 1 0 5152 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_52
timestamp 1676037725
transform 1 0 5888 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1676037725
transform 1 0 6348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_100
timestamp 1676037725
transform 1 0 10304 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_125
timestamp 1676037725
transform 1 0 12604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1676037725
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_147
timestamp 1676037725
transform 1 0 14628 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_164
timestamp 1676037725
transform 1 0 16192 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_184
timestamp 1676037725
transform 1 0 18032 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_206
timestamp 1676037725
transform 1 0 20056 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_214
timestamp 1676037725
transform 1 0 20792 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_237
timestamp 1676037725
transform 1 0 22908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp 1676037725
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_258
timestamp 1676037725
transform 1 0 24840 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_266
timestamp 1676037725
transform 1 0 25576 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_285
timestamp 1676037725
transform 1 0 27324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_292
timestamp 1676037725
transform 1 0 27968 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1676037725
transform 1 0 28520 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_21
timestamp 1676037725
transform 1 0 3036 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_25
timestamp 1676037725
transform 1 0 3404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50
timestamp 1676037725
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_63
timestamp 1676037725
transform 1 0 6900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_80
timestamp 1676037725
transform 1 0 8464 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_88
timestamp 1676037725
transform 1 0 9200 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_118
timestamp 1676037725
transform 1 0 11960 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_126
timestamp 1676037725
transform 1 0 12696 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_178
timestamp 1676037725
transform 1 0 17480 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_190
timestamp 1676037725
transform 1 0 18584 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_207
timestamp 1676037725
transform 1 0 20148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1676037725
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_256
timestamp 1676037725
transform 1 0 24656 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_274
timestamp 1676037725
transform 1 0 26312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_290
timestamp 1676037725
transform 1 0 27784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_297
timestamp 1676037725
transform 1 0 28428 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_40
timestamp 1676037725
transform 1 0 4784 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_52
timestamp 1676037725
transform 1 0 5888 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_69
timestamp 1676037725
transform 1 0 7452 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_76
timestamp 1676037725
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1676037725
transform 1 0 9660 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_114
timestamp 1676037725
transform 1 0 11592 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_126
timestamp 1676037725
transform 1 0 12696 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1676037725
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_230
timestamp 1676037725
transform 1 0 22264 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_273
timestamp 1676037725
transform 1 0 26220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_286
timestamp 1676037725
transform 1 0 27416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1676037725
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_36
timestamp 1676037725
transform 1 0 4416 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_48
timestamp 1676037725
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_64
timestamp 1676037725
transform 1 0 6992 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_73
timestamp 1676037725
transform 1 0 7820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_85
timestamp 1676037725
transform 1 0 8924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_97
timestamp 1676037725
transform 1 0 10028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp 1676037725
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_160
timestamp 1676037725
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_174
timestamp 1676037725
transform 1 0 17112 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_186
timestamp 1676037725
transform 1 0 18216 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_198
timestamp 1676037725
transform 1 0 19320 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_210
timestamp 1676037725
transform 1 0 20424 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_230
timestamp 1676037725
transform 1 0 22264 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_269
timestamp 1676037725
transform 1 0 25852 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_275
timestamp 1676037725
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_286
timestamp 1676037725
transform 1 0 27416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1676037725
transform 1 0 2116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1676037725
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_34
timestamp 1676037725
transform 1 0 4232 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_46
timestamp 1676037725
transform 1 0 5336 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_63
timestamp 1676037725
transform 1 0 6900 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_74
timestamp 1676037725
transform 1 0 7912 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1676037725
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1676037725
transform 1 0 9660 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_104
timestamp 1676037725
transform 1 0 10672 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_123
timestamp 1676037725
transform 1 0 12420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1676037725
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_147
timestamp 1676037725
transform 1 0 14628 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_151
timestamp 1676037725
transform 1 0 14996 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_176
timestamp 1676037725
transform 1 0 17296 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_188
timestamp 1676037725
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_220
timestamp 1676037725
transform 1 0 21344 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_227
timestamp 1676037725
transform 1 0 21988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_239
timestamp 1676037725
transform 1 0 23092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_273
timestamp 1676037725
transform 1 0 26220 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_291
timestamp 1676037725
transform 1 0 27876 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_18
timestamp 1676037725
transform 1 0 2760 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_25
timestamp 1676037725
transform 1 0 3404 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_37
timestamp 1676037725
transform 1 0 4508 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1676037725
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_65
timestamp 1676037725
transform 1 0 7084 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_76
timestamp 1676037725
transform 1 0 8096 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_88
timestamp 1676037725
transform 1 0 9200 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1676037725
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_133
timestamp 1676037725
transform 1 0 13340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_145
timestamp 1676037725
transform 1 0 14444 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_157
timestamp 1676037725
transform 1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1676037725
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_177
timestamp 1676037725
transform 1 0 17388 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_206
timestamp 1676037725
transform 1 0 20056 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_213
timestamp 1676037725
transform 1 0 20700 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp 1676037725
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_253
timestamp 1676037725
transform 1 0 24380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_265
timestamp 1676037725
transform 1 0 25484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1676037725
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_289
timestamp 1676037725
transform 1 0 27692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_297
timestamp 1676037725
transform 1 0 28428 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1676037725
transform 1 0 2116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1676037725
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_50
timestamp 1676037725
transform 1 0 5704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_63
timestamp 1676037725
transform 1 0 6900 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_78
timestamp 1676037725
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_107
timestamp 1676037725
transform 1 0 10948 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_119
timestamp 1676037725
transform 1 0 12052 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp 1676037725
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_191
timestamp 1676037725
transform 1 0 18676 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_202
timestamp 1676037725
transform 1 0 19688 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_214
timestamp 1676037725
transform 1 0 20792 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_226
timestamp 1676037725
transform 1 0 21896 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_270
timestamp 1676037725
transform 1 0 25944 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_290
timestamp 1676037725
transform 1 0 27784 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1676037725
transform 1 0 28520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_32
timestamp 1676037725
transform 1 0 4048 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1676037725
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_65
timestamp 1676037725
transform 1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_77
timestamp 1676037725
transform 1 0 8188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_89
timestamp 1676037725
transform 1 0 9292 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_95
timestamp 1676037725
transform 1 0 9844 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_152
timestamp 1676037725
transform 1 0 15088 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1676037725
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_185
timestamp 1676037725
transform 1 0 18124 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_206
timestamp 1676037725
transform 1 0 20056 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_214
timestamp 1676037725
transform 1 0 20792 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1676037725
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_267
timestamp 1676037725
transform 1 0 25668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1676037725
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_288
timestamp 1676037725
transform 1 0 27600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_295
timestamp 1676037725
transform 1 0 28244 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_18
timestamp 1676037725
transform 1 0 2760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1676037725
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_57
timestamp 1676037725
transform 1 0 6348 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp 1676037725
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_93
timestamp 1676037725
transform 1 0 9660 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_164
timestamp 1676037725
transform 1 0 16192 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_181
timestamp 1676037725
transform 1 0 17756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1676037725
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_205
timestamp 1676037725
transform 1 0 19964 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_225
timestamp 1676037725
transform 1 0 21804 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1676037725
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_258
timestamp 1676037725
transform 1 0 24840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_270
timestamp 1676037725
transform 1 0 25944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_280
timestamp 1676037725
transform 1 0 26864 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_291
timestamp 1676037725
transform 1 0 27876 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1676037725
transform 1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_34
timestamp 1676037725
transform 1 0 4232 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_46
timestamp 1676037725
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1676037725
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_77
timestamp 1676037725
transform 1 0 8188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_89
timestamp 1676037725
transform 1 0 9292 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_101
timestamp 1676037725
transform 1 0 10396 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1676037725
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_118
timestamp 1676037725
transform 1 0 11960 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_130
timestamp 1676037725
transform 1 0 13064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_162
timestamp 1676037725
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_192
timestamp 1676037725
transform 1 0 18768 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_204
timestamp 1676037725
transform 1 0 19872 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_216
timestamp 1676037725
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_233
timestamp 1676037725
transform 1 0 22540 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_257
timestamp 1676037725
transform 1 0 24748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1676037725
transform 1 0 25852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp 1676037725
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_290
timestamp 1676037725
transform 1 0 27784 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_298
timestamp 1676037725
transform 1 0 28520 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1676037725
transform 1 0 2116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1676037725
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_68
timestamp 1676037725
transform 1 0 7360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1676037725
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_94
timestamp 1676037725
transform 1 0 9752 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_103
timestamp 1676037725
transform 1 0 10580 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_107
timestamp 1676037725
transform 1 0 10948 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_117
timestamp 1676037725
transform 1 0 11868 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_129
timestamp 1676037725
transform 1 0 12972 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1676037725
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_156
timestamp 1676037725
transform 1 0 15456 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_160
timestamp 1676037725
transform 1 0 15824 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_164
timestamp 1676037725
transform 1 0 16192 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_170
timestamp 1676037725
transform 1 0 16744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_187
timestamp 1676037725
transform 1 0 18308 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_212
timestamp 1676037725
transform 1 0 20608 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_224
timestamp 1676037725
transform 1 0 21712 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_232
timestamp 1676037725
transform 1 0 22448 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_237
timestamp 1676037725
transform 1 0 22908 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_287
timestamp 1676037725
transform 1 0 27508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_297
timestamp 1676037725
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_19
timestamp 1676037725
transform 1 0 2852 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_31
timestamp 1676037725
transform 1 0 3956 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_40
timestamp 1676037725
transform 1 0 4784 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1676037725
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_89
timestamp 1676037725
transform 1 0 9292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_95
timestamp 1676037725
transform 1 0 9844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1676037725
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_145
timestamp 1676037725
transform 1 0 14444 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_151
timestamp 1676037725
transform 1 0 14996 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp 1676037725
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_175
timestamp 1676037725
transform 1 0 17204 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_179
timestamp 1676037725
transform 1 0 17572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_191
timestamp 1676037725
transform 1 0 18676 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1676037725
transform 1 0 20884 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1676037725
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_273
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1676037725
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_289
timestamp 1676037725
transform 1 0 27692 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_297
timestamp 1676037725
transform 1 0 28428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_11
timestamp 1676037725
transform 1 0 2116 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_44
timestamp 1676037725
transform 1 0 5152 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_50
timestamp 1676037725
transform 1 0 5704 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_58
timestamp 1676037725
transform 1 0 6440 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1676037725
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_93
timestamp 1676037725
transform 1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_112
timestamp 1676037725
transform 1 0 11408 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_125
timestamp 1676037725
transform 1 0 12604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1676037725
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_183
timestamp 1676037725
transform 1 0 17940 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_204
timestamp 1676037725
transform 1 0 19872 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_229
timestamp 1676037725
transform 1 0 22172 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1676037725
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_277
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_281
timestamp 1676037725
transform 1 0 26956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_289
timestamp 1676037725
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp 1676037725
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_11
timestamp 1676037725
transform 1 0 2116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_16
timestamp 1676037725
transform 1 0 2576 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_23
timestamp 1676037725
transform 1 0 3220 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_48
timestamp 1676037725
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_88
timestamp 1676037725
transform 1 0 9200 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_100
timestamp 1676037725
transform 1 0 10304 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_131
timestamp 1676037725
transform 1 0 13156 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_148
timestamp 1676037725
transform 1 0 14720 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_160
timestamp 1676037725
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_180
timestamp 1676037725
transform 1 0 17664 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_192
timestamp 1676037725
transform 1 0 18768 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1676037725
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_233
timestamp 1676037725
transform 1 0 22540 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_257
timestamp 1676037725
transform 1 0 24748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1676037725
transform 1 0 25852 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1676037725
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_289
timestamp 1676037725
transform 1 0 27692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_297
timestamp 1676037725
transform 1 0 28428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1676037725
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_49
timestamp 1676037725
transform 1 0 5612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_64
timestamp 1676037725
transform 1 0 6992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_71
timestamp 1676037725
transform 1 0 7636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_75
timestamp 1676037725
transform 1 0 8004 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1676037725
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_94
timestamp 1676037725
transform 1 0 9752 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_102
timestamp 1676037725
transform 1 0 10488 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_107
timestamp 1676037725
transform 1 0 10948 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_117
timestamp 1676037725
transform 1 0 11868 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_129
timestamp 1676037725
transform 1 0 12972 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1676037725
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_152
timestamp 1676037725
transform 1 0 15088 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_164
timestamp 1676037725
transform 1 0 16192 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_175
timestamp 1676037725
transform 1 0 17204 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_187
timestamp 1676037725
transform 1 0 18308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1676037725
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_205
timestamp 1676037725
transform 1 0 19964 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_213
timestamp 1676037725
transform 1 0 20700 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_237
timestamp 1676037725
transform 1 0 22908 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 1676037725
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_259
timestamp 1676037725
transform 1 0 24932 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_265
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_279
timestamp 1676037725
transform 1 0 26772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_291
timestamp 1676037725
transform 1 0 27876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_11
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_25
timestamp 1676037725
transform 1 0 3404 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1676037725
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_68
timestamp 1676037725
transform 1 0 7360 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_80
timestamp 1676037725
transform 1 0 8464 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_92
timestamp 1676037725
transform 1 0 9568 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_100
timestamp 1676037725
transform 1 0 10304 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1676037725
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_138
timestamp 1676037725
transform 1 0 13800 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_146
timestamp 1676037725
transform 1 0 14536 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_156
timestamp 1676037725
transform 1 0 15456 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_187
timestamp 1676037725
transform 1 0 18308 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_195
timestamp 1676037725
transform 1 0 19044 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_205
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_233
timestamp 1676037725
transform 1 0 22540 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_243
timestamp 1676037725
transform 1 0 23460 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_250
timestamp 1676037725
transform 1 0 24104 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_256
timestamp 1676037725
transform 1 0 24656 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1676037725
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_296
timestamp 1676037725
transform 1 0 28336 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_40
timestamp 1676037725
transform 1 0 4784 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_48
timestamp 1676037725
transform 1 0 5520 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_66
timestamp 1676037725
transform 1 0 7176 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_78
timestamp 1676037725
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_96
timestamp 1676037725
transform 1 0 9936 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_104
timestamp 1676037725
transform 1 0 10672 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_111
timestamp 1676037725
transform 1 0 11316 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_117
timestamp 1676037725
transform 1 0 11868 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_128
timestamp 1676037725
transform 1 0 12880 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_152
timestamp 1676037725
transform 1 0 15088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_159
timestamp 1676037725
transform 1 0 15732 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1676037725
transform 1 0 16468 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_176
timestamp 1676037725
transform 1 0 17296 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_188
timestamp 1676037725
transform 1 0 18400 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_208
timestamp 1676037725
transform 1 0 20240 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_219
timestamp 1676037725
transform 1 0 21252 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_231
timestamp 1676037725
transform 1 0 22356 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_243
timestamp 1676037725
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_268
timestamp 1676037725
transform 1 0 25760 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_274
timestamp 1676037725
transform 1 0 26312 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_296
timestamp 1676037725
transform 1 0 28336 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_28
timestamp 1676037725
transform 1 0 3680 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_48
timestamp 1676037725
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_68
timestamp 1676037725
transform 1 0 7360 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_96
timestamp 1676037725
transform 1 0 9936 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1676037725
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp 1676037725
transform 1 0 15824 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_180
timestamp 1676037725
transform 1 0 17664 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_192
timestamp 1676037725
transform 1 0 18768 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_209
timestamp 1676037725
transform 1 0 20332 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_215
timestamp 1676037725
transform 1 0 20884 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_229
timestamp 1676037725
transform 1 0 22172 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_246
timestamp 1676037725
transform 1 0 23736 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_258
timestamp 1676037725
transform 1 0 24840 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_270
timestamp 1676037725
transform 1 0 25944 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1676037725
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_286
timestamp 1676037725
transform 1 0 27416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_290
timestamp 1676037725
transform 1 0 27784 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_297
timestamp 1676037725
transform 1 0 28428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_8
timestamp 1676037725
transform 1 0 1840 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_22
timestamp 1676037725
transform 1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_55
timestamp 1676037725
transform 1 0 6164 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_75
timestamp 1676037725
transform 1 0 8004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1676037725
transform 1 0 9660 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_108
timestamp 1676037725
transform 1 0 11040 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_114
timestamp 1676037725
transform 1 0 11592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_130
timestamp 1676037725
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1676037725
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_151
timestamp 1676037725
transform 1 0 14996 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_175
timestamp 1676037725
transform 1 0 17204 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_187
timestamp 1676037725
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_207
timestamp 1676037725
transform 1 0 20148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_219
timestamp 1676037725
transform 1 0 21252 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_227
timestamp 1676037725
transform 1 0 21988 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_235
timestamp 1676037725
transform 1 0 22724 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1676037725
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_262
timestamp 1676037725
transform 1 0 25208 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_270
timestamp 1676037725
transform 1 0 25944 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_294
timestamp 1676037725
transform 1 0 28152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_298
timestamp 1676037725
transform 1 0 28520 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_9
timestamp 1676037725
transform 1 0 1932 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_33
timestamp 1676037725
transform 1 0 4140 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_43
timestamp 1676037725
transform 1 0 5060 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_50
timestamp 1676037725
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_62
timestamp 1676037725
transform 1 0 6808 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_95
timestamp 1676037725
transform 1 0 9844 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 1676037725
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_129
timestamp 1676037725
transform 1 0 12972 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_155
timestamp 1676037725
transform 1 0 15364 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1676037725
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_175
timestamp 1676037725
transform 1 0 17204 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_188
timestamp 1676037725
transform 1 0 18400 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_200
timestamp 1676037725
transform 1 0 19504 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_208
timestamp 1676037725
transform 1 0 20240 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_233
timestamp 1676037725
transform 1 0 22540 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_252
timestamp 1676037725
transform 1 0 24288 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_272
timestamp 1676037725
transform 1 0 26128 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1676037725
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_296
timestamp 1676037725
transform 1 0 28336 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_12
timestamp 1676037725
transform 1 0 2208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_19
timestamp 1676037725
transform 1 0 2852 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1676037725
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_45
timestamp 1676037725
transform 1 0 5244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_72
timestamp 1676037725
transform 1 0 7728 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1676037725
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_118
timestamp 1676037725
transform 1 0 11960 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_125
timestamp 1676037725
transform 1 0 12604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_152
timestamp 1676037725
transform 1 0 15088 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_161
timestamp 1676037725
transform 1 0 15916 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_173
timestamp 1676037725
transform 1 0 17020 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_185
timestamp 1676037725
transform 1 0 18124 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1676037725
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_232
timestamp 1676037725
transform 1 0 22448 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_244
timestamp 1676037725
transform 1 0 23552 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_288
timestamp 1676037725
transform 1 0 27600 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_296
timestamp 1676037725
transform 1 0 28336 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_32
timestamp 1676037725
transform 1 0 4048 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp 1676037725
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1676037725
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_62
timestamp 1676037725
transform 1 0 6808 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_68
timestamp 1676037725
transform 1 0 7360 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_72
timestamp 1676037725
transform 1 0 7728 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_84
timestamp 1676037725
transform 1 0 8832 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_92
timestamp 1676037725
transform 1 0 9568 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_144
timestamp 1676037725
transform 1 0 14352 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_159
timestamp 1676037725
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_191
timestamp 1676037725
transform 1 0 18676 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_202
timestamp 1676037725
transform 1 0 19688 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_210
timestamp 1676037725
transform 1 0 20424 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_214
timestamp 1676037725
transform 1 0 20792 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1676037725
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1676037725
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_249
timestamp 1676037725
transform 1 0 24012 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_257
timestamp 1676037725
transform 1 0 24748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_261
timestamp 1676037725
transform 1 0 25116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1676037725
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_286
timestamp 1676037725
transform 1 0 27416 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_298
timestamp 1676037725
transform 1 0 28520 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_10
timestamp 1676037725
transform 1 0 2024 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_17
timestamp 1676037725
transform 1 0 2668 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_21
timestamp 1676037725
transform 1 0 3036 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1676037725
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_47
timestamp 1676037725
transform 1 0 5428 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_69
timestamp 1676037725
transform 1 0 7452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1676037725
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_99
timestamp 1676037725
transform 1 0 10212 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_114
timestamp 1676037725
transform 1 0 11592 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_122
timestamp 1676037725
transform 1 0 12328 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_132
timestamp 1676037725
transform 1 0 13248 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_163
timestamp 1676037725
transform 1 0 16100 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_183
timestamp 1676037725
transform 1 0 17940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_205
timestamp 1676037725
transform 1 0 19964 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_213
timestamp 1676037725
transform 1 0 20700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_225
timestamp 1676037725
transform 1 0 21804 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_233
timestamp 1676037725
transform 1 0 22540 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_238
timestamp 1676037725
transform 1 0 23000 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_269
timestamp 1676037725
transform 1 0 25852 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_273
timestamp 1676037725
transform 1 0 26220 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_285
timestamp 1676037725
transform 1 0 27324 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1676037725
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1676037725
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1676037725
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1676037725
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1676037725
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_72
timestamp 1676037725
transform 1 0 7728 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_84
timestamp 1676037725
transform 1 0 8832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_96
timestamp 1676037725
transform 1 0 9936 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_102
timestamp 1676037725
transform 1 0 10488 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_124
timestamp 1676037725
transform 1 0 12512 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_128
timestamp 1676037725
transform 1 0 12880 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_177
timestamp 1676037725
transform 1 0 17388 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_194
timestamp 1676037725
transform 1 0 18952 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_214
timestamp 1676037725
transform 1 0 20792 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_234
timestamp 1676037725
transform 1 0 22632 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_247
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_259
timestamp 1676037725
transform 1 0 24932 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_271
timestamp 1676037725
transform 1 0 26036 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1676037725
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_293
timestamp 1676037725
transform 1 0 28060 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_11
timestamp 1676037725
transform 1 0 2116 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_16
timestamp 1676037725
transform 1 0 2576 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_26_25
timestamp 1676037725
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1676037725
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_103
timestamp 1676037725
transform 1 0 10580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_111
timestamp 1676037725
transform 1 0 11316 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_123
timestamp 1676037725
transform 1 0 12420 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_152
timestamp 1676037725
transform 1 0 15088 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_160
timestamp 1676037725
transform 1 0 15824 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_172
timestamp 1676037725
transform 1 0 16928 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_184
timestamp 1676037725
transform 1 0 18032 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_221
timestamp 1676037725
transform 1 0 21436 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_229
timestamp 1676037725
transform 1 0 22172 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_263
timestamp 1676037725
transform 1 0 25300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_275
timestamp 1676037725
transform 1 0 26404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_281
timestamp 1676037725
transform 1 0 26956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_289
timestamp 1676037725
transform 1 0 27692 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_297
timestamp 1676037725
transform 1 0 28428 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_19
timestamp 1676037725
transform 1 0 2852 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_31
timestamp 1676037725
transform 1 0 3956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_37
timestamp 1676037725
transform 1 0 4508 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1676037725
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_65
timestamp 1676037725
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1676037725
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_132
timestamp 1676037725
transform 1 0 13248 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_147
timestamp 1676037725
transform 1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_156
timestamp 1676037725
transform 1 0 15456 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_174
timestamp 1676037725
transform 1 0 17112 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_186
timestamp 1676037725
transform 1 0 18216 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_198
timestamp 1676037725
transform 1 0 19320 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_210
timestamp 1676037725
transform 1 0 20424 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_250
timestamp 1676037725
transform 1 0 24104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_264
timestamp 1676037725
transform 1 0 25392 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_275
timestamp 1676037725
transform 1 0 26404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1676037725
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_289
timestamp 1676037725
transform 1 0 27692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_297
timestamp 1676037725
transform 1 0 28428 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1676037725
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_34
timestamp 1676037725
transform 1 0 4232 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_49
timestamp 1676037725
transform 1 0 5612 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_69
timestamp 1676037725
transform 1 0 7452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1676037725
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_94
timestamp 1676037725
transform 1 0 9752 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_106
timestamp 1676037725
transform 1 0 10856 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_114
timestamp 1676037725
transform 1 0 11592 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1676037725
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_156
timestamp 1676037725
transform 1 0 15456 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_174
timestamp 1676037725
transform 1 0 17112 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_186
timestamp 1676037725
transform 1 0 18216 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_206
timestamp 1676037725
transform 1 0 20056 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_218
timestamp 1676037725
transform 1 0 21160 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_226
timestamp 1676037725
transform 1 0 21896 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_237
timestamp 1676037725
transform 1 0 22908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1676037725
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_271
timestamp 1676037725
transform 1 0 26036 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_283
timestamp 1676037725
transform 1 0 27140 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_297
timestamp 1676037725
transform 1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_36
timestamp 1676037725
transform 1 0 4416 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1676037725
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_62
timestamp 1676037725
transform 1 0 6808 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_70
timestamp 1676037725
transform 1 0 7544 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_144
timestamp 1676037725
transform 1 0 14352 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_151
timestamp 1676037725
transform 1 0 14996 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1676037725
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_178
timestamp 1676037725
transform 1 0 17480 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_190
timestamp 1676037725
transform 1 0 18584 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_212
timestamp 1676037725
transform 1 0 20608 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_249
timestamp 1676037725
transform 1 0 24012 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_260
timestamp 1676037725
transform 1 0 25024 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_264
timestamp 1676037725
transform 1 0 25392 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1676037725
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_36
timestamp 1676037725
transform 1 0 4416 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_48
timestamp 1676037725
transform 1 0 5520 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_62
timestamp 1676037725
transform 1 0 6808 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_74
timestamp 1676037725
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1676037725
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_103
timestamp 1676037725
transform 1 0 10580 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_115
timestamp 1676037725
transform 1 0 11684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_127
timestamp 1676037725
transform 1 0 12788 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_166
timestamp 1676037725
transform 1 0 16376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1676037725
transform 1 0 20884 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_228
timestamp 1676037725
transform 1 0 22080 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_236
timestamp 1676037725
transform 1 0 22816 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1676037725
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_262
timestamp 1676037725
transform 1 0 25208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_266
timestamp 1676037725
transform 1 0 25576 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_288
timestamp 1676037725
transform 1 0 27600 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_296
timestamp 1676037725
transform 1 0 28336 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_24
timestamp 1676037725
transform 1 0 3312 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_30
timestamp 1676037725
transform 1 0 3864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_37
timestamp 1676037725
transform 1 0 4508 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_45
timestamp 1676037725
transform 1 0 5244 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1676037725
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_62
timestamp 1676037725
transform 1 0 6808 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_82
timestamp 1676037725
transform 1 0 8648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_86
timestamp 1676037725
transform 1 0 9016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_96
timestamp 1676037725
transform 1 0 9936 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 1676037725
transform 1 0 10672 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_124
timestamp 1676037725
transform 1 0 12512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_133
timestamp 1676037725
transform 1 0 13340 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_144
timestamp 1676037725
transform 1 0 14352 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_156
timestamp 1676037725
transform 1 0 15456 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1676037725
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_176
timestamp 1676037725
transform 1 0 17296 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_188
timestamp 1676037725
transform 1 0 18400 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_200
timestamp 1676037725
transform 1 0 19504 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_218
timestamp 1676037725
transform 1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_230
timestamp 1676037725
transform 1 0 22264 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_250
timestamp 1676037725
transform 1 0 24104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_254
timestamp 1676037725
transform 1 0 24472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_262
timestamp 1676037725
transform 1 0 25208 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1676037725
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1676037725
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_296
timestamp 1676037725
transform 1 0 28336 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_9
timestamp 1676037725
transform 1 0 1932 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1676037725
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_57
timestamp 1676037725
transform 1 0 6348 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1676037725
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_94
timestamp 1676037725
transform 1 0 9752 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_118
timestamp 1676037725
transform 1 0 11960 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_126
timestamp 1676037725
transform 1 0 12696 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1676037725
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_156
timestamp 1676037725
transform 1 0 15456 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_164
timestamp 1676037725
transform 1 0 16192 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_175
timestamp 1676037725
transform 1 0 17204 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_184
timestamp 1676037725
transform 1 0 18032 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_201
timestamp 1676037725
transform 1 0 19596 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_208
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_214
timestamp 1676037725
transform 1 0 20792 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_220
timestamp 1676037725
transform 1 0 21344 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_232
timestamp 1676037725
transform 1 0 22448 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_264
timestamp 1676037725
transform 1 0 25392 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_268
timestamp 1676037725
transform 1 0 25760 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_272
timestamp 1676037725
transform 1 0 26128 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp 1676037725
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_9
timestamp 1676037725
transform 1 0 1932 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_26
timestamp 1676037725
transform 1 0 3496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_36
timestamp 1676037725
transform 1 0 4416 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_45
timestamp 1676037725
transform 1 0 5244 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_49
timestamp 1676037725
transform 1 0 5612 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1676037725
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_82
timestamp 1676037725
transform 1 0 8648 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_90
timestamp 1676037725
transform 1 0 9384 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_98
timestamp 1676037725
transform 1 0 10120 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1676037725
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_123
timestamp 1676037725
transform 1 0 12420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_133
timestamp 1676037725
transform 1 0 13340 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_153
timestamp 1676037725
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1676037725
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_187
timestamp 1676037725
transform 1 0 18308 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_199
timestamp 1676037725
transform 1 0 19412 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_207
timestamp 1676037725
transform 1 0 20148 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_219
timestamp 1676037725
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_232
timestamp 1676037725
transform 1 0 22448 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_240
timestamp 1676037725
transform 1 0 23184 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_262
timestamp 1676037725
transform 1 0 25208 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_274
timestamp 1676037725
transform 1 0 26312 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_286
timestamp 1676037725
transform 1 0 27416 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_298
timestamp 1676037725
transform 1 0 28520 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_25
timestamp 1676037725
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_45
timestamp 1676037725
transform 1 0 5244 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_67
timestamp 1676037725
transform 1 0 7268 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1676037725
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_121
timestamp 1676037725
transform 1 0 12236 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_152
timestamp 1676037725
transform 1 0 15088 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_164
timestamp 1676037725
transform 1 0 16192 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_185
timestamp 1676037725
transform 1 0 18124 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1676037725
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_221
timestamp 1676037725
transform 1 0 21436 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_233
timestamp 1676037725
transform 1 0 22540 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_241
timestamp 1676037725
transform 1 0 23276 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_263
timestamp 1676037725
transform 1 0 25300 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_275
timestamp 1676037725
transform 1 0 26404 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_287
timestamp 1676037725
transform 1 0 27508 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp 1676037725
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_14
timestamp 1676037725
transform 1 0 2392 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_24
timestamp 1676037725
transform 1 0 3312 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_34
timestamp 1676037725
transform 1 0 4232 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_46
timestamp 1676037725
transform 1 0 5336 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_62
timestamp 1676037725
transform 1 0 6808 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_74
timestamp 1676037725
transform 1 0 7912 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_86
timestamp 1676037725
transform 1 0 9016 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_103
timestamp 1676037725
transform 1 0 10580 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_121
timestamp 1676037725
transform 1 0 12236 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_138
timestamp 1676037725
transform 1 0 13800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_142
timestamp 1676037725
transform 1 0 14168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_150
timestamp 1676037725
transform 1 0 14904 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_157
timestamp 1676037725
transform 1 0 15548 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1676037725
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_188
timestamp 1676037725
transform 1 0 18400 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_194
timestamp 1676037725
transform 1 0 18952 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_202
timestamp 1676037725
transform 1 0 19688 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_214
timestamp 1676037725
transform 1 0 20792 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_230
timestamp 1676037725
transform 1 0 22264 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_238
timestamp 1676037725
transform 1 0 23000 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_249
timestamp 1676037725
transform 1 0 24012 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_260
timestamp 1676037725
transform 1 0 25024 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_272
timestamp 1676037725
transform 1 0 26128 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1676037725
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_296
timestamp 1676037725
transform 1 0 28336 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_9
timestamp 1676037725
transform 1 0 1932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1676037725
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_36
timestamp 1676037725
transform 1 0 4416 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_61
timestamp 1676037725
transform 1 0 6716 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_69
timestamp 1676037725
transform 1 0 7452 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1676037725
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_119
timestamp 1676037725
transform 1 0 12052 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_128
timestamp 1676037725
transform 1 0 12880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_156
timestamp 1676037725
transform 1 0 15456 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_168
timestamp 1676037725
transform 1 0 16560 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_174
timestamp 1676037725
transform 1 0 17112 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_191
timestamp 1676037725
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1676037725
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_206
timestamp 1676037725
transform 1 0 20056 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_218
timestamp 1676037725
transform 1 0 21160 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_230
timestamp 1676037725
transform 1 0 22264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_265
timestamp 1676037725
transform 1 0 25484 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_294
timestamp 1676037725
transform 1 0 28152 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_298
timestamp 1676037725
transform 1 0 28520 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_11
timestamp 1676037725
transform 1 0 2116 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_28
timestamp 1676037725
transform 1 0 3680 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_37
timestamp 1676037725
transform 1 0 4508 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_48
timestamp 1676037725
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_89
timestamp 1676037725
transform 1 0 9292 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_106
timestamp 1676037725
transform 1 0 10856 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_123
timestamp 1676037725
transform 1 0 12420 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_138
timestamp 1676037725
transform 1 0 13800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_165
timestamp 1676037725
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_177
timestamp 1676037725
transform 1 0 17388 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_187
timestamp 1676037725
transform 1 0 18308 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_212
timestamp 1676037725
transform 1 0 20608 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_233
timestamp 1676037725
transform 1 0 22540 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_254
timestamp 1676037725
transform 1 0 24472 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_266
timestamp 1676037725
transform 1 0 25576 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_274
timestamp 1676037725
transform 1 0 26312 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1676037725
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_286
timestamp 1676037725
transform 1 0 27416 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_298
timestamp 1676037725
transform 1 0 28520 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_11
timestamp 1676037725
transform 1 0 2116 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_16
timestamp 1676037725
transform 1 0 2576 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1676037725
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_51
timestamp 1676037725
transform 1 0 5796 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_68
timestamp 1676037725
transform 1 0 7360 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_72
timestamp 1676037725
transform 1 0 7728 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1676037725
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_97
timestamp 1676037725
transform 1 0 10028 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_110
timestamp 1676037725
transform 1 0 11224 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_118
timestamp 1676037725
transform 1 0 11960 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_124
timestamp 1676037725
transform 1 0 12512 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1676037725
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_152
timestamp 1676037725
transform 1 0 15088 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_159
timestamp 1676037725
transform 1 0 15732 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_171
timestamp 1676037725
transform 1 0 16836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_183
timestamp 1676037725
transform 1 0 17940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1676037725
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_213
timestamp 1676037725
transform 1 0 20700 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_234
timestamp 1676037725
transform 1 0 22632 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_242
timestamp 1676037725
transform 1 0 23368 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_262
timestamp 1676037725
transform 1 0 25208 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_274
timestamp 1676037725
transform 1 0 26312 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_296
timestamp 1676037725
transform 1 0 28336 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_36
timestamp 1676037725
transform 1 0 4416 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_48
timestamp 1676037725
transform 1 0 5520 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_80
timestamp 1676037725
transform 1 0 8464 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_92
timestamp 1676037725
transform 1 0 9568 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_104
timestamp 1676037725
transform 1 0 10672 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_137
timestamp 1676037725
transform 1 0 13708 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_154
timestamp 1676037725
transform 1 0 15272 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_189
timestamp 1676037725
transform 1 0 18492 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_213
timestamp 1676037725
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1676037725
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_243
timestamp 1676037725
transform 1 0 23460 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_255
timestamp 1676037725
transform 1 0 24564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_267
timestamp 1676037725
transform 1 0 25668 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_296
timestamp 1676037725
transform 1 0 28336 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_22
timestamp 1676037725
transform 1 0 3128 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_34
timestamp 1676037725
transform 1 0 4232 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_46
timestamp 1676037725
transform 1 0 5336 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_54
timestamp 1676037725
transform 1 0 6072 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_60
timestamp 1676037725
transform 1 0 6624 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_72
timestamp 1676037725
transform 1 0 7728 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_117
timestamp 1676037725
transform 1 0 11868 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_127
timestamp 1676037725
transform 1 0 12788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1676037725
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_159
timestamp 1676037725
transform 1 0 15732 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_171
timestamp 1676037725
transform 1 0 16836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_182
timestamp 1676037725
transform 1 0 17848 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_188
timestamp 1676037725
transform 1 0 18400 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1676037725
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_202
timestamp 1676037725
transform 1 0 19688 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_214
timestamp 1676037725
transform 1 0 20792 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_226
timestamp 1676037725
transform 1 0 21896 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_236
timestamp 1676037725
transform 1 0 22816 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1676037725
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1676037725
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1676037725
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_289
timestamp 1676037725
transform 1 0 27692 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_297
timestamp 1676037725
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_35
timestamp 1676037725
transform 1 0 4324 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_47
timestamp 1676037725
transform 1 0 5428 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_78
timestamp 1676037725
transform 1 0 8280 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_90
timestamp 1676037725
transform 1 0 9384 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_102
timestamp 1676037725
transform 1 0 10488 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1676037725
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_124
timestamp 1676037725
transform 1 0 12512 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_136
timestamp 1676037725
transform 1 0 13616 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_142
timestamp 1676037725
transform 1 0 14168 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_150
timestamp 1676037725
transform 1 0 14904 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_162
timestamp 1676037725
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_187
timestamp 1676037725
transform 1 0 18308 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_198
timestamp 1676037725
transform 1 0 19320 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_210
timestamp 1676037725
transform 1 0 20424 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1676037725
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_233
timestamp 1676037725
transform 1 0 22540 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_252
timestamp 1676037725
transform 1 0 24288 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_262
timestamp 1676037725
transform 1 0 25208 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1676037725
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1676037725
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1676037725
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_19
timestamp 1676037725
transform 1 0 2852 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1676037725
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_38
timestamp 1676037725
transform 1 0 4600 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_46
timestamp 1676037725
transform 1 0 5336 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_57
timestamp 1676037725
transform 1 0 6348 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_94
timestamp 1676037725
transform 1 0 9752 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_102
timestamp 1676037725
transform 1 0 10488 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_118
timestamp 1676037725
transform 1 0 11960 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_130
timestamp 1676037725
transform 1 0 13064 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_134
timestamp 1676037725
transform 1 0 13432 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1676037725
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_156
timestamp 1676037725
transform 1 0 15456 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_168
timestamp 1676037725
transform 1 0 16560 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1676037725
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1676037725
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_209
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_217
timestamp 1676037725
transform 1 0 21068 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_235
timestamp 1676037725
transform 1 0 22724 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1676037725
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_262
timestamp 1676037725
transform 1 0 25208 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_291
timestamp 1676037725
transform 1 0 27876 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_17
timestamp 1676037725
transform 1 0 2668 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_37
timestamp 1676037725
transform 1 0 4508 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_45
timestamp 1676037725
transform 1 0 5244 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_53
timestamp 1676037725
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_72
timestamp 1676037725
transform 1 0 7728 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_78
timestamp 1676037725
transform 1 0 8280 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_100
timestamp 1676037725
transform 1 0 10304 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_119
timestamp 1676037725
transform 1 0 12052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_123
timestamp 1676037725
transform 1 0 12420 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_131
timestamp 1676037725
transform 1 0 13156 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_137
timestamp 1676037725
transform 1 0 13708 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_162
timestamp 1676037725
transform 1 0 16008 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_196
timestamp 1676037725
transform 1 0 19136 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_203
timestamp 1676037725
transform 1 0 19780 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_210
timestamp 1676037725
transform 1 0 20424 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1676037725
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1676037725
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_240
timestamp 1676037725
transform 1 0 23184 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_253
timestamp 1676037725
transform 1 0 24380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1676037725
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_286
timestamp 1676037725
transform 1 0 27416 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_298
timestamp 1676037725
transform 1 0 28520 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_9
timestamp 1676037725
transform 1 0 1932 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1676037725
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_36
timestamp 1676037725
transform 1 0 4416 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_44
timestamp 1676037725
transform 1 0 5152 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_89
timestamp 1676037725
transform 1 0 9292 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_93
timestamp 1676037725
transform 1 0 9660 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_101
timestamp 1676037725
transform 1 0 10396 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_123
timestamp 1676037725
transform 1 0 12420 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_127
timestamp 1676037725
transform 1 0 12788 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_131
timestamp 1676037725
transform 1 0 13156 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_156
timestamp 1676037725
transform 1 0 15456 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_164
timestamp 1676037725
transform 1 0 16192 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_181
timestamp 1676037725
transform 1 0 17756 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_188
timestamp 1676037725
transform 1 0 18400 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_220
timestamp 1676037725
transform 1 0 21344 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1676037725
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1676037725
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_261
timestamp 1676037725
transform 1 0 25116 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_266
timestamp 1676037725
transform 1 0 25576 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_291
timestamp 1676037725
transform 1 0 27876 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_32
timestamp 1676037725
transform 1 0 4048 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_45
timestamp 1676037725
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1676037725
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_68
timestamp 1676037725
transform 1 0 7360 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_72
timestamp 1676037725
transform 1 0 7728 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_76
timestamp 1676037725
transform 1 0 8096 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_93
timestamp 1676037725
transform 1 0 9660 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1676037725
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_118
timestamp 1676037725
transform 1 0 11960 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_145
timestamp 1676037725
transform 1 0 14444 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_157
timestamp 1676037725
transform 1 0 15548 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_165
timestamp 1676037725
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_177
timestamp 1676037725
transform 1 0 17388 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_189
timestamp 1676037725
transform 1 0 18492 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_197
timestamp 1676037725
transform 1 0 19228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_211
timestamp 1676037725
transform 1 0 20516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1676037725
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_230
timestamp 1676037725
transform 1 0 22264 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_243
timestamp 1676037725
transform 1 0 23460 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_255
timestamp 1676037725
transform 1 0 24564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_263
timestamp 1676037725
transform 1 0 25300 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1676037725
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_286
timestamp 1676037725
transform 1 0 27416 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_290
timestamp 1676037725
transform 1 0 27784 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_297
timestamp 1676037725
transform 1 0 28428 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1676037725
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_57
timestamp 1676037725
transform 1 0 6348 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_100
timestamp 1676037725
transform 1 0 10304 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_113
timestamp 1676037725
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_125
timestamp 1676037725
transform 1 0 12604 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1676037725
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_165
timestamp 1676037725
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_169
timestamp 1676037725
transform 1 0 16652 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_175
timestamp 1676037725
transform 1 0 17204 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_187
timestamp 1676037725
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_217
timestamp 1676037725
transform 1 0 21068 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_223
timestamp 1676037725
transform 1 0 21620 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_225
timestamp 1676037725
transform 1 0 21804 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_230
timestamp 1676037725
transform 1 0 22264 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_242
timestamp 1676037725
transform 1 0 23368 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1676037725
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_261
timestamp 1676037725
transform 1 0 25116 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_273
timestamp 1676037725
transform 1 0 26220 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_279
timestamp 1676037725
transform 1 0 26772 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_281
timestamp 1676037725
transform 1 0 26956 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_287
timestamp 1676037725
transform 1 0 27508 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_297
timestamp 1676037725
transform 1 0 28428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9752 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1676037725
transform 1 0 12328 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1676037725
transform 1 0 4784 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1676037725
transform -1 0 25760 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1676037725
transform -1 0 24104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1676037725
transform -1 0 20700 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1676037725
transform -1 0 19872 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1676037725
transform -1 0 17572 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1676037725
transform -1 0 14996 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1676037725
transform -1 0 13800 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1676037725
transform -1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1676037725
transform -1 0 26220 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1676037725
transform -1 0 27416 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1676037725
transform -1 0 27416 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1676037725
transform -1 0 21344 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1676037725
transform -1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1676037725
transform 1 0 27968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1676037725
transform 1 0 27140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1676037725
transform -1 0 2852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1676037725
transform -1 0 2576 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1676037725
transform -1 0 4784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1676037725
transform -1 0 8372 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1676037725
transform 1 0 11684 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1676037725
transform -1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1676037725
transform -1 0 6348 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1676037725
transform 1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1676037725
transform -1 0 3404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1676037725
transform 1 0 3128 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1676037725
transform -1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1676037725
transform -1 0 25024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1676037725
transform -1 0 22264 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1676037725
transform 1 0 20148 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1676037725
transform 1 0 18124 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1676037725
transform -1 0 19688 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1676037725
transform -1 0 20056 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1676037725
transform -1 0 26220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1676037725
transform -1 0 27416 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1676037725
transform -1 0 27416 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1676037725
transform 1 0 26404 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1676037725
transform 1 0 27140 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1676037725
transform -1 0 27416 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1676037725
transform -1 0 17112 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1676037725
transform -1 0 11960 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1676037725
transform -1 0 13156 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1676037725
transform -1 0 13708 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1676037725
transform 1 0 15272 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1676037725
transform -1 0 4508 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1676037725
transform -1 0 5612 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1676037725
transform -1 0 6072 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1676037725
transform -1 0 6808 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1676037725
transform 1 0 6348 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1676037725
transform -1 0 7360 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1676037725
transform -1 0 9660 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1676037725
transform -1 0 6808 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1676037725
transform 1 0 4784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1676037725
transform -1 0 10948 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1676037725
transform -1 0 2852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1676037725
transform -1 0 2668 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1676037725
transform -1 0 2852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1676037725
transform -1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1676037725
transform -1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _370_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _371_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _372_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16100 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _373_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23276 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1676037725
transform 1 0 23184 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp 1676037725
transform 1 0 23000 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1676037725
transform 1 0 22080 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_8  _377_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4048 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_2  _378_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _379__1
timestamp 1676037725
transform -1 0 12880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379__2
timestamp 1676037725
transform -1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _380_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10580 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _381_
timestamp 1676037725
transform -1 0 14904 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _382_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10672 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _383_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10948 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _384_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _385_
timestamp 1676037725
transform 1 0 7820 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _386_
timestamp 1676037725
transform 1 0 7820 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _387_
timestamp 1676037725
transform -1 0 12880 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _388_
timestamp 1676037725
transform -1 0 12512 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _389_
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _390_
timestamp 1676037725
transform -1 0 14904 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _391_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9568 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _392_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12420 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _393_
timestamp 1676037725
transform 1 0 10580 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _394_
timestamp 1676037725
transform 1 0 9108 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _395_
timestamp 1676037725
transform -1 0 12788 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _396_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_4  _397_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14352 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__o211ai_4  _398_
timestamp 1676037725
transform 1 0 12788 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 1676037725
transform -1 0 14996 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_2  _400_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_2  _401_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8464 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _402_
timestamp 1676037725
transform 1 0 19044 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _403_
timestamp 1676037725
transform -1 0 25208 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _404_
timestamp 1676037725
transform 1 0 18676 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _405_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _406_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _407_
timestamp 1676037725
transform 1 0 24564 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _408_
timestamp 1676037725
transform 1 0 22816 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _409_
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _410_
timestamp 1676037725
transform -1 0 24104 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _411_
timestamp 1676037725
transform -1 0 25024 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _412_
timestamp 1676037725
transform 1 0 23552 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _413_
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _414_
timestamp 1676037725
transform 1 0 20884 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _415_
timestamp 1676037725
transform 1 0 21804 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _416_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _417_
timestamp 1676037725
transform -1 0 25208 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _418_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_4  _419_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14628 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__and3b_1  _420_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _421_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _422_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25484 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _423_
timestamp 1676037725
transform 1 0 6716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _424_
timestamp 1676037725
transform 1 0 6624 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _425_
timestamp 1676037725
transform -1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _426_
timestamp 1676037725
transform -1 0 7820 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _427_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7268 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _428_
timestamp 1676037725
transform 1 0 6348 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _429_
timestamp 1676037725
transform 1 0 6716 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _430_
timestamp 1676037725
transform 1 0 4876 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _431_
timestamp 1676037725
transform -1 0 9752 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _432_
timestamp 1676037725
transform 1 0 10488 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _433_
timestamp 1676037725
transform 1 0 5796 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _434_
timestamp 1676037725
transform -1 0 12420 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _435_
timestamp 1676037725
transform 1 0 10120 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _436_
timestamp 1676037725
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _437_
timestamp 1676037725
transform 1 0 9108 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _438_
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _439_
timestamp 1676037725
transform 1 0 10212 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _440_
timestamp 1676037725
transform -1 0 9660 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _441_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7636 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _442_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11960 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _443_
timestamp 1676037725
transform -1 0 15088 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_4  _444_
timestamp 1676037725
transform -1 0 13800 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__a21boi_1  _445_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_2  _446_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10396 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _447_
timestamp 1676037725
transform 1 0 2300 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _448_
timestamp 1676037725
transform 1 0 17296 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _449_
timestamp 1676037725
transform 1 0 18124 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _450_
timestamp 1676037725
transform -1 0 25208 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _451_
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _452_
timestamp 1676037725
transform 1 0 20056 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _453_
timestamp 1676037725
transform 1 0 16652 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _454_
timestamp 1676037725
transform 1 0 20608 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _455_
timestamp 1676037725
transform 1 0 19044 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _456_
timestamp 1676037725
transform -1 0 19964 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _457_
timestamp 1676037725
transform 1 0 18308 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _458_
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _459_
timestamp 1676037725
transform 1 0 15456 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _460_
timestamp 1676037725
transform 1 0 15364 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _461_
timestamp 1676037725
transform 1 0 17572 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _462_
timestamp 1676037725
transform -1 0 23460 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _463_
timestamp 1676037725
transform -1 0 21528 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _464_
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _465_
timestamp 1676037725
transform 1 0 14996 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _466_
timestamp 1676037725
transform 1 0 14444 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _467_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15456 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _468_
timestamp 1676037725
transform 1 0 27140 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_2  _469_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _470_
timestamp 1676037725
transform 1 0 27140 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _471_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 26404 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _472_
timestamp 1676037725
transform -1 0 28428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _473_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 28428 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _474_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26036 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _475_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _476_
timestamp 1676037725
transform 1 0 27140 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _477_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26680 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _478_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 28428 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _479_
timestamp 1676037725
transform 1 0 27140 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _480_
timestamp 1676037725
transform 1 0 26220 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _481_
timestamp 1676037725
transform 1 0 27232 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _482_
timestamp 1676037725
transform 1 0 27140 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _483_
timestamp 1676037725
transform -1 0 26680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _484_
timestamp 1676037725
transform 1 0 27048 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_2  _485_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24472 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _486_
timestamp 1676037725
transform 1 0 24656 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _487_
timestamp 1676037725
transform -1 0 26404 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _488_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _489_
timestamp 1676037725
transform 1 0 27048 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27692 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_2  _491_
timestamp 1676037725
transform -1 0 26312 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _492_
timestamp 1676037725
transform 1 0 27140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _493_
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _494_
timestamp 1676037725
transform -1 0 20056 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _495_
timestamp 1676037725
transform -1 0 17480 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _496_
timestamp 1676037725
transform 1 0 12420 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _497_
timestamp 1676037725
transform -1 0 13064 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _498_
timestamp 1676037725
transform 1 0 6532 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _499_
timestamp 1676037725
transform 1 0 6532 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _500_
timestamp 1676037725
transform -1 0 9936 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _501_
timestamp 1676037725
transform 1 0 3036 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _502_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5336 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _503_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2668 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _504_
timestamp 1676037725
transform 1 0 4784 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _505_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _506_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4876 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _507_
timestamp 1676037725
transform -1 0 4600 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _508_
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _509_
timestamp 1676037725
transform 1 0 2944 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _510_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4416 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _511_
timestamp 1676037725
transform -1 0 2576 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _512_
timestamp 1676037725
transform 1 0 2944 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _513_
timestamp 1676037725
transform 1 0 4048 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _514_
timestamp 1676037725
transform -1 0 3128 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _515_
timestamp 1676037725
transform 1 0 3680 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _516_
timestamp 1676037725
transform 1 0 4784 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _517_
timestamp 1676037725
transform -1 0 2392 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _518_
timestamp 1676037725
transform 1 0 2760 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _519_
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _520_
timestamp 1676037725
transform 1 0 2760 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _521_
timestamp 1676037725
transform 1 0 15456 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _522_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _523_
timestamp 1676037725
transform 1 0 22632 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _524_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _525_
timestamp 1676037725
transform 1 0 23092 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_4  _526_
timestamp 1676037725
transform -1 0 15732 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2_2  _527_
timestamp 1676037725
transform -1 0 14996 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _528_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _529_
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _530_
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _531_
timestamp 1676037725
transform -1 0 17204 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_2  _532_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10580 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _533_
timestamp 1676037725
transform 1 0 10396 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _534_
timestamp 1676037725
transform 1 0 10764 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _535_
timestamp 1676037725
transform 1 0 11684 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _536_
timestamp 1676037725
transform -1 0 12420 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _537_
timestamp 1676037725
transform 1 0 13892 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _538_
timestamp 1676037725
transform 1 0 12972 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _539_
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _540_
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _541_
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _542_
timestamp 1676037725
transform 1 0 9844 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _543_
timestamp 1676037725
transform 1 0 9936 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _544_
timestamp 1676037725
transform 1 0 11040 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _545_
timestamp 1676037725
transform 1 0 12144 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _546_
timestamp 1676037725
transform 1 0 6072 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _547_
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _548_
timestamp 1676037725
transform 1 0 7360 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _549_
timestamp 1676037725
transform 1 0 11776 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _550_
timestamp 1676037725
transform -1 0 16376 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _551_
timestamp 1676037725
transform -1 0 18952 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _552_
timestamp 1676037725
transform 1 0 17848 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _553_
timestamp 1676037725
transform 1 0 15916 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _554_
timestamp 1676037725
transform 1 0 21252 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _555_
timestamp 1676037725
transform 1 0 22908 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _556_
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _557_
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _558_
timestamp 1676037725
transform 1 0 16376 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _559_
timestamp 1676037725
transform 1 0 21988 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _560_
timestamp 1676037725
transform 1 0 23552 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _561_
timestamp 1676037725
transform 1 0 20424 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _562_
timestamp 1676037725
transform 1 0 23092 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _563_
timestamp 1676037725
transform 1 0 17572 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _564_
timestamp 1676037725
transform 1 0 17296 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _565_
timestamp 1676037725
transform 1 0 17020 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _566_
timestamp 1676037725
transform 1 0 17480 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _567_
timestamp 1676037725
transform -1 0 13340 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _568_
timestamp 1676037725
transform 1 0 9108 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _569_
timestamp 1676037725
transform 1 0 9108 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _570_
timestamp 1676037725
transform 1 0 7820 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _571_
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _572_
timestamp 1676037725
transform -1 0 13616 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _573_
timestamp 1676037725
transform 1 0 7636 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _574_
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _575_
timestamp 1676037725
transform 1 0 9752 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _576_
timestamp 1676037725
transform 1 0 11684 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _577_
timestamp 1676037725
transform 1 0 15824 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _578_
timestamp 1676037725
transform -1 0 17296 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _579_
timestamp 1676037725
transform -1 0 3128 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _580_
timestamp 1676037725
transform -1 0 3496 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _581_
timestamp 1676037725
transform -1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _582_
timestamp 1676037725
transform -1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _583_
timestamp 1676037725
transform -1 0 4232 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _584_
timestamp 1676037725
transform -1 0 5244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _585_
timestamp 1676037725
transform 1 0 6532 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _586_
timestamp 1676037725
transform 1 0 6532 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _587_
timestamp 1676037725
transform 1 0 6164 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _588_
timestamp 1676037725
transform 1 0 5520 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _589_
timestamp 1676037725
transform 1 0 5612 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _590_
timestamp 1676037725
transform -1 0 6072 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _591_
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _592_
timestamp 1676037725
transform 1 0 14260 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _593_
timestamp 1676037725
transform 1 0 14260 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _594_
timestamp 1676037725
transform 1 0 10764 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _595_
timestamp 1676037725
transform 1 0 25484 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _596_
timestamp 1676037725
transform 1 0 27140 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _597_
timestamp 1676037725
transform 1 0 27140 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _598_
timestamp 1676037725
transform 1 0 27140 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _599_
timestamp 1676037725
transform 1 0 25484 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _600_
timestamp 1676037725
transform -1 0 20608 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _601_
timestamp 1676037725
transform 1 0 17296 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _602_
timestamp 1676037725
transform 1 0 19320 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _603_
timestamp 1676037725
transform 1 0 21988 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _604_
timestamp 1676037725
transform 1 0 2300 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _605_
timestamp 1676037725
transform 1 0 3956 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _606_
timestamp 1676037725
transform 1 0 7268 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _607_
timestamp 1676037725
transform 1 0 6256 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _608_
timestamp 1676037725
transform 1 0 9752 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _609_
timestamp 1676037725
transform 1 0 7176 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _610_
timestamp 1676037725
transform 1 0 3956 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _611_
timestamp 1676037725
transform -1 0 3404 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _612_
timestamp 1676037725
transform 1 0 2300 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _613_
timestamp 1676037725
transform 1 0 27140 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _614_
timestamp 1676037725
transform 1 0 25484 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _615_
timestamp 1676037725
transform 1 0 20332 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _616_
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _617_
timestamp 1676037725
transform 1 0 16560 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _618_
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _619_
timestamp 1676037725
transform 1 0 20332 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _620_
timestamp 1676037725
transform 1 0 22908 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _621_
timestamp 1676037725
transform -1 0 26772 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _622_
timestamp 1676037725
transform 1 0 14720 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _623_
timestamp 1676037725
transform -1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _624_
timestamp 1676037725
transform 1 0 17480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _625_
timestamp 1676037725
transform 1 0 19412 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _626_
timestamp 1676037725
transform 1 0 20424 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _627_
timestamp 1676037725
transform -1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _628_
timestamp 1676037725
transform -1 0 22264 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _629_
timestamp 1676037725
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _630_
timestamp 1676037725
transform 1 0 24656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _631_
timestamp 1676037725
transform 1 0 23276 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _632_
timestamp 1676037725
transform -1 0 19320 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _633_
timestamp 1676037725
transform 1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _634_
timestamp 1676037725
transform 1 0 15916 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _635_
timestamp 1676037725
transform -1 0 13708 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _636_
timestamp 1676037725
transform 1 0 13892 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _637_
timestamp 1676037725
transform -1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _638_
timestamp 1676037725
transform 1 0 24840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _639_
timestamp 1676037725
transform -1 0 26496 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _640_
timestamp 1676037725
transform 1 0 26312 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _641_
timestamp 1676037725
transform -1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _642_
timestamp 1676037725
transform -1 0 2484 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _643_
timestamp 1676037725
transform 1 0 2944 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _644_
timestamp 1676037725
transform 1 0 7360 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _645_
timestamp 1676037725
transform 1 0 10396 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _646_
timestamp 1676037725
transform -1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _647_
timestamp 1676037725
transform 1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _648_
timestamp 1676037725
transform -1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _649_
timestamp 1676037725
transform -1 0 4784 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _650_
timestamp 1676037725
transform 1 0 3956 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _651_
timestamp 1676037725
transform -1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _652_
timestamp 1676037725
transform 1 0 25668 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _653_
timestamp 1676037725
transform 1 0 27784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _654_
timestamp 1676037725
transform 1 0 26128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _655_
timestamp 1676037725
transform -1 0 22264 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _656_
timestamp 1676037725
transform -1 0 21068 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _657_
timestamp 1676037725
transform -1 0 19780 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _658_
timestamp 1676037725
transform 1 0 18492 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _659_
timestamp 1676037725
transform 1 0 17756 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _660_
timestamp 1676037725
transform 1 0 24932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _661_
timestamp 1676037725
transform 1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _662_
timestamp 1676037725
transform -1 0 26496 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _663_
timestamp 1676037725
transform -1 0 26680 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _664_
timestamp 1676037725
transform -1 0 26220 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _665_
timestamp 1676037725
transform 1 0 25300 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _666_
timestamp 1676037725
transform 1 0 10396 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _667_
timestamp 1676037725
transform 1 0 12144 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _668_
timestamp 1676037725
transform 1 0 13524 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _669_
timestamp 1676037725
transform -1 0 15732 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _670_
timestamp 1676037725
transform -1 0 7728 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _671_
timestamp 1676037725
transform -1 0 6808 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _672_
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _673_
timestamp 1676037725
transform -1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _674_
timestamp 1676037725
transform -1 0 5520 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _675_
timestamp 1676037725
transform -1 0 6348 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _676_
timestamp 1676037725
transform 1 0 7820 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _677_
timestamp 1676037725
transform 1 0 22356 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _678_
timestamp 1676037725
transform 1 0 22724 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _679_
timestamp 1676037725
transform -1 0 24840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _680_
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _681_
timestamp 1676037725
transform 1 0 5428 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _682_
timestamp 1676037725
transform -1 0 11040 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _683_
timestamp 1676037725
transform 1 0 11960 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _684_
timestamp 1676037725
transform -1 0 3036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _685_
timestamp 1676037725
transform -1 0 2576 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _686_
timestamp 1676037725
transform -1 0 2024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _687_
timestamp 1676037725
transform -1 0 2484 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _688_
timestamp 1676037725
transform -1 0 2208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _689_
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _690_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _691_
timestamp 1676037725
transform 1 0 5704 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _692_
timestamp 1676037725
transform -1 0 9936 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _693_
timestamp 1676037725
transform -1 0 3496 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _694_
timestamp 1676037725
transform 1 0 2576 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _695_
timestamp 1676037725
transform 1 0 3036 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _696_
timestamp 1676037725
transform 1 0 2852 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _697_
timestamp 1676037725
transform 1 0 2024 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _698_
timestamp 1676037725
transform 1 0 2208 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _699_
timestamp 1676037725
transform 1 0 2024 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _700_
timestamp 1676037725
transform 1 0 2024 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _701_
timestamp 1676037725
transform 1 0 16560 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _702_
timestamp 1676037725
transform 1 0 24288 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _703_
timestamp 1676037725
transform 1 0 22632 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _704_
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _705_
timestamp 1676037725
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _706_
timestamp 1676037725
transform 1 0 17572 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _707_
timestamp 1676037725
transform -1 0 20148 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _708_
timestamp 1676037725
transform -1 0 16376 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _709_
timestamp 1676037725
transform 1 0 14720 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _710_
timestamp 1676037725
transform -1 0 13800 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _711_
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _712_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12880 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13984 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _714_
timestamp 1676037725
transform 1 0 15364 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _715_
timestamp 1676037725
transform 1 0 16836 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _716_
timestamp 1676037725
transform 1 0 18124 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _717_
timestamp 1676037725
transform 1 0 19504 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _718_
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _719_
timestamp 1676037725
transform 1 0 20976 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _720_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _721_
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _722_
timestamp 1676037725
transform 1 0 22264 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _723_
timestamp 1676037725
transform 1 0 15732 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _724_
timestamp 1676037725
transform 1 0 22816 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _725_
timestamp 1676037725
transform 1 0 13340 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _726_
timestamp 1676037725
transform 1 0 13248 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _727_
timestamp 1676037725
transform 1 0 16468 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _728_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _729_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _730_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10212 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _731_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _732_
timestamp 1676037725
transform 1 0 11776 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _733_
timestamp 1676037725
transform 1 0 20240 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_2  _734_
timestamp 1676037725
transform 1 0 24748 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _735_
timestamp 1676037725
transform 1 0 22816 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _736_
timestamp 1676037725
transform 1 0 20240 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _737_
timestamp 1676037725
transform 1 0 18952 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _738_
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _739_
timestamp 1676037725
transform 1 0 14076 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _740_
timestamp 1676037725
transform 1 0 14260 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _741_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _742_
timestamp 1676037725
transform 1 0 25668 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _743_
timestamp 1676037725
transform 1 0 26220 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _744_
timestamp 1676037725
transform 1 0 26404 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _745_
timestamp 1676037725
transform 1 0 2300 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _746_
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _747_
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _748_
timestamp 1676037725
transform 1 0 7084 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _749_
timestamp 1676037725
transform -1 0 12604 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _750_
timestamp 1676037725
transform 1 0 9292 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _751_
timestamp 1676037725
transform -1 0 8464 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _752_
timestamp 1676037725
transform 1 0 6716 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _753_
timestamp 1676037725
transform 1 0 3772 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _754_
timestamp 1676037725
transform -1 0 4416 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _755_
timestamp 1676037725
transform 1 0 2116 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_2  _756_
timestamp 1676037725
transform 1 0 23092 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _757_
timestamp 1676037725
transform 1 0 26312 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _758_
timestamp 1676037725
transform -1 0 27876 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _759_
timestamp 1676037725
transform -1 0 27324 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _760_
timestamp 1676037725
transform 1 0 12328 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _761_
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _762_
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _763_
timestamp 1676037725
transform 1 0 11868 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _764_
timestamp 1676037725
transform -1 0 10856 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _765_
timestamp 1676037725
transform -1 0 10948 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _766_
timestamp 1676037725
transform 1 0 10764 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _767_
timestamp 1676037725
transform 1 0 5428 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _768_
timestamp 1676037725
transform 1 0 4416 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _769_
timestamp 1676037725
transform 1 0 6716 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _770_
timestamp 1676037725
transform -1 0 11408 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _771_
timestamp 1676037725
transform 1 0 21712 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _772_
timestamp 1676037725
transform -1 0 21344 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _773_
timestamp 1676037725
transform -1 0 19136 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _774_
timestamp 1676037725
transform 1 0 18584 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _775_
timestamp 1676037725
transform 1 0 18676 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _776_
timestamp 1676037725
transform 1 0 25668 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _777_
timestamp 1676037725
transform 1 0 26496 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _778_
timestamp 1676037725
transform 1 0 26220 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _779_
timestamp 1676037725
transform 1 0 26404 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _780_
timestamp 1676037725
transform -1 0 27876 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _781_
timestamp 1676037725
transform 1 0 25944 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _782_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _783_
timestamp 1676037725
transform 1 0 16468 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _784_
timestamp 1676037725
transform 1 0 19320 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _785_
timestamp 1676037725
transform 1 0 17480 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _786_
timestamp 1676037725
transform 1 0 19688 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _787_
timestamp 1676037725
transform 1 0 22632 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _788_
timestamp 1676037725
transform 1 0 22632 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _789_
timestamp 1676037725
transform 1 0 22632 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _790_
timestamp 1676037725
transform 1 0 21988 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _791_
timestamp 1676037725
transform 1 0 22816 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _792_
timestamp 1676037725
transform 1 0 19964 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _793_
timestamp 1676037725
transform 1 0 21252 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _794_
timestamp 1676037725
transform 1 0 10488 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _795_
timestamp 1676037725
transform 1 0 12512 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _796_
timestamp 1676037725
transform 1 0 14076 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _797_
timestamp 1676037725
transform -1 0 16284 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _798_
timestamp 1676037725
transform 1 0 5520 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _799_
timestamp 1676037725
transform 1 0 6532 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _800_
timestamp 1676037725
transform 1 0 6716 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _801_
timestamp 1676037725
transform 1 0 5336 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _802_
timestamp 1676037725
transform 1 0 6532 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _803_
timestamp 1676037725
transform 1 0 6256 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _804_
timestamp 1676037725
transform 1 0 8372 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_2  _805_
timestamp 1676037725
transform 1 0 15548 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _806_
timestamp 1676037725
transform 1 0 16928 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _807_
timestamp 1676037725
transform 1 0 16836 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _808_
timestamp 1676037725
transform 1 0 17204 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _809_
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _810_
timestamp 1676037725
transform 1 0 9108 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _811_
timestamp 1676037725
transform 1 0 7176 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _812_
timestamp 1676037725
transform -1 0 11960 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _813_
timestamp 1676037725
transform 1 0 7084 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _814_
timestamp 1676037725
transform 1 0 6716 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _815_
timestamp 1676037725
transform 1 0 9384 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _816_
timestamp 1676037725
transform 1 0 10396 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _817_
timestamp 1676037725
transform 1 0 16284 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _818_
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _819_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _820_
timestamp 1676037725
transform 1 0 22264 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _821_
timestamp 1676037725
transform 1 0 22172 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _822_
timestamp 1676037725
transform 1 0 22816 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _823_
timestamp 1676037725
transform 1 0 5612 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _824_
timestamp 1676037725
transform -1 0 6164 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _825_
timestamp 1676037725
transform 1 0 11684 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _826_
timestamp 1676037725
transform 1 0 2576 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _827_
timestamp 1676037725
transform 1 0 2024 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _828_
timestamp 1676037725
transform 1 0 1932 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _829_
timestamp 1676037725
transform 1 0 2024 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _830_
timestamp 1676037725
transform 1 0 1564 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _831_
timestamp 1676037725
transform 1 0 7912 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__203_
timestamp 1676037725
transform -1 0 12052 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__222_
timestamp 1676037725
transform 1 0 22632 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__245_
timestamp 1676037725
transform -1 0 8556 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__264_
timestamp 1676037725
transform 1 0 21068 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1676037725
transform 1 0 3956 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__183_
timestamp 1676037725
transform -1 0 14812 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__203_
timestamp 1676037725
transform -1 0 9660 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__222_
timestamp 1676037725
transform -1 0 22632 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__245_
timestamp 1676037725
transform -1 0 6072 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__264_
timestamp 1676037725
transform -1 0 20056 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1676037725
transform -1 0 3404 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__183_
timestamp 1676037725
transform -1 0 14812 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__203_
timestamp 1676037725
transform 1 0 10396 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__222_
timestamp 1676037725
transform 1 0 23368 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__245_
timestamp 1676037725
transform 1 0 4508 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__264_
timestamp 1676037725
transform 1 0 19688 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11316 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout17
timestamp 1676037725
transform -1 0 11868 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  fanout18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5428 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  fanout19
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  fanout20
timestamp 1676037725
transform -1 0 5612 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  fanout21
timestamp 1676037725
transform -1 0 20884 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  fanout22
timestamp 1676037725
transform -1 0 18308 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  fanout23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5244 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout24
timestamp 1676037725
transform 1 0 9660 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout25
timestamp 1676037725
transform -1 0 4416 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10304 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22172 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout28
timestamp 1676037725
transform -1 0 12604 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout29
timestamp 1676037725
transform 1 0 19688 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout30
timestamp 1676037725
transform 1 0 12788 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout31
timestamp 1676037725
transform 1 0 13248 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout32
timestamp 1676037725
transform -1 0 4508 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout33
timestamp 1676037725
transform 1 0 3956 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout34
timestamp 1676037725
transform -1 0 5244 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  fanout35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15456 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout36
timestamp 1676037725
transform -1 0 15272 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout37
timestamp 1676037725
transform -1 0 13800 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout38
timestamp 1676037725
transform 1 0 16836 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__bufbuf_16  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold2
timestamp 1676037725
transform 1 0 7268 0 -1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__buf_6  input1
timestamp 1676037725
transform 1 0 9476 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input2
timestamp 1676037725
transform 1 0 12972 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17204 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1676037725
transform 1 0 20516 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1676037725
transform 1 0 24564 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input6
timestamp 1676037725
transform 1 0 27600 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 1676037725
transform 1 0 6532 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output8
timestamp 1676037725
transform 1 0 27876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output9
timestamp 1676037725
transform 1 0 27876 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output10
timestamp 1676037725
transform 1 0 27876 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output11
timestamp 1676037725
transform 1 0 27876 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1676037725
transform 1 0 27876 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output13
timestamp 1676037725
transform 1 0 27876 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output14
timestamp 1676037725
transform 1 0 27876 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output15
timestamp 1676037725
transform 1 0 27876 0 -1 27200
box -38 -48 590 592
<< labels >>
flabel metal2 s 2042 29200 2098 30000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 9402 29200 9458 30000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 13082 29200 13138 30000 0 FreeSans 224 90 0 0 io_in[1]
port 2 nsew signal input
flabel metal2 s 16762 29200 16818 30000 0 FreeSans 224 90 0 0 io_in[2]
port 3 nsew signal input
flabel metal2 s 20442 29200 20498 30000 0 FreeSans 224 90 0 0 io_in[3]
port 4 nsew signal input
flabel metal2 s 24122 29200 24178 30000 0 FreeSans 224 90 0 0 io_in[4]
port 5 nsew signal input
flabel metal2 s 27802 29200 27858 30000 0 FreeSans 224 90 0 0 io_in[5]
port 6 nsew signal input
flabel metal3 s 29200 2048 30000 2168 0 FreeSans 480 0 0 0 io_out[0]
port 7 nsew signal tristate
flabel metal3 s 29200 5720 30000 5840 0 FreeSans 480 0 0 0 io_out[1]
port 8 nsew signal tristate
flabel metal3 s 29200 9392 30000 9512 0 FreeSans 480 0 0 0 io_out[2]
port 9 nsew signal tristate
flabel metal3 s 29200 13064 30000 13184 0 FreeSans 480 0 0 0 io_out[3]
port 10 nsew signal tristate
flabel metal3 s 29200 16736 30000 16856 0 FreeSans 480 0 0 0 io_out[4]
port 11 nsew signal tristate
flabel metal3 s 29200 20408 30000 20528 0 FreeSans 480 0 0 0 io_out[5]
port 12 nsew signal tristate
flabel metal3 s 29200 24080 30000 24200 0 FreeSans 480 0 0 0 io_out[6]
port 13 nsew signal tristate
flabel metal3 s 29200 27752 30000 27872 0 FreeSans 480 0 0 0 io_out[7]
port 14 nsew signal tristate
flabel metal2 s 5722 29200 5778 30000 0 FreeSans 224 90 0 0 rst
port 15 nsew signal input
flabel metal4 s 4417 2128 4737 27792 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 11363 2128 11683 27792 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 18309 2128 18629 27792 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 25255 2128 25575 27792 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 7890 2128 8210 27792 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 14836 2128 15156 27792 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 21782 2128 22102 27792 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 28728 2128 29048 27792 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
