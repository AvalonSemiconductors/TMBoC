VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_as2650
  CLASS BLOCK ;
  FOREIGN wrapped_as2650 ;
  ORIGIN 0.000 0.000 ;
  SIZE 425.000 BY 400.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END io_in[7]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.720 4.000 307.320 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 4.000 335.880 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END io_out[26]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END io_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 389.200 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 419.060 389.045 ;
      LAYER met1 ;
        RECT 4.670 10.640 419.060 389.200 ;
      LAYER met2 ;
        RECT 4.690 4.280 415.280 392.885 ;
        RECT 4.690 4.000 21.430 4.280 ;
        RECT 22.270 4.000 63.750 4.280 ;
        RECT 64.590 4.000 106.070 4.280 ;
        RECT 106.910 4.000 148.390 4.280 ;
        RECT 149.230 4.000 190.710 4.280 ;
        RECT 191.550 4.000 233.030 4.280 ;
        RECT 233.870 4.000 275.350 4.280 ;
        RECT 276.190 4.000 317.670 4.280 ;
        RECT 318.510 4.000 359.990 4.280 ;
        RECT 360.830 4.000 402.310 4.280 ;
        RECT 403.150 4.000 415.280 4.280 ;
      LAYER met3 ;
        RECT 4.400 392.000 406.630 392.865 ;
        RECT 4.000 379.120 406.630 392.000 ;
        RECT 4.400 377.720 406.630 379.120 ;
        RECT 4.000 364.840 406.630 377.720 ;
        RECT 4.400 363.440 406.630 364.840 ;
        RECT 4.000 350.560 406.630 363.440 ;
        RECT 4.400 349.160 406.630 350.560 ;
        RECT 4.000 336.280 406.630 349.160 ;
        RECT 4.400 334.880 406.630 336.280 ;
        RECT 4.000 322.000 406.630 334.880 ;
        RECT 4.400 320.600 406.630 322.000 ;
        RECT 4.000 307.720 406.630 320.600 ;
        RECT 4.400 306.320 406.630 307.720 ;
        RECT 4.000 293.440 406.630 306.320 ;
        RECT 4.400 292.040 406.630 293.440 ;
        RECT 4.000 279.160 406.630 292.040 ;
        RECT 4.400 277.760 406.630 279.160 ;
        RECT 4.000 264.880 406.630 277.760 ;
        RECT 4.400 263.480 406.630 264.880 ;
        RECT 4.000 250.600 406.630 263.480 ;
        RECT 4.400 249.200 406.630 250.600 ;
        RECT 4.000 236.320 406.630 249.200 ;
        RECT 4.400 234.920 406.630 236.320 ;
        RECT 4.000 222.040 406.630 234.920 ;
        RECT 4.400 220.640 406.630 222.040 ;
        RECT 4.000 207.760 406.630 220.640 ;
        RECT 4.400 206.360 406.630 207.760 ;
        RECT 4.000 193.480 406.630 206.360 ;
        RECT 4.400 192.080 406.630 193.480 ;
        RECT 4.000 179.200 406.630 192.080 ;
        RECT 4.400 177.800 406.630 179.200 ;
        RECT 4.000 164.920 406.630 177.800 ;
        RECT 4.400 163.520 406.630 164.920 ;
        RECT 4.000 150.640 406.630 163.520 ;
        RECT 4.400 149.240 406.630 150.640 ;
        RECT 4.000 136.360 406.630 149.240 ;
        RECT 4.400 134.960 406.630 136.360 ;
        RECT 4.000 122.080 406.630 134.960 ;
        RECT 4.400 120.680 406.630 122.080 ;
        RECT 4.000 107.800 406.630 120.680 ;
        RECT 4.400 106.400 406.630 107.800 ;
        RECT 4.000 93.520 406.630 106.400 ;
        RECT 4.400 92.120 406.630 93.520 ;
        RECT 4.000 79.240 406.630 92.120 ;
        RECT 4.400 77.840 406.630 79.240 ;
        RECT 4.000 64.960 406.630 77.840 ;
        RECT 4.400 63.560 406.630 64.960 ;
        RECT 4.000 50.680 406.630 63.560 ;
        RECT 4.400 49.280 406.630 50.680 ;
        RECT 4.000 36.400 406.630 49.280 ;
        RECT 4.400 35.000 406.630 36.400 ;
        RECT 4.000 22.120 406.630 35.000 ;
        RECT 4.400 20.720 406.630 22.120 ;
        RECT 4.000 7.840 406.630 20.720 ;
        RECT 4.400 6.975 406.630 7.840 ;
      LAYER met4 ;
        RECT 11.335 55.255 20.640 318.745 ;
        RECT 23.040 55.255 97.440 318.745 ;
        RECT 99.840 55.255 174.240 318.745 ;
        RECT 176.640 55.255 251.040 318.745 ;
        RECT 253.440 55.255 318.025 318.745 ;
  END
END wrapped_as2650
END LIBRARY

