magic
tech sky130B
magscale 1 2
timestamp 1680008313
<< nwell >>
rect 1066 20933 22854 21499
rect 1066 19845 22854 20411
rect 1066 18757 22854 19323
rect 1066 17669 22854 18235
rect 1066 16581 22854 17147
rect 1066 15493 22854 16059
rect 1066 14405 22854 14971
rect 1066 13317 22854 13883
rect 1066 12229 22854 12795
rect 1066 11141 22854 11707
rect 1066 10053 22854 10619
rect 1066 8965 22854 9531
rect 1066 7877 22854 8443
rect 1066 6789 22854 7355
rect 1066 5701 22854 6267
rect 1066 4613 22854 5179
rect 1066 3525 22854 4091
rect 1066 2437 22854 3003
<< obsli1 >>
rect 1104 2159 22816 21777
<< obsm1 >>
rect 1104 2128 22976 21808
<< metal2 >>
rect 3974 23200 4030 24000
rect 11978 23200 12034 24000
rect 19982 23200 20038 24000
rect 1674 0 1730 800
rect 4618 0 4674 800
rect 7562 0 7618 800
rect 10506 0 10562 800
rect 13450 0 13506 800
rect 16394 0 16450 800
rect 19338 0 19394 800
rect 22282 0 22338 800
<< obsm2 >>
rect 1676 23144 3918 23338
rect 4086 23144 11922 23338
rect 12090 23144 19926 23338
rect 20094 23144 22970 23338
rect 1676 856 22970 23144
rect 1786 800 4562 856
rect 4730 800 7506 856
rect 7674 800 10450 856
rect 10618 800 13394 856
rect 13562 800 16338 856
rect 16506 800 19282 856
rect 19450 800 22226 856
rect 22394 800 22970 856
<< obsm3 >>
rect 3660 2143 22974 21793
<< metal4 >>
rect 3658 2128 3978 21808
rect 6372 2128 6692 21808
rect 9086 2128 9406 21808
rect 11800 2128 12120 21808
rect 14514 2128 14834 21808
rect 17228 2128 17548 21808
rect 19942 2128 20262 21808
rect 22656 2128 22976 21808
<< labels >>
rlabel metal2 s 3974 23200 4030 24000 6 clk
port 1 nsew signal input
rlabel metal2 s 19982 23200 20038 24000 6 io_in
port 2 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 io_out[0]
port 3 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 io_out[1]
port 4 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 io_out[2]
port 5 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 io_out[3]
port 6 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 io_out[4]
port 7 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 io_out[5]
port 8 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 io_out[6]
port 9 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 io_out[7]
port 10 nsew signal output
rlabel metal2 s 11978 23200 12034 24000 6 rst
port 11 nsew signal input
rlabel metal4 s 3658 2128 3978 21808 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 9086 2128 9406 21808 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 14514 2128 14834 21808 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 19942 2128 20262 21808 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 6372 2128 6692 21808 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 11800 2128 12120 21808 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 17228 2128 17548 21808 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 22656 2128 22976 21808 6 vssd1
port 13 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 24000 24000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1282772
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/Diceroll/runs/23_03_28_14_57/results/signoff/tt2_tholin_diceroll.magic.gds
string GDS_START 520274
<< end >>

