* NGSPICE file created from posit_unit.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

.subckt posit_unit clk io_in[0] io_in[1] io_in[2] io_out[0] io_out[1] io_out[2] io_out[3]
+ rst vccd1 vssd1
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7963_ _8046_/Q _7964_/C _7962_/Y vssd1 vssd1 vccd1 vccd1 _8046_/D sky130_fd_sc_hd__a21oi_1
XFILLER_82_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6914_ _6914_/A _6914_/B vssd1 vssd1 vccd1 vccd1 _6923_/A sky130_fd_sc_hd__xnor2_4
X_7894_ _7894_/A _7894_/B vssd1 vssd1 vccd1 vccd1 _7895_/C sky130_fd_sc_hd__or2_1
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6845_ _6845_/A _6845_/B vssd1 vssd1 vccd1 vccd1 _6866_/B sky130_fd_sc_hd__xor2_4
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6776_ _6776_/A _6776_/B vssd1 vssd1 vccd1 vccd1 _6776_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5727_ _5728_/A _5728_/B vssd1 vssd1 vccd1 vccd1 _5727_/X sky130_fd_sc_hd__and2_1
X_5658_ _5662_/B _5662_/A vssd1 vssd1 vccd1 vccd1 _5658_/Y sky130_fd_sc_hd__nand2b_1
X_5589_ _5589_/A _5589_/B vssd1 vssd1 vccd1 vccd1 _5643_/B sky130_fd_sc_hd__xnor2_4
X_4609_ _7001_/A _4605_/B _4603_/Y vssd1 vssd1 vccd1 vccd1 _4611_/B sky130_fd_sc_hd__o21ai_4
X_7328_ _7328_/A _7328_/B vssd1 vssd1 vccd1 vccd1 _7345_/A sky130_fd_sc_hd__or2_4
X_7259_ _7263_/A _7263_/B vssd1 vssd1 vccd1 vccd1 _7259_/X sky130_fd_sc_hd__and2b_1
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4960_ _4960_/A _4960_/B vssd1 vssd1 vccd1 vccd1 _4995_/B sky130_fd_sc_hd__xor2_4
XFILLER_83_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4891_ _5013_/C _4991_/A vssd1 vssd1 vccd1 vccd1 _4892_/B sky130_fd_sc_hd__nand2b_4
X_6630_ _6749_/S vssd1 vssd1 vccd1 vccd1 _7616_/S sky130_fd_sc_hd__clkinv_4
X_6561_ _6548_/B _6556_/B _6540_/B vssd1 vssd1 vccd1 vccd1 _6562_/B sky130_fd_sc_hd__a21oi_1
X_5512_ _5303_/Y _5566_/A _5511_/X vssd1 vssd1 vccd1 vccd1 _5563_/B sky130_fd_sc_hd__a21oi_4
XFILLER_118_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6492_ _6492_/A _6492_/B vssd1 vssd1 vccd1 vccd1 _6495_/B sky130_fd_sc_hd__nor2_1
X_5443_ _5443_/A _5443_/B vssd1 vssd1 vccd1 vccd1 _5451_/A sky130_fd_sc_hd__xor2_4
X_5374_ _5541_/A _5796_/B vssd1 vssd1 vccd1 vccd1 _5375_/B sky130_fd_sc_hd__nor2_4
X_4325_ _4322_/X _4323_/X _4324_/X vssd1 vssd1 vccd1 vccd1 _4325_/Y sky130_fd_sc_hd__o21ai_2
X_7113_ _7334_/B _7235_/B vssd1 vssd1 vccd1 vccd1 _7113_/X sky130_fd_sc_hd__or2_1
XFILLER_99_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout138 _7294_/A vssd1 vssd1 vccd1 vccd1 _4662_/A sky130_fd_sc_hd__clkbuf_16
Xfanout105 _5362_/Y vssd1 vssd1 vccd1 vccd1 _7366_/B sky130_fd_sc_hd__buf_8
Xfanout116 _4920_/A vssd1 vssd1 vccd1 vccd1 _4991_/A sky130_fd_sc_hd__buf_8
Xfanout127 _4320_/X vssd1 vssd1 vccd1 vccd1 _6916_/A sky130_fd_sc_hd__buf_8
XFILLER_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4256_ _4356_/A _4406_/A vssd1 vssd1 vccd1 vccd1 _4256_/Y sky130_fd_sc_hd__nor2_1
Xfanout149 _4334_/Y vssd1 vssd1 vccd1 vccd1 _7012_/A sky130_fd_sc_hd__buf_4
X_7044_ _7045_/B _7045_/A vssd1 vssd1 vccd1 vccd1 _7048_/B sky130_fd_sc_hd__nand2b_1
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4187_ _4216_/B _4187_/B vssd1 vssd1 vccd1 vccd1 _4193_/A sky130_fd_sc_hd__xnor2_4
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7946_ _7649_/A _6774_/C _6771_/X vssd1 vssd1 vccd1 vccd1 _7947_/C sky130_fd_sc_hd__o21ai_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7877_ _7876_/X _7877_/B vssd1 vssd1 vccd1 vccd1 _7877_/X sky130_fd_sc_hd__and2b_1
X_6828_ _6828_/A _6828_/B vssd1 vssd1 vccd1 vccd1 _7392_/C sky130_fd_sc_hd__nor2_1
XFILLER_11_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6759_ _6757_/D _7788_/B _7718_/S vssd1 vssd1 vccd1 vccd1 _7580_/C sky130_fd_sc_hd__mux2_2
XFILLER_11_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4110_ _4111_/A _6018_/A vssd1 vssd1 vccd1 vccd1 _4110_/Y sky130_fd_sc_hd__nor2_2
X_5090_ _5090_/A _5090_/B vssd1 vssd1 vccd1 vccd1 _5090_/X sky130_fd_sc_hd__and2_1
X_4041_ _8058_/Q _4052_/B vssd1 vssd1 vccd1 vccd1 _4080_/B sky130_fd_sc_hd__or2_4
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5992_ _5995_/A vssd1 vssd1 vccd1 vccd1 _6018_/B sky130_fd_sc_hd__inv_2
X_7800_ _7817_/A _7800_/B vssd1 vssd1 vccd1 vccd1 _7874_/B sky130_fd_sc_hd__and2_4
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7731_ _7731_/A _7731_/B _7703_/B vssd1 vssd1 vccd1 vccd1 _7757_/B sky130_fd_sc_hd__nor3b_1
X_4943_ _4976_/A _4976_/B _4940_/Y vssd1 vssd1 vccd1 vccd1 _4945_/B sky130_fd_sc_hd__a21oi_4
XFILLER_17_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7662_ _7837_/A _7684_/A _7684_/B _7802_/B2 vssd1 vssd1 vccd1 vccd1 _7663_/B sky130_fd_sc_hd__a31o_1
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6613_ _6615_/A _6613_/B vssd1 vssd1 vccd1 vccd1 _6616_/C sky130_fd_sc_hd__xor2_2
X_4874_ _4874_/A _4874_/B vssd1 vssd1 vccd1 vccd1 _4876_/A sky130_fd_sc_hd__or2_4
XFILLER_20_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7593_ _7657_/B _7460_/X _7592_/Y vssd1 vssd1 vccd1 vccd1 _7594_/A sky130_fd_sc_hd__o21ai_2
XFILLER_118_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6544_ _6457_/X _6500_/Y _6544_/S vssd1 vssd1 vccd1 vccd1 _6545_/B sky130_fd_sc_hd__mux2_4
X_6475_ _6475_/A _6475_/B vssd1 vssd1 vccd1 vccd1 _6475_/X sky130_fd_sc_hd__or2_2
X_5426_ _5426_/A _5426_/B vssd1 vssd1 vccd1 vccd1 _5556_/B sky130_fd_sc_hd__xor2_2
XFILLER_114_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5357_ _5357_/A _5357_/B vssd1 vssd1 vccd1 vccd1 _5358_/B sky130_fd_sc_hd__xor2_4
XFILLER_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8076_ _8077_/CLK _8076_/D vssd1 vssd1 vccd1 vccd1 _8076_/Q sky130_fd_sc_hd__dfxtp_4
X_5288_ _5288_/A _5288_/B vssd1 vssd1 vccd1 vccd1 _6173_/A sky130_fd_sc_hd__nand2_1
X_4308_ _4302_/X _5322_/B _5322_/A vssd1 vssd1 vccd1 vccd1 _4308_/X sky130_fd_sc_hd__mux2_4
XFILLER_75_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4239_ _4322_/A _4239_/B _4239_/C vssd1 vssd1 vccd1 vccd1 _4239_/Y sky130_fd_sc_hd__nand3_1
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7027_ _7027_/A _7344_/B _7027_/C vssd1 vssd1 vccd1 vccd1 _7084_/A sky130_fd_sc_hd__or3_4
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7929_ _7929_/A _7929_/B vssd1 vssd1 vccd1 vccd1 _7929_/X sky130_fd_sc_hd__or2_1
XFILLER_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4590_ _7116_/A _5033_/A vssd1 vssd1 vccd1 vccd1 _4594_/A sky130_fd_sc_hd__nor2_2
XFILLER_115_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6260_ _7930_/A _7639_/B _6259_/X vssd1 vssd1 vccd1 vccd1 _6260_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6191_ _6081_/Y _6111_/B _6111_/C _6151_/X vssd1 vssd1 vccd1 vccd1 _6200_/B sky130_fd_sc_hd__a31o_1
X_5211_ _5151_/C _5264_/A _6783_/A _5210_/X vssd1 vssd1 vccd1 vccd1 _5212_/B sky130_fd_sc_hd__o31a_4
X_5142_ _5166_/B _6807_/A _5208_/A vssd1 vssd1 vccd1 vccd1 _5172_/A sky130_fd_sc_hd__and3_1
XFILLER_96_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5073_ _5074_/B _5074_/C _5074_/A vssd1 vssd1 vccd1 vccd1 _5352_/A sky130_fd_sc_hd__a21o_4
X_4024_ _8013_/Q _8014_/Q _7955_/S vssd1 vssd1 vccd1 vccd1 _8014_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5975_ _4050_/Y _4303_/C _4130_/X _4303_/B vssd1 vssd1 vccd1 vccd1 _5975_/X sky130_fd_sc_hd__o211a_1
X_7714_ _7837_/A _7744_/A _7744_/B vssd1 vssd1 vccd1 vccd1 _7714_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4926_ _4926_/A _4963_/A vssd1 vssd1 vccd1 vccd1 _4936_/A sky130_fd_sc_hd__nor2_4
X_7645_ _7607_/B _7612_/X _7607_/A vssd1 vssd1 vccd1 vccd1 _7645_/X sky130_fd_sc_hd__o21a_1
X_4857_ _4857_/A _4867_/A _4857_/C vssd1 vssd1 vccd1 vccd1 _4858_/B sky130_fd_sc_hd__and3_1
X_7576_ _7576_/A _7611_/B vssd1 vssd1 vccd1 vccd1 _7576_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6527_ _6527_/A _6527_/B vssd1 vssd1 vccd1 vccd1 _6539_/A sky130_fd_sc_hd__xnor2_4
X_4788_ _4783_/B _4832_/A vssd1 vssd1 vccd1 vccd1 _4789_/B sky130_fd_sc_hd__and2b_1
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6458_ _6446_/Y _6457_/X _6480_/B vssd1 vssd1 vccd1 vccd1 _6541_/B sky130_fd_sc_hd__o21a_2
XFILLER_69_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6389_ _6379_/X _6388_/X _6431_/S vssd1 vssd1 vccd1 vccd1 _6390_/B sky130_fd_sc_hd__mux2_1
X_5409_ _5410_/A _5410_/B vssd1 vssd1 vccd1 vccd1 _5409_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8059_ _8077_/CLK _8059_/D vssd1 vssd1 vccd1 vccd1 _8059_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5760_ _5759_/A _5759_/B _5759_/C vssd1 vssd1 vccd1 vccd1 _5761_/C sky130_fd_sc_hd__a21o_2
XFILLER_91_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _5692_/B _5691_/B vssd1 vssd1 vccd1 vccd1 _5695_/A sky130_fd_sc_hd__nand2_4
X_4711_ _4689_/A _4689_/B _4689_/C vssd1 vssd1 vccd1 vccd1 _4712_/B sky130_fd_sc_hd__a21oi_1
X_7430_ _7430_/A _7430_/B vssd1 vssd1 vccd1 vccd1 _7430_/X sky130_fd_sc_hd__or2_1
X_4642_ _4642_/A _4642_/B vssd1 vssd1 vccd1 vccd1 _4644_/B sky130_fd_sc_hd__nor2_4
XFILLER_30_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7361_ _7359_/A _7370_/A _7369_/A _7364_/A vssd1 vssd1 vccd1 vccd1 _7374_/B sky130_fd_sc_hd__a31o_2
X_4573_ _4574_/A _4574_/B _4574_/C vssd1 vssd1 vccd1 vccd1 _4573_/Y sky130_fd_sc_hd__nor3_2
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout7 _6166_/S vssd1 vssd1 vccd1 vccd1 _6226_/S sky130_fd_sc_hd__buf_2
X_6312_ _6349_/B _6766_/S _6311_/Y vssd1 vssd1 vccd1 vccd1 _6590_/A sky130_fd_sc_hd__a21o_2
X_7292_ _7300_/A _7300_/B vssd1 vssd1 vccd1 vccd1 _7293_/B sky130_fd_sc_hd__and2b_1
XFILLER_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6243_ _5897_/Y _6239_/B _6238_/X _6242_/X vssd1 vssd1 vccd1 vccd1 _6243_/X sky130_fd_sc_hd__a211o_2
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6174_ _6174_/A _6174_/B vssd1 vssd1 vccd1 vccd1 _6175_/A sky130_fd_sc_hd__or2_1
XFILLER_111_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5125_ _5198_/B _5386_/A vssd1 vssd1 vccd1 vccd1 _5165_/B sky130_fd_sc_hd__or2_1
X_5056_ _5247_/B _5247_/C _5247_/A vssd1 vssd1 vccd1 vccd1 _5248_/A sky130_fd_sc_hd__a21oi_4
X_4007_ _6770_/A vssd1 vssd1 vccd1 vccd1 _7949_/A sky130_fd_sc_hd__inv_2
XFILLER_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5958_ _5959_/A _5959_/B _5959_/C vssd1 vssd1 vccd1 vccd1 _5960_/A sky130_fd_sc_hd__a21o_1
XFILLER_40_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4909_ _4909_/A _4909_/B vssd1 vssd1 vccd1 vccd1 _4916_/B sky130_fd_sc_hd__xor2_4
XFILLER_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5889_ _5889_/A _5889_/B vssd1 vssd1 vccd1 vccd1 _5902_/B sky130_fd_sc_hd__xnor2_4
X_7628_ _7629_/A _7629_/B vssd1 vssd1 vccd1 vccd1 _7687_/A sky130_fd_sc_hd__nor2_4
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7559_ _7554_/B _7590_/A _7939_/A vssd1 vssd1 vccd1 vccd1 _7559_/X sky130_fd_sc_hd__and3b_1
XFILLER_107_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_5 _7306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6930_ _6925_/A _6925_/B _6912_/X vssd1 vssd1 vccd1 vccd1 _6939_/A sky130_fd_sc_hd__a21bo_2
X_6861_ _6861_/A _6861_/B vssd1 vssd1 vccd1 vccd1 _6892_/A sky130_fd_sc_hd__xnor2_2
X_6792_ _6916_/A _5782_/A _5128_/Y vssd1 vssd1 vccd1 vccd1 _6793_/B sky130_fd_sc_hd__a21oi_1
X_5812_ _5817_/A _5817_/B vssd1 vssd1 vccd1 vccd1 _5815_/B sky130_fd_sc_hd__nand2b_1
X_5743_ _5743_/A _5743_/B vssd1 vssd1 vccd1 vccd1 _5746_/B sky130_fd_sc_hd__xnor2_4
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5674_ _5723_/A _7285_/B vssd1 vssd1 vccd1 vccd1 _5724_/A sky130_fd_sc_hd__nand2_2
X_7413_ _7413_/A _7413_/B vssd1 vssd1 vccd1 vccd1 _7421_/B sky130_fd_sc_hd__xor2_4
X_4625_ _4625_/A _4625_/B _4625_/C vssd1 vssd1 vccd1 vccd1 _4660_/A sky130_fd_sc_hd__and3_2
X_7344_ _7371_/A _7344_/B vssd1 vssd1 vccd1 vccd1 _7349_/A sky130_fd_sc_hd__nor2_2
X_4556_ _4556_/A _4556_/B vssd1 vssd1 vccd1 vccd1 _4563_/A sky130_fd_sc_hd__xnor2_4
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7275_ _7275_/A _7275_/B vssd1 vssd1 vccd1 vccd1 _7293_/A sky130_fd_sc_hd__xor2_2
X_4487_ _4501_/A _4480_/X _4481_/X _4486_/X _6916_/A vssd1 vssd1 vccd1 vccd1 _4487_/X
+ sky130_fd_sc_hd__a311o_4
X_6226_ _6165_/Y _6184_/X _6226_/S vssd1 vssd1 vccd1 vccd1 _6226_/X sky130_fd_sc_hd__mux2_2
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6157_ _7269_/B _5969_/Y _6146_/A _6148_/Y _6156_/Y vssd1 vssd1 vccd1 vccd1 _6163_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _5582_/A _7046_/B vssd1 vssd1 vccd1 vccd1 _5156_/C sky130_fd_sc_hd__or2_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6088_ _6088_/A _6088_/B vssd1 vssd1 vccd1 vccd1 _6088_/Y sky130_fd_sc_hd__nand2_2
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5039_ _5039_/A _5039_/B vssd1 vssd1 vccd1 vccd1 _5039_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4410_ _4360_/A _4401_/X _4404_/Y _4409_/X vssd1 vssd1 vccd1 vccd1 _4411_/B sky130_fd_sc_hd__o22a_1
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5390_ _5391_/A _5391_/B vssd1 vssd1 vccd1 vccd1 _5422_/A sky130_fd_sc_hd__nand2_4
X_4341_ _4341_/A1 _4266_/A _4266_/B _4267_/X _4354_/A vssd1 vssd1 vccd1 vccd1 _6951_/A
+ sky130_fd_sc_hd__a311oi_4
X_4272_ _4180_/Y _4259_/B _4271_/X vssd1 vssd1 vccd1 vccd1 _4272_/Y sky130_fd_sc_hd__a21oi_1
X_7060_ _7072_/A _7072_/B _7059_/X vssd1 vssd1 vccd1 vccd1 _7112_/B sky130_fd_sc_hd__o21ba_1
XFILLER_113_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6011_ _6310_/B _6011_/B vssd1 vssd1 vccd1 vccd1 _6012_/B sky130_fd_sc_hd__xnor2_4
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7962_ _8046_/Q _7964_/C _7971_/B vssd1 vssd1 vccd1 vccd1 _7962_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_94_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6913_ _6913_/A _6913_/B vssd1 vssd1 vccd1 vccd1 _6925_/A sky130_fd_sc_hd__xnor2_2
X_7893_ _7939_/A _7877_/B _7891_/Y _7892_/Y _7918_/B vssd1 vssd1 vccd1 vccd1 _7893_/X
+ sky130_fd_sc_hd__a311o_1
X_6844_ _6878_/C _7114_/B vssd1 vssd1 vccd1 vccd1 _6866_/A sky130_fd_sc_hd__nand2_4
XFILLER_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6775_ _7580_/C _7579_/A _7935_/A _7923_/A vssd1 vssd1 vccd1 vccd1 _6776_/B sky130_fd_sc_hd__o31a_1
XFILLER_22_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5726_ _5726_/A _5726_/B vssd1 vssd1 vccd1 vccd1 _5728_/B sky130_fd_sc_hd__xor2_4
XFILLER_22_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5657_ _5657_/A _5657_/B vssd1 vssd1 vccd1 vccd1 _5662_/B sky130_fd_sc_hd__xnor2_4
X_5588_ _5588_/A _5588_/B vssd1 vssd1 vccd1 vccd1 _5589_/B sky130_fd_sc_hd__xor2_4
X_4608_ _4606_/A _4606_/Y _4607_/Y _4574_/X vssd1 vssd1 vccd1 vccd1 _4611_/A sky130_fd_sc_hd__o211ai_4
X_7327_ _7327_/A _7327_/B vssd1 vssd1 vccd1 vccd1 _7328_/B sky130_fd_sc_hd__and2_1
X_4539_ _4662_/A _4539_/B vssd1 vssd1 vccd1 vccd1 _4540_/B sky130_fd_sc_hd__xnor2_4
XFILLER_116_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7258_ _7277_/A _7277_/B _7250_/Y vssd1 vssd1 vccd1 vccd1 _7263_/B sky130_fd_sc_hd__o21ai_4
XFILLER_89_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6209_ _6262_/S _6206_/X _6207_/X _6193_/A vssd1 vssd1 vccd1 vccd1 _6209_/X sky130_fd_sc_hd__o211a_1
XFILLER_58_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7189_ _7203_/A _7203_/B _7180_/X vssd1 vssd1 vccd1 vccd1 _7190_/B sky130_fd_sc_hd__o21bai_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _8065_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4890_ _4890_/A _4919_/C vssd1 vssd1 vccd1 vccd1 _4892_/A sky130_fd_sc_hd__xnor2_4
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6560_ _6626_/B _6560_/B vssd1 vssd1 vccd1 vccd1 _6617_/A sky130_fd_sc_hd__nor2_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5511_ _5858_/B _6951_/D _5541_/A _5880_/A vssd1 vssd1 vccd1 vccd1 _5511_/X sky130_fd_sc_hd__o2bb2a_2
XFILLER_118_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6491_ _6584_/A _6583_/B vssd1 vssd1 vccd1 vccd1 _6571_/B sky130_fd_sc_hd__nand2_4
X_5442_ _5443_/A _5443_/B vssd1 vssd1 vccd1 vccd1 _5442_/Y sky130_fd_sc_hd__nor2_1
X_5373_ _7026_/A _5373_/B vssd1 vssd1 vccd1 vccd1 _5375_/A sky130_fd_sc_hd__xor2_4
XFILLER_99_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4324_ _4341_/A1 _4315_/B _4547_/D _4356_/A vssd1 vssd1 vccd1 vccd1 _4324_/X sky130_fd_sc_hd__a31o_1
X_7112_ _7112_/A _7112_/B vssd1 vssd1 vccd1 vccd1 _7119_/A sky130_fd_sc_hd__xnor2_1
XFILLER_101_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout128 _5993_/B vssd1 vssd1 vccd1 vccd1 _5134_/A2 sky130_fd_sc_hd__buf_4
Xfanout106 _7358_/B vssd1 vssd1 vccd1 vccd1 _7210_/B sky130_fd_sc_hd__buf_12
X_7043_ _7041_/A _7041_/B _7042_/X vssd1 vssd1 vccd1 vccd1 _7045_/B sky130_fd_sc_hd__o21ba_1
Xfanout117 _4920_/A vssd1 vssd1 vccd1 vccd1 _4585_/B sky130_fd_sc_hd__buf_4
X_4255_ _4341_/A1 _4322_/B _4322_/C _4248_/X vssd1 vssd1 vccd1 vccd1 _4406_/A sky130_fd_sc_hd__a31o_4
Xfanout139 _4343_/Y vssd1 vssd1 vccd1 vccd1 _7319_/A sky130_fd_sc_hd__buf_12
XFILLER_101_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4186_ _4187_/B vssd1 vssd1 vccd1 vccd1 _6274_/B sky130_fd_sc_hd__inv_2
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7945_ _7943_/X _7944_/Y _7856_/A vssd1 vssd1 vccd1 vccd1 _8042_/D sky130_fd_sc_hd__a21oi_1
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7876_ _7837_/A _7873_/Y _7874_/X _7918_/B vssd1 vssd1 vccd1 vccd1 _7876_/X sky130_fd_sc_hd__a31o_1
XFILLER_70_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6827_ _7558_/A _6827_/B _7392_/A vssd1 vssd1 vccd1 vccd1 _7392_/B sky130_fd_sc_hd__nor3_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6758_ _6732_/X _6757_/X _7894_/A vssd1 vssd1 vccd1 vccd1 _6760_/B sky130_fd_sc_hd__o21a_1
XFILLER_10_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6689_ _6688_/X _6677_/A _6689_/S vssd1 vssd1 vccd1 vccd1 _6689_/X sky130_fd_sc_hd__mux2_1
X_5709_ _5941_/B _5709_/B vssd1 vssd1 vccd1 vccd1 _5942_/A sky130_fd_sc_hd__and2b_1
XFILLER_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4040_ _8057_/Q _8056_/Q _8055_/Q _4096_/B vssd1 vssd1 vccd1 vccd1 _4052_/B sky130_fd_sc_hd__or4_2
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5991_ _6289_/A _4119_/Y _6272_/A _4071_/B vssd1 vssd1 vccd1 vccd1 _5995_/A sky130_fd_sc_hd__a211o_1
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7730_ _6255_/D _7729_/X _7930_/A vssd1 vssd1 vccd1 vccd1 _7731_/B sky130_fd_sc_hd__mux2_1
X_4942_ _4942_/A _4942_/B vssd1 vssd1 vccd1 vccd1 _4976_/B sky130_fd_sc_hd__xor2_4
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7661_ _7837_/A _7684_/A _7684_/B vssd1 vssd1 vccd1 vccd1 _7663_/A sky130_fd_sc_hd__a21oi_1
X_6612_ _6612_/A _6612_/B vssd1 vssd1 vccd1 vccd1 _6616_/B sky130_fd_sc_hd__nor2_1
XFILLER_60_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4873_ _4897_/A _4873_/B vssd1 vssd1 vccd1 vccd1 _4878_/A sky130_fd_sc_hd__xnor2_4
X_7592_ _7657_/B _7592_/B vssd1 vssd1 vccd1 vccd1 _7592_/Y sky130_fd_sc_hd__nand2_1
X_6543_ _6543_/A _6543_/B vssd1 vssd1 vccd1 vccd1 _6547_/A sky130_fd_sc_hd__xor2_4
X_6474_ _6406_/X _6474_/B vssd1 vssd1 vccd1 vccd1 _6529_/A sky130_fd_sc_hd__nand2b_4
XFILLER_118_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5425_ _5395_/A _5393_/Y _5392_/Y vssd1 vssd1 vccd1 vccd1 _5556_/A sky130_fd_sc_hd__a21o_1
XFILLER_102_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5356_ _5356_/A _5356_/B vssd1 vssd1 vccd1 vccd1 _5357_/B sky130_fd_sc_hd__xnor2_4
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8075_ _8075_/CLK _8075_/D vssd1 vssd1 vccd1 vccd1 _8075_/Q sky130_fd_sc_hd__dfxtp_4
X_4307_ _5145_/B _5145_/C _5268_/A vssd1 vssd1 vccd1 vccd1 _5322_/B sky130_fd_sc_hd__a21o_2
X_5287_ _5287_/A _5287_/B vssd1 vssd1 vccd1 vccd1 _5288_/B sky130_fd_sc_hd__or2_1
X_4238_ _4178_/X _4260_/C _4235_/X _4315_/B vssd1 vssd1 vccd1 vccd1 _4239_/C sky130_fd_sc_hd__a211o_1
XFILLER_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7026_ _7026_/A _7086_/A vssd1 vssd1 vccd1 vccd1 _7027_/C sky130_fd_sc_hd__xor2_2
XFILLER_101_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4169_ _8076_/Q _4170_/B vssd1 vssd1 vccd1 vccd1 _4169_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7928_ _7928_/A _7928_/B vssd1 vssd1 vccd1 vccd1 _8041_/D sky130_fd_sc_hd__nor2_1
XFILLER_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7859_ _7883_/A _7883_/B vssd1 vssd1 vccd1 vccd1 _7886_/C sky130_fd_sc_hd__xnor2_1
XFILLER_23_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5210_ _5208_/A _5465_/A _5166_/B vssd1 vssd1 vccd1 vccd1 _5210_/X sky130_fd_sc_hd__a21o_1
X_6190_ _6199_/S _6149_/X _6189_/X vssd1 vssd1 vccd1 vccd1 _6190_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5141_ _5207_/A _6778_/B vssd1 vssd1 vccd1 vccd1 _6780_/A sky130_fd_sc_hd__or2_1
X_5072_ _5071_/A _5071_/B _5184_/A vssd1 vssd1 vccd1 vccd1 _5074_/C sky130_fd_sc_hd__a21o_2
XFILLER_96_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4023_ _8012_/Q _8013_/Q _7955_/S vssd1 vssd1 vccd1 vccd1 _8013_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7713_ _7749_/A _7713_/B vssd1 vssd1 vccd1 vccd1 _7744_/B sky130_fd_sc_hd__nor2_1
X_5974_ _4059_/B _4303_/C _4135_/X _6021_/A0 vssd1 vssd1 vccd1 vccd1 _5974_/X sky130_fd_sc_hd__o211a_1
XFILLER_52_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4925_ _4931_/B _4925_/B _4925_/C vssd1 vssd1 vccd1 vccd1 _4963_/A sky130_fd_sc_hd__and3_2
X_7644_ _7757_/D _7702_/A vssd1 vssd1 vccd1 vccd1 _7644_/Y sky130_fd_sc_hd__xnor2_4
X_4856_ _4850_/A _4947_/C _4748_/B vssd1 vssd1 vccd1 vccd1 _4865_/A sky130_fd_sc_hd__a21o_2
XFILLER_33_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7575_ _7611_/D _7611_/C _7611_/B vssd1 vssd1 vccd1 vccd1 _7643_/A sky130_fd_sc_hd__nand3_4
X_6526_ _6463_/X _6506_/X _6544_/S vssd1 vssd1 vccd1 vccd1 _6527_/B sky130_fd_sc_hd__mux2_4
X_4787_ _4787_/A vssd1 vssd1 vccd1 vccd1 _5063_/A sky130_fd_sc_hd__inv_2
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6457_ _6482_/B _6482_/A vssd1 vssd1 vccd1 vccd1 _6457_/X sky130_fd_sc_hd__and2b_1
X_6388_ _5842_/B _7123_/A _6456_/S vssd1 vssd1 vccd1 vccd1 _6388_/X sky130_fd_sc_hd__mux2_1
X_5408_ _5408_/A _5408_/B vssd1 vssd1 vccd1 vccd1 _5410_/B sky130_fd_sc_hd__xor2_4
XFILLER_114_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5339_ _5621_/A _5516_/A _5338_/Y vssd1 vssd1 vccd1 vccd1 _5339_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_102_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8058_ _8075_/CLK _8058_/D vssd1 vssd1 vccd1 vccd1 _8058_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_75_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7009_ _7213_/B _7195_/B vssd1 vssd1 vccd1 vccd1 _7122_/A sky130_fd_sc_hd__nand2_2
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4710_ _4709_/B _4708_/A _4708_/B vssd1 vssd1 vccd1 vccd1 _4710_/Y sky130_fd_sc_hd__o21bai_2
X_5690_ _5715_/A _5796_/B vssd1 vssd1 vccd1 vccd1 _5736_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4641_ _4641_/A _4641_/B vssd1 vssd1 vccd1 vccd1 _4644_/A sky130_fd_sc_hd__nand2_4
XFILLER_30_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7360_ _7363_/A _7363_/B vssd1 vssd1 vccd1 vccd1 _7364_/A sky130_fd_sc_hd__nor2_1
X_4572_ _4654_/A _4572_/B vssd1 vssd1 vccd1 vccd1 _4574_/C sky130_fd_sc_hd__xnor2_4
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout8 _6134_/X vssd1 vssd1 vccd1 vccd1 _6166_/S sky130_fd_sc_hd__clkbuf_4
X_6311_ _6311_/A _6766_/S vssd1 vssd1 vccd1 vccd1 _6311_/Y sky130_fd_sc_hd__nor2_1
X_7291_ _7301_/A _7301_/B _7288_/Y vssd1 vssd1 vccd1 vccd1 _7300_/B sky130_fd_sc_hd__a21o_2
X_6242_ _6240_/Y _6241_/Y _6242_/S vssd1 vssd1 vccd1 vccd1 _6242_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6173_ _6173_/A _6173_/B vssd1 vssd1 vccd1 vccd1 _6174_/B sky130_fd_sc_hd__xor2_1
XFILLER_111_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5124_ _5621_/A _5386_/A vssd1 vssd1 vccd1 vccd1 _5166_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5055_ _4913_/Y _4944_/X _4915_/B vssd1 vssd1 vccd1 vccd1 _5247_/C sky130_fd_sc_hd__a21o_2
XFILLER_38_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4006_ _8067_/Q vssd1 vssd1 vccd1 vccd1 _4315_/A sky130_fd_sc_hd__inv_2
XFILLER_65_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5957_ _5957_/A _5957_/B vssd1 vssd1 vccd1 vccd1 _5959_/C sky130_fd_sc_hd__xor2_1
X_4908_ _5090_/A _4878_/A _4900_/A _4901_/Y vssd1 vssd1 vccd1 vccd1 _4916_/A sky130_fd_sc_hd__o31ai_4
XFILLER_40_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7627_ _7847_/A _7544_/C _7626_/X vssd1 vssd1 vccd1 vccd1 _7629_/B sky130_fd_sc_hd__o21ai_4
X_5888_ _5904_/A _5888_/B vssd1 vssd1 vccd1 vccd1 _5902_/A sky130_fd_sc_hd__xor2_4
X_4839_ _4654_/A _7001_/A _5013_/B vssd1 vssd1 vccd1 vccd1 _4839_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7558_ _7558_/A _8010_/Q _8009_/Q vssd1 vssd1 vccd1 vccd1 _7558_/X sky130_fd_sc_hd__or3b_2
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6509_ _6387_/A _6387_/B _6508_/X vssd1 vssd1 vccd1 vccd1 _6509_/X sky130_fd_sc_hd__o21a_1
X_7489_ _7487_/Y _7488_/X _7513_/S vssd1 vssd1 vccd1 vccd1 _7489_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_6 _7085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6860_ _6861_/A _6861_/B vssd1 vssd1 vccd1 vccd1 _6860_/Y sky130_fd_sc_hd__nand2_2
X_6791_ _6791_/A _6791_/B vssd1 vssd1 vccd1 vccd1 _6812_/A sky130_fd_sc_hd__nor2_2
XFILLER_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5811_ _5811_/A _5811_/B vssd1 vssd1 vccd1 vccd1 _5817_/B sky130_fd_sc_hd__xor2_4
X_5742_ _5741_/A _5741_/B _5779_/B _5779_/A vssd1 vssd1 vccd1 vccd1 _5746_/A sky130_fd_sc_hd__a22o_4
XFILLER_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5673_ _5722_/A _5722_/B _7285_/B vssd1 vssd1 vccd1 vccd1 _5676_/B sky130_fd_sc_hd__nand3_4
X_7412_ _7419_/A _7438_/A vssd1 vssd1 vccd1 vccd1 _7436_/A sky130_fd_sc_hd__nor2_2
X_4624_ _4620_/A _4619_/C _4619_/B vssd1 vssd1 vccd1 vccd1 _4625_/C sky130_fd_sc_hd__a21o_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7343_ _7345_/A _7345_/B vssd1 vssd1 vccd1 vccd1 _7343_/X sky130_fd_sc_hd__and2b_1
X_4555_ _4555_/A _4556_/A _4555_/C vssd1 vssd1 vccd1 vccd1 _4555_/X sky130_fd_sc_hd__and3_1
XFILLER_104_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7274_ _7274_/A _7274_/B vssd1 vssd1 vccd1 vccd1 _7297_/A sky130_fd_sc_hd__xnor2_4
X_4486_ _5969_/B _4482_/Y _4602_/A vssd1 vssd1 vccd1 vccd1 _4486_/X sky130_fd_sc_hd__o21a_1
X_6225_ _6220_/Y _6250_/B _6225_/S vssd1 vssd1 vccd1 vccd1 _6225_/X sky130_fd_sc_hd__mux2_1
X_6156_ _6156_/A _6160_/B vssd1 vssd1 vccd1 vccd1 _6156_/Y sky130_fd_sc_hd__nand2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5107_ _8065_/Q _5107_/B _5107_/C vssd1 vssd1 vccd1 vccd1 _5107_/X sky130_fd_sc_hd__or3_4
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6087_ _6110_/A _6093_/B vssd1 vssd1 vccd1 vccd1 _6132_/A sky130_fd_sc_hd__nor2_2
XFILLER_57_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5038_ _5038_/A _5038_/B vssd1 vssd1 vccd1 vccd1 _5039_/B sky130_fd_sc_hd__xor2_1
XFILLER_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6989_ _6992_/A _6990_/B vssd1 vssd1 vccd1 vccd1 _6989_/X sky130_fd_sc_hd__and2b_1
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4340_ _4340_/A _4340_/B vssd1 vssd1 vccd1 vccd1 _4340_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4271_ _4241_/B _4227_/X _4231_/X _4178_/X vssd1 vssd1 vccd1 vccd1 _4271_/X sky130_fd_sc_hd__o211a_1
X_6010_ _6349_/B _6010_/B vssd1 vssd1 vccd1 vccd1 _6012_/A sky130_fd_sc_hd__xor2_4
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7961_ _7961_/A _7961_/B vssd1 vssd1 vccd1 vccd1 _7971_/B sky130_fd_sc_hd__nor2_1
XFILLER_94_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7892_ _7939_/A _7877_/B _7891_/Y vssd1 vssd1 vccd1 vccd1 _7892_/Y sky130_fd_sc_hd__a21oi_1
X_6912_ _6912_/A _6913_/A _6912_/C vssd1 vssd1 vccd1 vccd1 _6912_/X sky130_fd_sc_hd__or3_1
XFILLER_62_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6843_ _6843_/A _6870_/A vssd1 vssd1 vccd1 vccd1 _6845_/B sky130_fd_sc_hd__nand2_2
XFILLER_35_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6774_ _8010_/Q _8009_/Q _6774_/C vssd1 vssd1 vccd1 vccd1 _6774_/X sky130_fd_sc_hd__or3_4
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5725_ _5763_/A _5763_/B _5719_/X vssd1 vssd1 vccd1 vccd1 _5728_/A sky130_fd_sc_hd__a21o_2
XFILLER_22_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5656_ _5652_/A _5651_/Y _5653_/Y vssd1 vssd1 vccd1 vccd1 _5662_/A sky130_fd_sc_hd__o21ai_4
XFILLER_108_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4607_ _4574_/A _4574_/B _4574_/C vssd1 vssd1 vccd1 vccd1 _4607_/Y sky130_fd_sc_hd__o21ai_4
X_5587_ _5588_/A _5588_/B vssd1 vssd1 vccd1 vccd1 _5587_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7326_ _7326_/A _7326_/B vssd1 vssd1 vccd1 vccd1 _7348_/A sky130_fd_sc_hd__xnor2_2
X_4538_ _4506_/A _4506_/B _4510_/Y vssd1 vssd1 vccd1 vccd1 _4539_/B sky130_fd_sc_hd__a21oi_4
XFILLER_2_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7257_ _7257_/A _7257_/B vssd1 vssd1 vccd1 vccd1 _7277_/B sky130_fd_sc_hd__xnor2_4
X_4469_ _4394_/Y _4566_/A _4467_/X _4468_/Y vssd1 vssd1 vccd1 vccd1 _4497_/A sky130_fd_sc_hd__a211oi_4
XFILLER_104_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6208_ _6262_/S _6206_/X _6207_/X vssd1 vssd1 vccd1 vccd1 _6208_/X sky130_fd_sc_hd__o21a_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7188_ _7188_/A _7227_/A vssd1 vssd1 vccd1 vccd1 _7203_/B sky130_fd_sc_hd__xnor2_4
XFILLER_112_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6139_ _7085_/B _6139_/B vssd1 vssd1 vccd1 vccd1 _6139_/Y sky130_fd_sc_hd__nor2_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5510_ _5715_/A _5755_/A vssd1 vssd1 vccd1 vccd1 _5563_/A sky130_fd_sc_hd__nor2_2
X_6490_ _6485_/B _6488_/Y _6443_/A _6425_/B vssd1 vssd1 vccd1 vccd1 _6583_/B sky130_fd_sc_hd__o2bb2a_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5441_ _5441_/A _5441_/B vssd1 vssd1 vccd1 vccd1 _5443_/B sky130_fd_sc_hd__xnor2_4
X_5372_ _5123_/A _5123_/B _7285_/B vssd1 vssd1 vccd1 vccd1 _5373_/B sky130_fd_sc_hd__o21a_4
XFILLER_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4323_ _4341_/A1 _4239_/B _4239_/C _4548_/C vssd1 vssd1 vccd1 vccd1 _4323_/X sky130_fd_sc_hd__a31o_2
X_7111_ _7111_/A _7111_/B vssd1 vssd1 vccd1 vccd1 _7135_/A sky130_fd_sc_hd__xnor2_4
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout129 _4121_/X vssd1 vssd1 vccd1 vccd1 _5993_/B sky130_fd_sc_hd__buf_4
X_7042_ _7052_/B _7052_/A vssd1 vssd1 vccd1 vccd1 _7042_/X sky130_fd_sc_hd__and2b_1
Xfanout107 _7358_/B vssd1 vssd1 vccd1 vccd1 _5855_/A sky130_fd_sc_hd__buf_6
Xfanout118 _4367_/X vssd1 vssd1 vccd1 vccd1 _4920_/A sky130_fd_sc_hd__buf_4
XFILLER_113_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4254_ _4341_/A1 _4322_/B _4322_/C _4248_/X vssd1 vssd1 vccd1 vccd1 _4376_/A sky130_fd_sc_hd__a31oi_4
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4185_ _8073_/Q _4185_/B vssd1 vssd1 vccd1 vccd1 _4187_/B sky130_fd_sc_hd__xor2_4
XFILLER_79_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7944_ _8042_/Q _7944_/B vssd1 vssd1 vccd1 vccd1 _7944_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7875_ _7939_/A _7874_/X _7873_/Y vssd1 vssd1 vccd1 vccd1 _7877_/B sky130_fd_sc_hd__a21o_1
X_6826_ _7558_/A _7392_/A _6827_/B vssd1 vssd1 vccd1 vccd1 _6828_/B sky130_fd_sc_hd__o21a_1
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6757_ _6757_/A _6757_/B _6757_/C _6757_/D vssd1 vssd1 vccd1 vccd1 _6757_/X sky130_fd_sc_hd__or4_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5708_ _5708_/A _5708_/B vssd1 vssd1 vccd1 vccd1 _5941_/B sky130_fd_sc_hd__xor2_1
X_6688_ _6524_/A _6539_/A _6688_/S vssd1 vssd1 vccd1 vccd1 _6688_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5639_ _5639_/A _5639_/B vssd1 vssd1 vccd1 vccd1 _5641_/B sky130_fd_sc_hd__xnor2_4
X_7309_ _7332_/A _7310_/B vssd1 vssd1 vccd1 vccd1 _7309_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5990_ _6326_/B _5990_/B vssd1 vssd1 vccd1 vccd1 _5996_/A sky130_fd_sc_hd__xnor2_2
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4941_ _4998_/A _5040_/B _4933_/A _4934_/X vssd1 vssd1 vccd1 vccd1 _4976_/A sky130_fd_sc_hd__a31o_4
X_7660_ _7687_/A _7687_/B vssd1 vssd1 vccd1 vccd1 _7684_/B sky130_fd_sc_hd__xor2_2
X_4872_ _4879_/A _4879_/B vssd1 vssd1 vccd1 vccd1 _4872_/Y sky130_fd_sc_hd__nor2_1
X_6611_ _6611_/A _6611_/B vssd1 vssd1 vccd1 vccd1 _6612_/B sky130_fd_sc_hd__and2_1
XFILLER_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7591_ _7657_/A _7549_/Y _7624_/S vssd1 vssd1 vccd1 vccd1 _7592_/B sky130_fd_sc_hd__mux2_1
X_6542_ _6544_/S _6502_/Y _6541_/Y vssd1 vssd1 vccd1 vccd1 _6543_/B sky130_fd_sc_hd__a21oi_4
X_6473_ _6443_/A _6404_/B _6407_/B vssd1 vssd1 vccd1 vccd1 _6473_/Y sky130_fd_sc_hd__a21oi_1
X_5424_ _5426_/A _5426_/B vssd1 vssd1 vccd1 vccd1 _5612_/A sky130_fd_sc_hd__or2_1
X_5355_ _5356_/A _5356_/B vssd1 vssd1 vccd1 vccd1 _5355_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_102_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8074_ _8075_/CLK _8074_/D vssd1 vssd1 vccd1 vccd1 _8074_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4306_ _4087_/B _4303_/C _4304_/X _5135_/C1 vssd1 vssd1 vccd1 vccd1 _5145_/C sky130_fd_sc_hd__o211ai_4
X_5286_ _5287_/A _5287_/B vssd1 vssd1 vccd1 vccd1 _5288_/A sky130_fd_sc_hd__nand2_1
X_4237_ _4170_/X _4260_/C _4236_/X _4548_/B vssd1 vssd1 vccd1 vccd1 _4239_/B sky130_fd_sc_hd__a211o_1
X_7025_ _7025_/A _7366_/B vssd1 vssd1 vccd1 vccd1 _7025_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4168_ _8075_/Q _4147_/A _4147_/B _4168_/B1 vssd1 vssd1 vccd1 vccd1 _4170_/B sky130_fd_sc_hd__o31a_4
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4099_ _4088_/A _8053_/Q _8052_/Q _4096_/A vssd1 vssd1 vccd1 vccd1 _4100_/B sky130_fd_sc_hd__o31a_2
XFILLER_83_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7927_ _7991_/D _7925_/X _7926_/X vssd1 vssd1 vccd1 vccd1 _7928_/B sky130_fd_sc_hd__o21ba_1
X_7858_ _7930_/A _7858_/B vssd1 vssd1 vccd1 vccd1 _7883_/B sky130_fd_sc_hd__or2_2
X_6809_ _6809_/A _6809_/B vssd1 vssd1 vccd1 vccd1 _6810_/B sky130_fd_sc_hd__or2_1
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7789_ _7789_/A _7789_/B _7789_/C vssd1 vssd1 vccd1 vccd1 _7822_/A sky130_fd_sc_hd__and3_2
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5140_ _5207_/A _6842_/B vssd1 vssd1 vccd1 vccd1 _5208_/A sky130_fd_sc_hd__nor2_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5071_ _5071_/A _5071_/B vssd1 vssd1 vccd1 vccd1 _5184_/B sky130_fd_sc_hd__nand2_2
X_4022_ _8011_/Q _8012_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _8012_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5973_ _5133_/A _5133_/B _5087_/B vssd1 vssd1 vccd1 vccd1 _5973_/Y sky130_fd_sc_hd__a21oi_4
X_7712_ _7748_/A _7748_/B vssd1 vssd1 vccd1 vccd1 _7713_/B sky130_fd_sc_hd__and2_1
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4924_ _4798_/X _4927_/A _4923_/X vssd1 vssd1 vccd1 vccd1 _4925_/C sky130_fd_sc_hd__a21o_1
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7643_ _7643_/A _7643_/B _7702_/A vssd1 vssd1 vccd1 vccd1 _7671_/A sky130_fd_sc_hd__or3_4
X_4855_ _4857_/A _4867_/A _4857_/C vssd1 vssd1 vccd1 vccd1 _4860_/B sky130_fd_sc_hd__a21oi_4
X_7574_ _7831_/A _6255_/B _7573_/X vssd1 vssd1 vccd1 vccd1 _7611_/B sky130_fd_sc_hd__a21boi_4
X_4786_ _4786_/A _4786_/B vssd1 vssd1 vccd1 vccd1 _4787_/A sky130_fd_sc_hd__nand2_1
X_6525_ _6525_/A _6525_/B vssd1 vssd1 vccd1 vccd1 _6562_/A sky130_fd_sc_hd__or2_2
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6456_ _7366_/A _7366_/B _6456_/S vssd1 vssd1 vccd1 vccd1 _6482_/B sky130_fd_sc_hd__mux2_2
X_6387_ _6387_/A _6387_/B vssd1 vssd1 vccd1 vccd1 _6520_/A sky130_fd_sc_hd__xnor2_4
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5407_ _5407_/A _5407_/B vssd1 vssd1 vccd1 vccd1 _5408_/B sky130_fd_sc_hd__xor2_4
XFILLER_88_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5338_ _5782_/A _5338_/B vssd1 vssd1 vccd1 vccd1 _5338_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8057_ _8057_/CLK _8057_/D vssd1 vssd1 vccd1 vccd1 _8057_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5269_ _5977_/B _5083_/X _5084_/X _5268_/X vssd1 vssd1 vccd1 vccd1 _5271_/B sky130_fd_sc_hd__a31oi_4
X_7008_ _7008_/A _7008_/B vssd1 vssd1 vccd1 vccd1 _7015_/A sky130_fd_sc_hd__xnor2_4
XFILLER_47_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4640_ _4639_/B _4639_/C _4639_/A vssd1 vssd1 vccd1 vccd1 _4650_/A sky130_fd_sc_hd__a21bo_1
X_6310_ _6310_/A _6310_/B vssd1 vssd1 vccd1 vccd1 _7401_/A sky130_fd_sc_hd__xnor2_4
X_4571_ _4654_/A _4572_/B vssd1 vssd1 vccd1 vccd1 _4571_/Y sky130_fd_sc_hd__nor2_2
XFILLER_116_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout9 _6113_/X vssd1 vssd1 vccd1 vccd1 _6199_/S sky130_fd_sc_hd__buf_4
X_7290_ _7290_/A _7290_/B vssd1 vssd1 vccd1 vccd1 _7301_/B sky130_fd_sc_hd__xor2_4
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6241_ _6241_/A _6241_/B vssd1 vssd1 vccd1 vccd1 _6241_/Y sky130_fd_sc_hd__xnor2_1
X_6172_ _6172_/A _6172_/B vssd1 vssd1 vccd1 vccd1 _6172_/X sky130_fd_sc_hd__xor2_2
XFILLER_97_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5123_ _5123_/A _5123_/B vssd1 vssd1 vccd1 vccd1 _5273_/A sky130_fd_sc_hd__nor2_4
XFILLER_97_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _5290_/A _5054_/B _5054_/C _5054_/D vssd1 vssd1 vccd1 vccd1 _5247_/B sky130_fd_sc_hd__or4_4
X_4005_ _6188_/A vssd1 vssd1 vccd1 vccd1 _4005_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5956_ _5956_/A _6354_/A vssd1 vssd1 vccd1 vccd1 _5957_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4907_ _4909_/B _4909_/A vssd1 vssd1 vccd1 vccd1 _4914_/A sky130_fd_sc_hd__nand2b_1
XFILLER_21_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5887_ _5904_/A _5888_/B vssd1 vssd1 vccd1 vccd1 _5887_/Y sky130_fd_sc_hd__nor2_1
X_7626_ _7766_/B _7847_/B vssd1 vssd1 vccd1 vccd1 _7626_/X sky130_fd_sc_hd__or2_2
X_4838_ _4720_/X _4721_/Y _4726_/Y _4720_/C _4837_/X vssd1 vssd1 vccd1 vccd1 _4838_/X
+ sky130_fd_sc_hd__o221a_1
X_7557_ _7939_/A _7590_/A _7590_/B vssd1 vssd1 vccd1 vccd1 _7557_/Y sky130_fd_sc_hd__a21oi_1
X_4769_ _4991_/A _5090_/B _4868_/B _4868_/C vssd1 vssd1 vccd1 vccd1 _4775_/B sky130_fd_sc_hd__a22o_2
XFILLER_119_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6508_ _6387_/A _6387_/B _6399_/A _6506_/X _6398_/A vssd1 vssd1 vccd1 vccd1 _6508_/X
+ sky130_fd_sc_hd__a221o_1
X_7488_ _7488_/A _7488_/B vssd1 vssd1 vccd1 vccd1 _7488_/X sky130_fd_sc_hd__xor2_2
X_6439_ _6430_/X _6438_/X _6483_/A vssd1 vssd1 vccd1 vccd1 _6439_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_7 _6951_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6790_ _6806_/A _7027_/A vssd1 vssd1 vccd1 vccd1 _6795_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5810_ _6878_/B _5927_/B vssd1 vssd1 vccd1 vccd1 _5817_/A sky130_fd_sc_hd__nand2_2
X_5741_ _5741_/A _5741_/B vssd1 vssd1 vccd1 vccd1 _5779_/B sky130_fd_sc_hd__xor2_4
XFILLER_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7411_ _7411_/A _7766_/A vssd1 vssd1 vccd1 vccd1 _7438_/A sky130_fd_sc_hd__xnor2_4
X_5672_ _5672_/A _5925_/A vssd1 vssd1 vccd1 vccd1 _5677_/A sky130_fd_sc_hd__nor2_2
XFILLER_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4623_ _4654_/A _4989_/A vssd1 vssd1 vccd1 vccd1 _4625_/B sky130_fd_sc_hd__nor2_1
X_7342_ _7350_/A _7350_/B vssd1 vssd1 vccd1 vccd1 _7345_/B sky130_fd_sc_hd__and2b_2
X_4554_ _4555_/A _4555_/C vssd1 vssd1 vccd1 vccd1 _4556_/B sky130_fd_sc_hd__nand2_2
X_7273_ _7273_/A _7273_/B vssd1 vssd1 vccd1 vccd1 _7471_/A sky130_fd_sc_hd__nand2_4
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6224_ _6130_/Y _6153_/Y _6254_/S vssd1 vssd1 vccd1 vccd1 _6250_/B sky130_fd_sc_hd__mux2_1
X_4485_ _4406_/A _4441_/A _4472_/B _4472_/A vssd1 vssd1 vccd1 vccd1 _4485_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6155_ _6155_/A _6155_/B vssd1 vssd1 vccd1 vccd1 _6160_/B sky130_fd_sc_hd__xnor2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _8065_/Q _5107_/B _5107_/C vssd1 vssd1 vccd1 vccd1 _5106_/Y sky130_fd_sc_hd__nor3_2
XFILLER_97_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6086_ _6086_/A _6086_/B vssd1 vssd1 vccd1 vccd1 _6093_/B sky130_fd_sc_hd__xnor2_4
XFILLER_85_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5037_ _5038_/A _5038_/B vssd1 vssd1 vccd1 vccd1 _5037_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6988_ _6988_/A _6988_/B vssd1 vssd1 vccd1 vccd1 _6990_/B sky130_fd_sc_hd__and2_1
XFILLER_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5939_ _6205_/A _6205_/B _6137_/A _5785_/X vssd1 vssd1 vccd1 vccd1 _6135_/A sky130_fd_sc_hd__a31oi_4
XFILLER_21_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7609_ _6222_/Y _7608_/Y _7639_/B vssd1 vssd1 vccd1 vccd1 _7831_/B sky130_fd_sc_hd__mux2_1
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4270_ _4241_/B _4227_/X _4231_/X _4192_/B vssd1 vssd1 vccd1 vccd1 _4270_/X sky130_fd_sc_hd__o211a_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7960_ _7961_/B _7960_/B vssd1 vssd1 vccd1 vccd1 _8045_/D sky130_fd_sc_hd__nor2_1
XFILLER_82_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7891_ _7657_/A _7889_/A _7913_/A _7913_/B _7914_/A vssd1 vssd1 vccd1 vccd1 _7891_/Y
+ sky130_fd_sc_hd__a221oi_4
X_6911_ _6912_/A _6912_/C vssd1 vssd1 vccd1 vccd1 _6913_/B sky130_fd_sc_hd__nor2_1
X_6842_ _7027_/A _6842_/B _6842_/C vssd1 vssd1 vccd1 vccd1 _6870_/A sky130_fd_sc_hd__or3_2
X_6773_ _8010_/Q _8009_/Q _6774_/C vssd1 vssd1 vccd1 vccd1 _7923_/A sky130_fd_sc_hd__nor3_4
XFILLER_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5724_ _5724_/A _5724_/B vssd1 vssd1 vccd1 vccd1 _5763_/B sky130_fd_sc_hd__xnor2_4
XFILLER_109_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5655_ _5697_/A _5697_/B _5644_/X vssd1 vssd1 vccd1 vccd1 _5657_/B sky130_fd_sc_hd__a21oi_4
X_4606_ _4606_/A _4606_/B _4606_/C vssd1 vssd1 vccd1 vccd1 _4606_/Y sky130_fd_sc_hd__nor3_4
X_7325_ _7323_/Y _7325_/B vssd1 vssd1 vccd1 vccd1 _7487_/A sky130_fd_sc_hd__nand2b_1
X_5586_ _5588_/A _5588_/B vssd1 vssd1 vccd1 vccd1 _5586_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4537_ _4537_/A _4537_/B vssd1 vssd1 vccd1 vccd1 _4540_/A sky130_fd_sc_hd__xnor2_4
XFILLER_89_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7256_ _7256_/A _7256_/B vssd1 vssd1 vccd1 vccd1 _7277_/A sky130_fd_sc_hd__xnor2_4
X_4468_ _4516_/B _4467_/C _4467_/A vssd1 vssd1 vccd1 vccd1 _4468_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6207_ _6081_/Y _6111_/B _6111_/C _6138_/Y vssd1 vssd1 vccd1 vccd1 _6207_/X sky130_fd_sc_hd__a31o_1
X_7187_ _7187_/A _7262_/A vssd1 vssd1 vccd1 vccd1 _7227_/A sky130_fd_sc_hd__nand2_4
XFILLER_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6138_ _6127_/A _6135_/Y _6137_/X _6146_/A vssd1 vssd1 vccd1 vccd1 _6138_/Y sky130_fd_sc_hd__o22ai_2
X_4399_ _4412_/A _4413_/B _4430_/B vssd1 vssd1 vccd1 vccd1 _4399_/Y sky130_fd_sc_hd__a21oi_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _6096_/A _6102_/A vssd1 vssd1 vccd1 vccd1 _6069_/Y sky130_fd_sc_hd__nor2_2
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5440_ _5440_/A _5440_/B vssd1 vssd1 vccd1 vccd1 _5441_/B sky130_fd_sc_hd__xor2_4
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5371_ _5445_/A _5925_/A vssd1 vssd1 vccd1 vccd1 _7026_/A sky130_fd_sc_hd__nor2_8
X_4322_ _4322_/A _4322_/B _4322_/C vssd1 vssd1 vccd1 vccd1 _4322_/X sky130_fd_sc_hd__and3_2
X_7110_ _7110_/A _7110_/B vssd1 vssd1 vccd1 vccd1 _7146_/A sky130_fd_sc_hd__xnor2_4
XFILLER_113_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4253_ _4199_/X _4260_/C _4249_/X _4315_/B vssd1 vssd1 vccd1 vccd1 _4322_/C sky130_fd_sc_hd__a211o_4
Xfanout108 _5323_/X vssd1 vssd1 vccd1 vccd1 _7358_/B sky130_fd_sc_hd__buf_12
X_7041_ _7041_/A _7041_/B vssd1 vssd1 vccd1 vccd1 _7052_/B sky130_fd_sc_hd__xnor2_4
Xfanout119 _4350_/X vssd1 vssd1 vccd1 vccd1 _4998_/A sky130_fd_sc_hd__buf_6
XFILLER_99_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4184_ _4210_/B _4210_/C vssd1 vssd1 vccd1 vccd1 _4184_/Y sky130_fd_sc_hd__nand2_2
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7943_ _7934_/X _7937_/X _7941_/X _7942_/Y _7952_/B1 vssd1 vssd1 vccd1 vccd1 _7943_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7874_ _7874_/A _7874_/B _7874_/C _7874_/D vssd1 vssd1 vccd1 vccd1 _7874_/X sky130_fd_sc_hd__or4_2
XFILLER_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6825_ _6810_/A _6819_/B _6819_/A vssd1 vssd1 vccd1 vccd1 _7392_/A sky130_fd_sc_hd__o21bai_2
X_6756_ _6572_/Y _6737_/B _6755_/X vssd1 vssd1 vccd1 vccd1 _6756_/X sky130_fd_sc_hd__o21ba_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5707_ _5748_/A _5748_/B _5702_/Y vssd1 vssd1 vccd1 vccd1 _5709_/B sky130_fd_sc_hd__a21o_1
X_6687_ _6704_/B _6686_/X _6751_/S vssd1 vssd1 vccd1 vccd1 _6687_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5638_ _5185_/Y _7285_/B _5633_/B _5631_/X vssd1 vssd1 vccd1 vccd1 _5641_/A sky130_fd_sc_hd__a31oi_4
XFILLER_117_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5569_ _5568_/B _5569_/B vssd1 vssd1 vccd1 vccd1 _5570_/B sky130_fd_sc_hd__and2b_1
X_7308_ _7285_/A _7285_/B _7285_/C _7307_/X vssd1 vssd1 vccd1 vccd1 _7310_/B sky130_fd_sc_hd__a31oi_4
XFILLER_77_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7239_ _7239_/A _7239_/B vssd1 vssd1 vccd1 vccd1 _7271_/B sky130_fd_sc_hd__xor2_4
XFILLER_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4940_ _4942_/A _4942_/B vssd1 vssd1 vccd1 vccd1 _4940_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4871_ _4927_/A _4894_/B _4926_/A vssd1 vssd1 vccd1 vccd1 _4879_/B sky130_fd_sc_hd__a21oi_1
X_6610_ _6610_/A _6610_/B vssd1 vssd1 vccd1 vccd1 _6610_/Y sky130_fd_sc_hd__nand2_1
X_7590_ _7590_/A _7590_/B vssd1 vssd1 vccd1 vccd1 _7623_/A sky130_fd_sc_hd__or2_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6541_ _6544_/S _6541_/B vssd1 vssd1 vccd1 vccd1 _6541_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6472_ _6366_/Y _6472_/B vssd1 vssd1 vccd1 vccd1 _6517_/A sky130_fd_sc_hd__and2b_4
X_5423_ _5423_/A _5423_/B vssd1 vssd1 vccd1 vccd1 _5426_/B sky130_fd_sc_hd__xnor2_2
X_5354_ _5354_/A _5354_/B vssd1 vssd1 vccd1 vccd1 _5356_/B sky130_fd_sc_hd__xor2_4
X_4305_ _4074_/Y _4118_/X _4084_/B _4071_/Y vssd1 vssd1 vccd1 vccd1 _4305_/X sky130_fd_sc_hd__o211a_1
XFILLER_101_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8073_ _8080_/CLK _8073_/D vssd1 vssd1 vccd1 vccd1 _8073_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_99_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5285_ _5285_/A _5285_/B vssd1 vssd1 vccd1 vccd1 _5287_/B sky130_fd_sc_hd__and2_1
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4236_ _4241_/B _4227_/X _4231_/X _4180_/Y vssd1 vssd1 vccd1 vccd1 _4236_/X sky130_fd_sc_hd__o211a_1
X_7024_ _7024_/A _7024_/B vssd1 vssd1 vccd1 vccd1 _7031_/A sky130_fd_sc_hd__and2_2
XFILLER_83_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4167_ _4228_/A _4172_/B vssd1 vssd1 vccd1 vccd1 _4167_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4098_ _6326_/A _4098_/B vssd1 vssd1 vccd1 vccd1 _4102_/A sky130_fd_sc_hd__xnor2_2
X_7926_ _8040_/Q _4018_/X _7857_/B _8041_/Q vssd1 vssd1 vccd1 vccd1 _7926_/X sky130_fd_sc_hd__a22o_1
XFILLER_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7857_ _8039_/Q _7857_/B vssd1 vssd1 vccd1 vccd1 _7857_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6808_ _6809_/A _6809_/B vssd1 vssd1 vccd1 vccd1 _6810_/A sky130_fd_sc_hd__nand2_2
XFILLER_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7788_ _7894_/A _7788_/B vssd1 vssd1 vccd1 vccd1 _7789_/C sky130_fd_sc_hd__or2_1
X_6739_ _6738_/Y _6691_/Y _6739_/S vssd1 vssd1 vccd1 vccd1 _6739_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout90 _7124_/A2 vssd1 vssd1 vccd1 vccd1 _5198_/B sky130_fd_sc_hd__buf_2
XFILLER_10_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5070_ _5977_/A _5065_/Y _5066_/Y _5068_/Y vssd1 vssd1 vccd1 vccd1 _5070_/Y sky130_fd_sc_hd__o31ai_4
XFILLER_69_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4021_ input3/X _8011_/Q _7955_/S vssd1 vssd1 vccd1 vccd1 _8011_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5972_ _6349_/A _6177_/A vssd1 vssd1 vccd1 vccd1 _5972_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7711_ _7748_/A _7748_/B vssd1 vssd1 vccd1 vccd1 _7749_/A sky130_fd_sc_hd__nor2_2
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4923_ _5040_/A _4923_/B _4923_/C _4947_/C vssd1 vssd1 vccd1 vccd1 _4923_/X sky130_fd_sc_hd__and4_1
X_7642_ _6255_/A _7641_/Y _7930_/A vssd1 vssd1 vccd1 vccd1 _7702_/A sky130_fd_sc_hd__mux2_8
X_4854_ _4854_/A _4854_/B vssd1 vssd1 vccd1 vccd1 _4857_/C sky130_fd_sc_hd__xnor2_2
XFILLER_20_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7573_ _6225_/S _6216_/X _7572_/X _7831_/A vssd1 vssd1 vccd1 vccd1 _7573_/X sky130_fd_sc_hd__a211o_1
X_4785_ _4785_/A _4785_/B _4789_/A vssd1 vssd1 vccd1 vccd1 _4786_/B sky130_fd_sc_hd__or3_1
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6524_ _6524_/A _6524_/B vssd1 vssd1 vccd1 vccd1 _6525_/B sky130_fd_sc_hd__or2_1
XFILLER_118_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6455_ _6386_/A _6374_/B _6454_/X vssd1 vssd1 vccd1 vccd1 _6482_/A sky130_fd_sc_hd__o21bai_4
X_6386_ _6386_/A _6386_/B _6387_/B vssd1 vssd1 vccd1 vccd1 _6386_/X sky130_fd_sc_hd__and3_1
X_5406_ _5530_/A _6917_/B vssd1 vssd1 vccd1 vccd1 _5408_/A sky130_fd_sc_hd__nor2_4
XFILLER_102_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5337_ _5503_/A _5503_/B _5313_/Y vssd1 vssd1 vccd1 vccd1 _5360_/A sky130_fd_sc_hd__a21oi_4
X_8056_ _8080_/CLK _8056_/D vssd1 vssd1 vccd1 vccd1 _8056_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5268_ _5268_/A _5268_/B vssd1 vssd1 vccd1 vccd1 _5268_/X sky130_fd_sc_hd__and2_2
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4219_ _4209_/X _4217_/Y _4218_/Y _4230_/C vssd1 vssd1 vccd1 vccd1 _4219_/Y sky130_fd_sc_hd__a211oi_4
X_7007_ _7306_/A _7007_/B _7008_/B vssd1 vssd1 vccd1 vccd1 _7007_/X sky130_fd_sc_hd__and3_1
X_5199_ _5530_/A _6778_/B vssd1 vssd1 vccd1 vccd1 _5255_/A sky130_fd_sc_hd__nor2_4
XFILLER_71_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7909_ _7929_/A _7909_/B _7909_/C vssd1 vssd1 vccd1 vccd1 _7910_/D sky130_fd_sc_hd__or3_1
XFILLER_71_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4570_ _4570_/A _4570_/B vssd1 vssd1 vccd1 vccd1 _4572_/B sky130_fd_sc_hd__xor2_4
XFILLER_30_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6240_ _6240_/A _6240_/B vssd1 vssd1 vccd1 vccd1 _6240_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6171_ _6173_/A _6173_/B _5288_/A vssd1 vssd1 vccd1 vccd1 _6172_/B sky130_fd_sc_hd__o21a_1
X_5122_ _5121_/A _5121_/B _5121_/C vssd1 vssd1 vccd1 vccd1 _5123_/B sky130_fd_sc_hd__a21oi_4
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5053_ _5054_/B _5054_/C _5054_/D vssd1 vssd1 vccd1 vccd1 _5364_/A sky130_fd_sc_hd__or3_1
X_4004_ _8045_/Q vssd1 vssd1 vccd1 vccd1 _7956_/B sky130_fd_sc_hd__inv_2
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5955_ _7949_/B _6805_/B vssd1 vssd1 vccd1 vccd1 _7558_/A sky130_fd_sc_hd__or2_4
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4906_ _4906_/A _4906_/B vssd1 vssd1 vccd1 vccd1 _4909_/B sky130_fd_sc_hd__xor2_4
X_5886_ _5886_/A _5886_/B vssd1 vssd1 vccd1 vccd1 _5888_/B sky130_fd_sc_hd__or2_4
X_7625_ _7468_/X _7624_/X _7657_/B vssd1 vssd1 vccd1 vccd1 _7847_/B sky130_fd_sc_hd__mux2_1
X_4837_ _4837_/A _4837_/B vssd1 vssd1 vccd1 vccd1 _4837_/X sky130_fd_sc_hd__and2_1
X_7556_ _7597_/A _7556_/B vssd1 vssd1 vccd1 vccd1 _7590_/B sky130_fd_sc_hd__and2_1
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4768_ _4854_/A _4768_/B vssd1 vssd1 vccd1 vccd1 _4782_/A sky130_fd_sc_hd__xor2_2
X_6507_ _6399_/A _6506_/X _6398_/A vssd1 vssd1 vccd1 vccd1 _6507_/Y sky130_fd_sc_hd__a21oi_1
X_7487_ _7487_/A _7487_/B vssd1 vssd1 vccd1 vccd1 _7487_/Y sky130_fd_sc_hd__xnor2_1
X_4699_ _4652_/A _4652_/C _4652_/B vssd1 vssd1 vccd1 vccd1 _4700_/C sky130_fd_sc_hd__a21bo_1
X_6438_ _5923_/A _7285_/A _6445_/S vssd1 vssd1 vccd1 vccd1 _6438_/X sky130_fd_sc_hd__mux2_2
XFILLER_115_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6369_ _6431_/S _6360_/X _6368_/X vssd1 vssd1 vccd1 vccd1 _6369_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_29_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8039_ _8065_/CLK _8039_/D vssd1 vssd1 vccd1 vccd1 _8039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_8 _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5740_ _5740_/A _5740_/B vssd1 vssd1 vccd1 vccd1 _5741_/B sky130_fd_sc_hd__xor2_4
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7410_ _7766_/A vssd1 vssd1 vccd1 vccd1 _7657_/A sky130_fd_sc_hd__clkinv_2
X_5671_ _5671_/A _5671_/B vssd1 vssd1 vccd1 vccd1 _5726_/A sky130_fd_sc_hd__nor2_4
XFILLER_30_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4622_ _4638_/A _4638_/B vssd1 vssd1 vccd1 vccd1 _4652_/A sky130_fd_sc_hd__and2_1
XFILLER_116_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7341_ _7351_/A _7340_/B _7340_/A vssd1 vssd1 vccd1 vccd1 _7350_/B sky130_fd_sc_hd__a21boi_4
X_4553_ _7319_/A _4551_/B _4386_/D _4387_/A vssd1 vssd1 vccd1 vccd1 _4555_/C sky130_fd_sc_hd__a22o_1
X_4484_ _4475_/X _4483_/X _4436_/A vssd1 vssd1 vccd1 vccd1 _4488_/C sky130_fd_sc_hd__a21o_1
X_7272_ _7271_/B _7272_/B vssd1 vssd1 vccd1 vccd1 _7273_/B sky130_fd_sc_hd__nand2b_2
XFILLER_116_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6223_ _6220_/Y _6222_/Y _6226_/S vssd1 vssd1 vccd1 vccd1 _6255_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6154_ _6148_/A _6147_/B _5948_/Y vssd1 vssd1 vccd1 vccd1 _6155_/B sky130_fd_sc_hd__a21boi_2
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _6086_/A _6086_/B vssd1 vssd1 vccd1 vccd1 _6259_/B sky130_fd_sc_hd__xor2_2
X_5105_ _5367_/A _5244_/A vssd1 vssd1 vccd1 vccd1 _5113_/A sky130_fd_sc_hd__or2_4
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5040_/A _5020_/B _5035_/X _5034_/X vssd1 vssd1 vccd1 vccd1 _5038_/B sky130_fd_sc_hd__a31o_1
XFILLER_38_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6987_ _6987_/A _6987_/B _6987_/C vssd1 vssd1 vccd1 vccd1 _6988_/B sky130_fd_sc_hd__or3_1
XFILLER_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5938_ _5749_/X _5938_/B vssd1 vssd1 vccd1 vccd1 _6137_/A sky130_fd_sc_hd__and2b_4
X_5869_ _5869_/A _5893_/A vssd1 vssd1 vccd1 vccd1 _5871_/B sky130_fd_sc_hd__and2_2
X_7608_ _6078_/A _7570_/B _7570_/Y vssd1 vssd1 vccd1 vccd1 _7608_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_31_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7539_ _7889_/A _7542_/D vssd1 vssd1 vccd1 vccd1 _7539_/X sky130_fd_sc_hd__or2_2
XFILLER_107_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7890_ _7913_/A _7913_/B vssd1 vssd1 vccd1 vccd1 _7914_/A sky130_fd_sc_hd__nor2_4
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6910_ _7030_/A _5621_/A _6877_/Y vssd1 vssd1 vccd1 vccd1 _6912_/C sky130_fd_sc_hd__o21a_1
X_6841_ _6843_/A _6841_/B vssd1 vssd1 vccd1 vccd1 _6842_/C sky130_fd_sc_hd__nand2_1
XFILLER_90_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6772_ _6614_/A _6720_/X _6771_/X vssd1 vssd1 vccd1 vccd1 _6774_/C sky130_fd_sc_hd__o21ai_4
XFILLER_50_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5723_ _5723_/A _7285_/B _5724_/B vssd1 vssd1 vccd1 vccd1 _5765_/A sky130_fd_sc_hd__and3_4
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5654_ _5654_/A _5654_/B vssd1 vssd1 vccd1 vccd1 _5697_/B sky130_fd_sc_hd__xnor2_4
XFILLER_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4605_ _7001_/A _4605_/B vssd1 vssd1 vccd1 vccd1 _4606_/C sky130_fd_sc_hd__xnor2_4
X_7324_ _7324_/A _7324_/B vssd1 vssd1 vccd1 vccd1 _7325_/B sky130_fd_sc_hd__nand2_1
X_5585_ _5585_/A _5585_/B vssd1 vssd1 vccd1 vccd1 _5588_/B sky130_fd_sc_hd__xnor2_4
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4536_ _4536_/A _4536_/B vssd1 vssd1 vccd1 vccd1 _4537_/B sky130_fd_sc_hd__xnor2_4
XFILLER_104_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7255_ _7256_/A _7256_/B vssd1 vssd1 vccd1 vccd1 _7255_/X sky130_fd_sc_hd__or2_1
X_4467_ _4467_/A _4516_/B _4467_/C vssd1 vssd1 vccd1 vccd1 _4467_/X sky130_fd_sc_hd__and3_2
XFILLER_89_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6206_ _6127_/A _6137_/X _6205_/X _6177_/A vssd1 vssd1 vccd1 vccd1 _6206_/X sky130_fd_sc_hd__a2bb2o_1
X_4398_ _4376_/A _4268_/X _4340_/A _4340_/B _4354_/A vssd1 vssd1 vccd1 vccd1 _4413_/B
+ sky130_fd_sc_hd__a221o_2
X_7186_ _7261_/A _7371_/B vssd1 vssd1 vccd1 vccd1 _7262_/A sky130_fd_sc_hd__nor2_4
XFILLER_98_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6137_ _6137_/A _6137_/B vssd1 vssd1 vccd1 vccd1 _6137_/X sky130_fd_sc_hd__xor2_4
XFILLER_100_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6068_ _6068_/A _6068_/B vssd1 vssd1 vccd1 vccd1 _6102_/A sky130_fd_sc_hd__nand2_4
XFILLER_93_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5019_ _5019_/A _5020_/B vssd1 vssd1 vccd1 vccd1 _5039_/A sky130_fd_sc_hd__and2_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5370_ _5445_/A _7210_/B vssd1 vssd1 vccd1 vccd1 _6970_/A sky130_fd_sc_hd__nor2_8
XFILLER_113_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4321_ _4312_/X _4314_/Y _4355_/B _4354_/A vssd1 vssd1 vccd1 vccd1 _6969_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4252_ _4192_/B _4260_/C _4251_/Y _4548_/B vssd1 vssd1 vccd1 vccd1 _4322_/B sky130_fd_sc_hd__a211o_2
Xfanout109 _5316_/Y vssd1 vssd1 vccd1 vccd1 _7344_/B sky130_fd_sc_hd__clkbuf_16
X_7040_ _7022_/A _7022_/B _7035_/A vssd1 vssd1 vccd1 vccd1 _7052_/A sky130_fd_sc_hd__a21bo_4
XFILLER_101_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4183_ _4183_/A _4183_/B vssd1 vssd1 vccd1 vccd1 _4210_/C sky130_fd_sc_hd__nor2_2
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7942_ _8041_/Q _7964_/C vssd1 vssd1 vccd1 vccd1 _7942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7873_ _7873_/A vssd1 vssd1 vccd1 vccd1 _7873_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6824_ _6824_/A _6824_/B vssd1 vssd1 vccd1 vccd1 _6828_/A sky130_fd_sc_hd__or2_1
XFILLER_63_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6755_ _6739_/S _6738_/Y _6739_/X _6751_/S _6584_/Y vssd1 vssd1 vccd1 vccd1 _6755_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5706_ _5706_/A _5706_/B vssd1 vssd1 vccd1 vccd1 _5748_/B sky130_fd_sc_hd__xor2_4
X_6686_ _6681_/B _6685_/Y _6739_/S vssd1 vssd1 vccd1 vccd1 _6686_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5637_ _5637_/A _5637_/B vssd1 vssd1 vccd1 vccd1 _5686_/A sky130_fd_sc_hd__xor2_4
X_5568_ _5569_/B _5568_/B vssd1 vssd1 vccd1 vccd1 _5570_/A sky130_fd_sc_hd__and2b_2
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7307_ _5977_/A _7284_/A _5271_/B _7210_/B _7311_/A vssd1 vssd1 vccd1 vccd1 _7307_/X
+ sky130_fd_sc_hd__o32a_2
XFILLER_2_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4519_ _4519_/A _4519_/B vssd1 vssd1 vccd1 vccd1 _4521_/B sky130_fd_sc_hd__xnor2_4
X_5499_ _5499_/A _5499_/B vssd1 vssd1 vccd1 vccd1 _6159_/A sky130_fd_sc_hd__xnor2_4
X_7238_ _7238_/A _7238_/B vssd1 vssd1 vccd1 vccd1 _7472_/A sky130_fd_sc_hd__xnor2_4
XFILLER_104_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7169_ _7169_/A _7169_/B vssd1 vssd1 vccd1 vccd1 _7176_/A sky130_fd_sc_hd__xnor2_4
XFILLER_100_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4870_ _4874_/B _4870_/B vssd1 vssd1 vccd1 vccd1 _4894_/B sky130_fd_sc_hd__and2b_2
X_6540_ _6562_/A _6540_/B vssd1 vssd1 vccd1 vccd1 _6588_/S sky130_fd_sc_hd__or2_4
X_6471_ _6355_/X _6469_/Y _7728_/A vssd1 vssd1 vccd1 vccd1 _6614_/A sky130_fd_sc_hd__a21oi_4
XFILLER_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5422_ _5422_/A _5422_/B vssd1 vssd1 vccd1 vccd1 _5423_/B sky130_fd_sc_hd__xor2_4
X_5353_ _5353_/A _5353_/B vssd1 vssd1 vccd1 vccd1 _5354_/B sky130_fd_sc_hd__xnor2_4
X_4304_ _4078_/A _4119_/Y _4084_/B _4111_/A vssd1 vssd1 vccd1 vccd1 _4304_/X sky130_fd_sc_hd__a211o_1
X_8072_ _8080_/CLK _8072_/D vssd1 vssd1 vccd1 vccd1 _8072_/Q sky130_fd_sc_hd__dfxtp_4
X_5284_ _5284_/A _5284_/B vssd1 vssd1 vccd1 vccd1 _5285_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4235_ _4241_/B _4227_/X _4231_/X _4187_/B vssd1 vssd1 vccd1 vccd1 _4235_/X sky130_fd_sc_hd__o211a_1
XFILLER_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7023_ _6873_/A _7306_/B _6970_/X vssd1 vssd1 vccd1 vccd1 _7024_/B sky130_fd_sc_hd__a21o_1
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4166_ _8077_/Q _4166_/B vssd1 vssd1 vccd1 vccd1 _4172_/B sky130_fd_sc_hd__xnor2_4
XFILLER_95_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4097_ _8055_/Q _4097_/B vssd1 vssd1 vccd1 vccd1 _4098_/B sky130_fd_sc_hd__xnor2_4
X_7925_ _6269_/X _7911_/Y _7918_/X _7924_/X vssd1 vssd1 vccd1 vccd1 _7925_/X sky130_fd_sc_hd__o211a_1
XFILLER_83_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7856_ _7856_/A _7856_/B vssd1 vssd1 vccd1 vccd1 _8038_/D sky130_fd_sc_hd__nor2_1
XFILLER_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6807_ _6807_/A _6819_/A vssd1 vssd1 vccd1 vccd1 _6809_/B sky130_fd_sc_hd__xnor2_1
X_7787_ _7787_/A _7787_/B vssd1 vssd1 vccd1 vccd1 _7787_/X sky130_fd_sc_hd__xor2_2
X_4999_ _4998_/A _5020_/B _4998_/C vssd1 vssd1 vccd1 vccd1 _5000_/B sky130_fd_sc_hd__a21oi_2
XFILLER_109_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6738_ _6570_/Y _6737_/B _6737_/Y vssd1 vssd1 vccd1 vccd1 _6738_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6669_ _6669_/A vssd1 vssd1 vccd1 vccd1 _6669_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout80 _7247_/C vssd1 vssd1 vccd1 vccd1 _5715_/A sky130_fd_sc_hd__buf_12
Xfanout91 _5088_/Y vssd1 vssd1 vccd1 vccd1 _7124_/A2 sky130_fd_sc_hd__buf_4
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4020_ _7974_/A _4020_/B vssd1 vssd1 vccd1 vccd1 _4020_/X sky130_fd_sc_hd__or2_2
XFILLER_96_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5971_ _6242_/S _6139_/B vssd1 vssd1 vccd1 vccd1 _6146_/A sky130_fd_sc_hd__nand2_2
X_7710_ _7462_/Y _7709_/Y _7847_/A vssd1 vssd1 vccd1 vccd1 _7748_/B sky130_fd_sc_hd__mux2_2
XFILLER_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4922_ _4921_/A _4931_/A _4921_/C vssd1 vssd1 vccd1 vccd1 _4925_/B sky130_fd_sc_hd__a21o_1
X_7641_ _7858_/B vssd1 vssd1 vccd1 vccd1 _7641_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4853_ _4866_/A _4866_/B vssd1 vssd1 vccd1 vccd1 _4867_/A sky130_fd_sc_hd__nand2_2
X_7572_ _7570_/B _6262_/X _7570_/Y _7639_/B vssd1 vssd1 vccd1 vccd1 _7572_/X sky130_fd_sc_hd__o211a_1
X_4784_ _4785_/B _4789_/A _4785_/A vssd1 vssd1 vccd1 vccd1 _4786_/A sky130_fd_sc_hd__o21ai_2
X_6523_ _6523_/A _6523_/B vssd1 vssd1 vccd1 vccd1 _6524_/B sky130_fd_sc_hd__xnor2_4
XFILLER_20_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6454_ _6492_/A _6452_/Y _6453_/Y _6364_/A vssd1 vssd1 vccd1 vccd1 _6454_/X sky130_fd_sc_hd__o211a_1
XFILLER_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5405_ _5294_/B _5399_/B _5343_/A _5343_/B vssd1 vssd1 vccd1 vccd1 _5410_/A sky130_fd_sc_hd__a2bb2o_4
X_6385_ _6878_/C _6878_/B _6456_/S vssd1 vssd1 vccd1 vccd1 _6387_/B sky130_fd_sc_hd__mux2_8
XFILLER_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5336_ _5336_/A _5336_/B vssd1 vssd1 vccd1 vccd1 _5503_/B sky130_fd_sc_hd__xnor2_4
XFILLER_114_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8055_ _8079_/CLK _8055_/D vssd1 vssd1 vccd1 vccd1 _8055_/Q sky130_fd_sc_hd__dfxtp_4
X_5267_ _5267_/A _5267_/B vssd1 vssd1 vccd1 vccd1 _5276_/A sky130_fd_sc_hd__xor2_4
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4218_ _4158_/X _4159_/Y _4210_/B vssd1 vssd1 vccd1 vccd1 _4218_/Y sky130_fd_sc_hd__a21oi_4
X_7006_ _7006_/A _7006_/B vssd1 vssd1 vccd1 vccd1 _7008_/B sky130_fd_sc_hd__xnor2_4
X_5198_ _5582_/A _5198_/B vssd1 vssd1 vccd1 vccd1 _5200_/B sky130_fd_sc_hd__or2_4
XFILLER_28_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4149_ _8081_/Q _4149_/B vssd1 vssd1 vccd1 vccd1 _4149_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7908_ _7908_/A _7930_/B _7907_/X vssd1 vssd1 vccd1 vccd1 _7929_/B sky130_fd_sc_hd__or3b_4
XFILLER_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7839_ _7887_/A _7839_/B _7839_/C vssd1 vssd1 vccd1 vccd1 _7839_/X sky130_fd_sc_hd__or3_1
XFILLER_51_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6170_ _6168_/X _6169_/X _6254_/S vssd1 vssd1 vccd1 vccd1 _6170_/X sky130_fd_sc_hd__mux2_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5121_ _5121_/A _5121_/B _5121_/C vssd1 vssd1 vccd1 vccd1 _5123_/A sky130_fd_sc_hd__and3_2
XFILLER_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5052_ _5703_/A _5703_/B _4978_/X _5378_/A vssd1 vssd1 vccd1 vccd1 _5054_/D sky130_fd_sc_hd__o211a_2
XFILLER_38_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5954_ _7949_/B _6805_/B vssd1 vssd1 vccd1 vccd1 _6354_/A sky130_fd_sc_hd__nor2_8
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4905_ _4905_/A _4939_/A vssd1 vssd1 vccd1 vccd1 _4909_/A sky130_fd_sc_hd__nand2_4
XFILLER_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5885_ _5885_/A _5885_/B vssd1 vssd1 vccd1 vccd1 _5886_/B sky130_fd_sc_hd__and2_1
X_7624_ _7766_/A _7411_/A _7624_/S vssd1 vssd1 vccd1 vccd1 _7624_/X sky130_fd_sc_hd__mux2_1
X_4836_ _4836_/A _4836_/B vssd1 vssd1 vccd1 vccd1 _4929_/A sky130_fd_sc_hd__xnor2_4
XFILLER_21_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7555_ _7553_/B _7554_/C _7554_/B vssd1 vssd1 vccd1 vccd1 _7556_/B sky130_fd_sc_hd__o21ai_1
XFILLER_119_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6506_ _6529_/A _6505_/X _6473_/Y vssd1 vssd1 vccd1 vccd1 _6506_/X sky130_fd_sc_hd__a21o_1
X_4767_ _5095_/B _4767_/B vssd1 vssd1 vccd1 vccd1 _4785_/A sky130_fd_sc_hd__and2_1
XFILLER_21_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7486_ _7484_/X _7485_/X _7535_/A vssd1 vssd1 vccd1 vccd1 _7544_/B sky130_fd_sc_hd__mux2_1
X_4698_ _4697_/B _4697_/C _4697_/A vssd1 vssd1 vccd1 vccd1 _4700_/B sky130_fd_sc_hd__o21ai_1
X_6437_ _6437_/A _6478_/B vssd1 vssd1 vccd1 vccd1 _6479_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6368_ _6368_/A _6368_/B _6359_/A vssd1 vssd1 vccd1 vccd1 _6368_/X sky130_fd_sc_hd__or3b_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5319_ _5582_/A _5797_/A vssd1 vssd1 vccd1 vccd1 _5325_/A sky130_fd_sc_hd__or2_4
X_6299_ _6299_/A _6299_/B vssd1 vssd1 vccd1 vccd1 _6308_/A sky130_fd_sc_hd__xnor2_4
X_8038_ _8082_/CLK _8038_/D vssd1 vssd1 vccd1 vccd1 _8038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_9 _7085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5670_ _5669_/B _5670_/B vssd1 vssd1 vccd1 vccd1 _5671_/B sky130_fd_sc_hd__and2b_1
XFILLER_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4621_ _7116_/A _5013_/B vssd1 vssd1 vccd1 vccd1 _4638_/B sky130_fd_sc_hd__nor2_4
XFILLER_116_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7340_ _7340_/A _7340_/B vssd1 vssd1 vccd1 vccd1 _7351_/B sky130_fd_sc_hd__xnor2_4
X_4552_ _4552_/A _4587_/A vssd1 vssd1 vccd1 vccd1 _4556_/A sky130_fd_sc_hd__nand2_4
X_4483_ _4483_/A _6999_/A _4662_/A vssd1 vssd1 vccd1 vccd1 _4483_/X sky130_fd_sc_hd__or3_1
XFILLER_7_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7271_ _7272_/B _7271_/B vssd1 vssd1 vccd1 vccd1 _7273_/A sky130_fd_sc_hd__nand2b_4
X_6222_ _6193_/A _6183_/X _6221_/X vssd1 vssd1 vccd1 vccd1 _6222_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6153_ _6199_/S _6151_/X _6152_/X vssd1 vssd1 vccd1 vccd1 _6153_/Y sky130_fd_sc_hd__o21ai_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6084_ _6084_/A _6088_/B vssd1 vssd1 vccd1 vccd1 _6086_/B sky130_fd_sc_hd__xor2_4
X_5104_ _6878_/B _5174_/B _5187_/B vssd1 vssd1 vccd1 vccd1 _5182_/B sky130_fd_sc_hd__and3_2
XFILLER_58_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _5034_/A _5034_/B _5034_/C vssd1 vssd1 vccd1 vccd1 _5035_/X sky130_fd_sc_hd__a21o_1
XFILLER_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6986_ _6991_/B _6991_/C _6991_/A vssd1 vssd1 vccd1 vccd1 _6992_/A sky130_fd_sc_hd__o21ai_4
XFILLER_41_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5937_ _5847_/A _5847_/B _6227_/A _6227_/B _5846_/Y vssd1 vssd1 vccd1 vccd1 _6205_/B
+ sky130_fd_sc_hd__a41o_4
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7607_ _7607_/A _7607_/B vssd1 vssd1 vccd1 vccd1 _7607_/X sky130_fd_sc_hd__and2_1
X_5868_ _5868_/A _5869_/A _5868_/C vssd1 vssd1 vccd1 vccd1 _5893_/A sky130_fd_sc_hd__nand3_2
X_4819_ _5014_/A _4923_/B vssd1 vssd1 vccd1 vccd1 _4926_/A sky130_fd_sc_hd__nor2_8
X_5799_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5799_/Y sky130_fd_sc_hd__inv_2
X_7538_ _7484_/X _7531_/C _7538_/S vssd1 vssd1 vccd1 vccd1 _7542_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7469_ _7465_/X _7468_/X _7535_/A vssd1 vssd1 vccd1 vccd1 _7537_/C sky130_fd_sc_hd__mux2_1
XFILLER_115_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _8079_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6840_ _7025_/A _6839_/B _6871_/B vssd1 vssd1 vccd1 vccd1 _6841_/B sky130_fd_sc_hd__o21ai_1
XFILLER_35_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6771_ _4005_/Y _5107_/X _6770_/Y vssd1 vssd1 vccd1 vccd1 _6771_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5722_ _5722_/A _5722_/B _7085_/B vssd1 vssd1 vccd1 vccd1 _5724_/B sky130_fd_sc_hd__and3_2
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5653_ _5654_/A _5654_/B vssd1 vssd1 vccd1 vccd1 _5653_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_30_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5584_ _5185_/Y _5919_/A _5576_/B _5574_/Y vssd1 vssd1 vccd1 vccd1 _5588_/A sky130_fd_sc_hd__a31o_4
X_4604_ _4604_/A _4604_/B vssd1 vssd1 vccd1 vccd1 _4605_/B sky130_fd_sc_hd__xnor2_4
XFILLER_116_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7323_ _7324_/A _7324_/B vssd1 vssd1 vccd1 vccd1 _7323_/Y sky130_fd_sc_hd__nor2_1
X_4535_ _4508_/A _4508_/B _4509_/B _4509_/A vssd1 vssd1 vccd1 vccd1 _4536_/B sky130_fd_sc_hd__o2bb2ai_4
XFILLER_116_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7254_ _7311_/A _7294_/B _7311_/C vssd1 vssd1 vccd1 vccd1 _7256_/B sky130_fd_sc_hd__or3_4
X_4466_ _4516_/A _4465_/C _4465_/A vssd1 vssd1 vccd1 vccd1 _4467_/C sky130_fd_sc_hd__a21o_1
X_4397_ _4430_/C _4396_/B _4436_/A vssd1 vssd1 vccd1 vccd1 _4397_/Y sky130_fd_sc_hd__a21oi_2
X_7185_ _7185_/A _7185_/B vssd1 vssd1 vccd1 vccd1 _7188_/A sky130_fd_sc_hd__or2_4
X_6205_ _6205_/A _6205_/B vssd1 vssd1 vccd1 vccd1 _6205_/X sky130_fd_sc_hd__xor2_4
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _6205_/A _6205_/B _5787_/A vssd1 vssd1 vccd1 vccd1 _6137_/B sky130_fd_sc_hd__a21oi_4
XFILLER_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _6067_/A _7426_/A vssd1 vssd1 vccd1 vccd1 _6068_/B sky130_fd_sc_hd__nand2_2
XFILLER_54_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5018_ _5018_/A _5018_/B _5018_/C vssd1 vssd1 vccd1 vccd1 _5018_/X sky130_fd_sc_hd__and3_2
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6969_ _6969_/A _7210_/B vssd1 vssd1 vccd1 vccd1 _7086_/A sky130_fd_sc_hd__or2_4
XFILLER_41_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4320_ _4312_/X _4314_/Y _4356_/B _4356_/A vssd1 vssd1 vccd1 vccd1 _4320_/X sky130_fd_sc_hd__o22a_4
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4251_ _4209_/X _4226_/X _4232_/Y _4200_/B vssd1 vssd1 vccd1 vccd1 _4251_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_113_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4182_ _4228_/A _4228_/B _4178_/X vssd1 vssd1 vccd1 vccd1 _4183_/B sky130_fd_sc_hd__o21a_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7941_ _7918_/B _7940_/Y _7903_/B1 vssd1 vssd1 vccd1 vccd1 _7941_/X sky130_fd_sc_hd__o21ba_1
XFILLER_82_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7872_ _7872_/A _7872_/B vssd1 vssd1 vccd1 vccd1 _7873_/A sky130_fd_sc_hd__xnor2_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6823_ _6833_/A _6823_/B vssd1 vssd1 vccd1 vccd1 _6831_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6754_ _6745_/X _6753_/X _7616_/S vssd1 vssd1 vccd1 vccd1 _6757_/D sky130_fd_sc_hd__mux2_1
X_6685_ _6695_/S _6659_/B _6684_/X vssd1 vssd1 vccd1 vccd1 _6685_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5705_ _5908_/A _6951_/D _5908_/C vssd1 vssd1 vccd1 vccd1 _5748_/A sky130_fd_sc_hd__and3_2
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5636_ _5637_/A _5637_/B vssd1 vssd1 vccd1 vccd1 _5636_/Y sky130_fd_sc_hd__nand2_1
X_5567_ _5566_/A _5566_/B _5619_/A _5619_/B vssd1 vssd1 vccd1 vccd1 _5568_/B sky130_fd_sc_hd__a22o_1
XFILLER_117_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5498_ _5498_/A _5498_/B vssd1 vssd1 vccd1 vccd1 _5499_/B sky130_fd_sc_hd__xnor2_4
XFILLER_2_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4518_ _7214_/A _4518_/B vssd1 vssd1 vccd1 vccd1 _4519_/B sky130_fd_sc_hd__xnor2_4
X_7306_ _7306_/A _7306_/B _7306_/C vssd1 vssd1 vccd1 vccd1 _7332_/A sky130_fd_sc_hd__and3_4
X_4449_ _4642_/A _4630_/B _4448_/Y vssd1 vssd1 vccd1 vccd1 _4451_/B sky130_fd_sc_hd__or3b_2
X_7237_ _7238_/B _7238_/A vssd1 vssd1 vccd1 vccd1 _7237_/X sky130_fd_sc_hd__and2b_1
XFILLER_104_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7168_ _7169_/A _7169_/B vssd1 vssd1 vccd1 vccd1 _7184_/A sky130_fd_sc_hd__nand2_1
XFILLER_100_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ _7099_/A _7099_/B vssd1 vssd1 vccd1 vccd1 _7102_/B sky130_fd_sc_hd__and2_2
X_6119_ _6117_/X _6118_/Y _6174_/A vssd1 vssd1 vccd1 vccd1 _6120_/B sky130_fd_sc_hd__a21oi_2
XFILLER_100_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6470_ _7949_/B _6805_/B _6355_/X vssd1 vssd1 vccd1 vccd1 _6514_/A sky130_fd_sc_hd__a21bo_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5421_ _5421_/A _5421_/B vssd1 vssd1 vccd1 vccd1 _5422_/B sky130_fd_sc_hd__xor2_4
XFILLER_114_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5352_ _5352_/A _5352_/B _7269_/B vssd1 vssd1 vccd1 vccd1 _5353_/B sky130_fd_sc_hd__and3_2
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8071_ _8079_/CLK _8071_/D vssd1 vssd1 vccd1 vccd1 _8071_/Q sky130_fd_sc_hd__dfxtp_4
X_4303_ _8051_/Q _4303_/B _4303_/C vssd1 vssd1 vccd1 vccd1 _5145_/B sky130_fd_sc_hd__nand3_1
XFILLER_99_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5283_ _5498_/A _5498_/B vssd1 vssd1 vccd1 vccd1 _5287_/A sky130_fd_sc_hd__nor2_1
X_7022_ _7022_/A _7022_/B vssd1 vssd1 vccd1 vccd1 _7034_/A sky130_fd_sc_hd__xnor2_1
X_4234_ _4209_/X _4226_/X _4232_/Y vssd1 vssd1 vccd1 vccd1 _4234_/X sky130_fd_sc_hd__a21o_1
X_4165_ _8076_/Q _8075_/Q _4175_/B _4147_/B _4211_/B vssd1 vssd1 vccd1 vccd1 _4166_/B
+ sky130_fd_sc_hd__o41a_4
XFILLER_68_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4096_ _4096_/A _4096_/B vssd1 vssd1 vccd1 vccd1 _4097_/B sky130_fd_sc_hd__nand2_2
XFILLER_83_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7924_ _7935_/A _7900_/X _7921_/Y _7923_/Y vssd1 vssd1 vccd1 vccd1 _7924_/X sky130_fd_sc_hd__a31o_1
XFILLER_82_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7855_ _8038_/Q _7944_/B _7853_/X _7854_/X vssd1 vssd1 vccd1 vccd1 _7856_/B sky130_fd_sc_hd__a22oi_1
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6806_ _6806_/A _7025_/A vssd1 vssd1 vccd1 vccd1 _6819_/A sky130_fd_sc_hd__nor2_1
X_7786_ _7833_/A _7833_/B _7785_/Y vssd1 vssd1 vccd1 vccd1 _7787_/B sky130_fd_sc_hd__a21oi_4
XFILLER_51_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4998_ _4998_/A _5020_/B _4998_/C vssd1 vssd1 vccd1 vccd1 _5009_/A sky130_fd_sc_hd__and3_4
XFILLER_23_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6737_ _6572_/Y _6737_/B vssd1 vssd1 vccd1 vccd1 _6737_/Y sky130_fd_sc_hd__nand2b_1
X_6668_ _6667_/X _6664_/Y _6691_/A vssd1 vssd1 vccd1 vccd1 _6669_/A sky130_fd_sc_hd__mux2_1
X_6599_ _6626_/B _6626_/C _6626_/A vssd1 vssd1 vccd1 vccd1 _6627_/A sky130_fd_sc_hd__o21ai_4
X_5619_ _5619_/A _5619_/B vssd1 vssd1 vccd1 vccd1 _5627_/A sky130_fd_sc_hd__xnor2_4
XFILLER_3_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout81 _7247_/C vssd1 vssd1 vccd1 vccd1 _6839_/B sky130_fd_sc_hd__buf_2
Xfanout70 _4308_/X vssd1 vssd1 vccd1 vccd1 _7101_/A sky130_fd_sc_hd__buf_6
Xfanout92 _4447_/Y vssd1 vssd1 vccd1 vccd1 _5040_/A sky130_fd_sc_hd__buf_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5970_ _5970_/A _5970_/B _6139_/B vssd1 vssd1 vccd1 vccd1 _6177_/A sky130_fd_sc_hd__and3_4
XFILLER_18_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4921_ _4921_/A _4931_/A _4921_/C vssd1 vssd1 vccd1 vccd1 _4931_/B sky130_fd_sc_hd__nand3_4
X_7640_ _7639_/B _6263_/X _7639_/Y vssd1 vssd1 vccd1 vccd1 _7858_/B sky130_fd_sc_hd__o21a_2
X_4852_ _4857_/A _4852_/B vssd1 vssd1 vccd1 vccd1 _4866_/B sky130_fd_sc_hd__and2_1
XFILLER_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7571_ _7570_/B _6262_/X _7570_/Y vssd1 vssd1 vccd1 vccd1 _7571_/X sky130_fd_sc_hd__o21a_2
X_4783_ _4832_/A _4783_/B vssd1 vssd1 vccd1 vccd1 _4789_/A sky130_fd_sc_hd__and2b_1
XFILLER_118_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6522_ _6466_/Y _6509_/X _6522_/S vssd1 vssd1 vccd1 vccd1 _6523_/B sky130_fd_sc_hd__mux2_4
XFILLER_119_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6453_ _6492_/A _6453_/B vssd1 vssd1 vccd1 vccd1 _6453_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5404_ _5330_/B _5407_/B _5354_/B _5354_/A vssd1 vssd1 vccd1 vccd1 _5411_/A sky130_fd_sc_hd__a22oi_4
X_6384_ _6386_/A _6386_/B vssd1 vssd1 vccd1 vccd1 _6387_/A sky130_fd_sc_hd__nand2_4
X_5335_ _5335_/A _5335_/B vssd1 vssd1 vccd1 vccd1 _5336_/B sky130_fd_sc_hd__xor2_4
X_8054_ _8063_/CLK _8054_/D vssd1 vssd1 vccd1 vccd1 _8054_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5266_ _5264_/A _5275_/A _5265_/Y vssd1 vssd1 vccd1 vccd1 _5267_/B sky130_fd_sc_hd__a21o_2
XFILLER_102_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4217_ _4227_/S _4215_/Y _4216_/X _4193_/Y vssd1 vssd1 vccd1 vccd1 _4217_/Y sky130_fd_sc_hd__o31ai_4
X_7005_ _7016_/A _7016_/B vssd1 vssd1 vccd1 vccd1 _7036_/B sky130_fd_sc_hd__nand2_2
X_5197_ _5352_/A _5352_/B _6878_/B vssd1 vssd1 vccd1 vccd1 _5245_/A sky130_fd_sc_hd__and3_4
XFILLER_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4148_ _4147_/A _4147_/B _4147_/C _4147_/D _4168_/B1 vssd1 vssd1 vccd1 vccd1 _4149_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4079_ _4111_/A _4079_/B vssd1 vssd1 vccd1 vccd1 _4081_/B sky130_fd_sc_hd__or2_4
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7907_ _7858_/B _7883_/A _7883_/C _7698_/X _7930_/A vssd1 vssd1 vccd1 vccd1 _7907_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_70_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7838_ _7887_/A _7839_/C _7839_/B vssd1 vssd1 vccd1 vccd1 _7838_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7769_ _7769_/A _7769_/B vssd1 vssd1 vccd1 vccd1 _7770_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5120_ _4998_/A _4752_/Y _5119_/X vssd1 vssd1 vccd1 vccd1 _5121_/C sky130_fd_sc_hd__a21o_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5051_ _5378_/A _5908_/A _5378_/C vssd1 vssd1 vccd1 vccd1 _5379_/A sky130_fd_sc_hd__a21oi_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5953_ _5285_/A _5288_/A _5238_/B vssd1 vssd1 vccd1 vccd1 _6180_/B sky130_fd_sc_hd__a21bo_1
XFILLER_53_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4904_ _4938_/A _4938_/B vssd1 vssd1 vccd1 vccd1 _4939_/A sky130_fd_sc_hd__nand2_2
X_5884_ _5927_/C _5884_/B _5884_/C vssd1 vssd1 vccd1 vccd1 _5904_/A sky130_fd_sc_hd__or3_4
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7623_ _7623_/A _7623_/B vssd1 vssd1 vccd1 vccd1 _7656_/A sky130_fd_sc_hd__nor2_1
X_4835_ _4851_/A _4926_/A vssd1 vssd1 vccd1 vccd1 _4857_/A sky130_fd_sc_hd__nand2_2
X_7554_ _7554_/A _7554_/B _7554_/C vssd1 vssd1 vccd1 vccd1 _7597_/A sky130_fd_sc_hd__or3_4
X_4766_ _4832_/A _4766_/B vssd1 vssd1 vccd1 vccd1 _4767_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6505_ _6419_/A _6504_/Y _6417_/X vssd1 vssd1 vccd1 vccd1 _6505_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7485_ _7466_/X _7464_/X _7515_/S vssd1 vssd1 vccd1 vccd1 _7485_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4697_ _4697_/A _4697_/B _4697_/C vssd1 vssd1 vccd1 vccd1 _4700_/A sky130_fd_sc_hd__or3_4
X_6436_ _6437_/A _6478_/B vssd1 vssd1 vccd1 vccd1 _6479_/A sky130_fd_sc_hd__and2_2
XFILLER_20_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6367_ _7114_/B _7085_/A _6445_/S vssd1 vssd1 vccd1 vccd1 _6368_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5318_ _5582_/A _6971_/B vssd1 vssd1 vccd1 vccd1 _5330_/A sky130_fd_sc_hd__or2_4
XFILLER_114_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6298_ _6564_/A _6305_/A _6304_/A vssd1 vssd1 vccd1 vccd1 _6299_/B sky130_fd_sc_hd__a21o_2
XFILLER_102_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8037_ _8082_/CLK _8037_/D vssd1 vssd1 vccd1 vccd1 _8037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5249_ _5745_/A _5338_/B vssd1 vssd1 vccd1 vccd1 _5399_/A sky130_fd_sc_hd__nand2_4
XFILLER_56_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _4620_/A _4625_/A vssd1 vssd1 vccd1 vccd1 _4638_/A sky130_fd_sc_hd__nand2_4
XFILLER_30_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4551_ _4551_/A _4551_/B _4552_/A _4551_/D vssd1 vssd1 vccd1 vccd1 _4587_/A sky130_fd_sc_hd__nand4_4
XFILLER_116_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7270_ _7371_/A _7247_/C _7274_/A _7268_/B _7268_/A vssd1 vssd1 vccd1 vccd1 _7272_/B
+ sky130_fd_sc_hd__o32a_1
X_4482_ _4412_/A _4413_/B _4436_/A vssd1 vssd1 vccd1 vccd1 _4482_/Y sky130_fd_sc_hd__a21oi_1
X_6221_ _6012_/B _6262_/S _6167_/X _6254_/S vssd1 vssd1 vccd1 vccd1 _6221_/X sky130_fd_sc_hd__o211a_1
XFILLER_112_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6152_ _6081_/Y _6111_/B _6111_/C _6149_/X vssd1 vssd1 vccd1 vccd1 _6152_/X sky130_fd_sc_hd__a31o_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5103_ _5110_/A _5103_/B vssd1 vssd1 vccd1 vccd1 _5187_/B sky130_fd_sc_hd__xnor2_4
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6083_ _6077_/A _6077_/B _6088_/A vssd1 vssd1 vccd1 vccd1 _6086_/A sky130_fd_sc_hd__a21oi_4
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5034_/A _5034_/B _5034_/C vssd1 vssd1 vccd1 vccd1 _5034_/X sky130_fd_sc_hd__and3_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6985_ _6993_/B _6993_/A vssd1 vssd1 vccd1 vccd1 _6991_/C sky130_fd_sc_hd__and2b_1
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5936_ _6227_/A _6227_/B vssd1 vssd1 vccd1 vccd1 _6228_/B sky130_fd_sc_hd__nand2_1
X_7606_ _7576_/A _7569_/C _7576_/Y vssd1 vssd1 vccd1 vccd1 _7607_/B sky130_fd_sc_hd__a21o_1
X_5867_ _5866_/A _5866_/B _5866_/C vssd1 vssd1 vccd1 vccd1 _5868_/C sky130_fd_sc_hd__o21ai_2
X_4818_ _4851_/A _4818_/B vssd1 vssd1 vccd1 vccd1 _4818_/Y sky130_fd_sc_hd__nor2_1
X_5798_ _5855_/C _5798_/B _5798_/C vssd1 vssd1 vccd1 vccd1 _5840_/A sky130_fd_sc_hd__and3b_4
X_7537_ _7766_/B _7537_/B _7537_/C _7537_/D vssd1 vssd1 vccd1 vccd1 _7537_/X sky130_fd_sc_hd__or4_1
X_4749_ _5445_/A _4751_/C _4850_/A vssd1 vssd1 vccd1 vccd1 _4854_/A sky130_fd_sc_hd__or3_4
XFILLER_107_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7468_ _7467_/X _7466_/X _7624_/S vssd1 vssd1 vccd1 vccd1 _7468_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6419_ _6419_/A _6419_/B vssd1 vssd1 vccd1 vccd1 _6533_/A sky130_fd_sc_hd__nand2_4
X_7399_ _7403_/A vssd1 vssd1 vccd1 vccd1 _7411_/A sky130_fd_sc_hd__clkinv_2
XFILLER_103_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6770_ _6770_/A _7949_/B vssd1 vssd1 vccd1 vccd1 _6770_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5721_ _5723_/A _7085_/B vssd1 vssd1 vccd1 vccd1 _5761_/A sky130_fd_sc_hd__and2_2
X_5652_ _5652_/A _5652_/B vssd1 vssd1 vccd1 vccd1 _5654_/B sky130_fd_sc_hd__xnor2_4
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5583_ _5639_/A _5639_/B vssd1 vssd1 vccd1 vccd1 _5589_/A sky130_fd_sc_hd__or2_4
X_4603_ _4604_/A _4604_/B vssd1 vssd1 vccd1 vccd1 _4603_/Y sky130_fd_sc_hd__nand2_1
X_7322_ _7320_/A _7327_/A _7327_/B _7321_/Y vssd1 vssd1 vccd1 vccd1 _7324_/B sky130_fd_sc_hd__o31a_1
X_4534_ _4795_/B _4534_/B vssd1 vssd1 vccd1 vccd1 _4536_/A sky130_fd_sc_hd__xnor2_4
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7253_ _7285_/A _7281_/D vssd1 vssd1 vccd1 vccd1 _7311_/C sky130_fd_sc_hd__nand2_2
X_4465_ _4465_/A _4516_/A _4465_/C vssd1 vssd1 vccd1 vccd1 _4516_/B sky130_fd_sc_hd__nand3_4
X_6204_ _6250_/A _6203_/Y _6226_/S vssd1 vssd1 vccd1 vccd1 _6255_/B sky130_fd_sc_hd__mux2_2
X_7184_ _7184_/A _7184_/B _7184_/C vssd1 vssd1 vccd1 vccd1 _7185_/B sky130_fd_sc_hd__and3_1
X_4396_ _4436_/A _4396_/B vssd1 vssd1 vccd1 vccd1 _4396_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6135_ _6135_/A _6135_/B vssd1 vssd1 vccd1 vccd1 _6135_/Y sky130_fd_sc_hd__xnor2_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6066_ _6067_/A _7426_/A vssd1 vssd1 vccd1 vccd1 _6068_/A sky130_fd_sc_hd__or2_2
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _5016_/B _5016_/C _5016_/A vssd1 vssd1 vccd1 vccd1 _5018_/C sky130_fd_sc_hd__a21bo_1
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6968_ _6968_/A _6968_/B vssd1 vssd1 vccd1 vccd1 _6975_/A sky130_fd_sc_hd__xnor2_4
X_6899_ _7306_/A _6951_/D vssd1 vssd1 vccd1 vccd1 _6943_/B sky130_fd_sc_hd__nand2_1
XFILLER_42_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5919_ _5919_/A _5927_/B _5919_/C vssd1 vssd1 vccd1 vccd1 _5919_/X sky130_fd_sc_hd__and3_1
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4250_ _4209_/X _4226_/X _4232_/Y _4204_/Y vssd1 vssd1 vccd1 vccd1 _4250_/X sky130_fd_sc_hd__a211o_1
X_4181_ _4216_/B _4228_/B _4178_/X vssd1 vssd1 vccd1 vccd1 _4183_/A sky130_fd_sc_hd__a21oi_1
X_7940_ _7940_/A _7940_/B vssd1 vssd1 vccd1 vccd1 _7940_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7871_ _7872_/A _7872_/B vssd1 vssd1 vccd1 vccd1 _7913_/A sky130_fd_sc_hd__or2_4
X_6822_ _6824_/B _6822_/B vssd1 vssd1 vccd1 vccd1 _6823_/B sky130_fd_sc_hd__xor2_4
XFILLER_63_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6753_ _6751_/X _6703_/X _6753_/S vssd1 vssd1 vccd1 vccd1 _6753_/X sky130_fd_sc_hd__mux2_1
X_6684_ _6695_/S _6683_/X _6645_/B _6641_/B vssd1 vssd1 vccd1 vccd1 _6684_/X sky130_fd_sc_hd__a2bb2o_1
X_5704_ _5908_/A _5908_/C vssd1 vssd1 vccd1 vccd1 _5927_/B sky130_fd_sc_hd__and2_4
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5635_ _5635_/A _5635_/B vssd1 vssd1 vccd1 vccd1 _5637_/B sky130_fd_sc_hd__xor2_4
X_5566_ _5566_/A _5566_/B vssd1 vssd1 vccd1 vccd1 _5619_/B sky130_fd_sc_hd__xor2_4
X_5497_ _5497_/A _5497_/B vssd1 vssd1 vccd1 vccd1 _6155_/A sky130_fd_sc_hd__xnor2_2
X_4517_ _4517_/A _4517_/B vssd1 vssd1 vccd1 vccd1 _4518_/B sky130_fd_sc_hd__nand2_4
X_7305_ _7366_/A _7358_/B vssd1 vssd1 vccd1 vccd1 _7306_/C sky130_fd_sc_hd__nor2_1
X_4448_ _4662_/A _4988_/A vssd1 vssd1 vccd1 vccd1 _4448_/Y sky130_fd_sc_hd__nor2_1
X_7236_ _7239_/A _7239_/B _7234_/A _7234_/B vssd1 vssd1 vccd1 vccd1 _7238_/B sky130_fd_sc_hd__o2bb2a_2
XFILLER_58_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7167_ _7167_/A _7167_/B vssd1 vssd1 vccd1 vccd1 _7169_/B sky130_fd_sc_hd__xnor2_4
X_4379_ _4412_/A _4407_/B _4396_/B _4455_/A _4377_/A vssd1 vssd1 vccd1 vccd1 _4379_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_85_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6118_ _6118_/A _6118_/B vssd1 vssd1 vccd1 vccd1 _6118_/Y sky130_fd_sc_hd__nand2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ _7108_/A _7108_/B vssd1 vssd1 vccd1 vccd1 _7099_/B sky130_fd_sc_hd__nand2b_1
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6049_ _6031_/A _6031_/B _6060_/A vssd1 vssd1 vccd1 vccd1 _6051_/S sky130_fd_sc_hd__a21o_1
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5420_ _5421_/B _5421_/A vssd1 vssd1 vccd1 vccd1 _5420_/Y sky130_fd_sc_hd__nand2b_1
X_5351_ _5582_/A _5715_/A vssd1 vssd1 vccd1 vccd1 _5407_/B sky130_fd_sc_hd__nor2_8
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8070_ _8075_/CLK _8070_/D vssd1 vssd1 vccd1 vccd1 _8070_/Q sky130_fd_sc_hd__dfxtp_4
X_4302_ _4296_/Y _4301_/Y _5087_/B vssd1 vssd1 vccd1 vccd1 _4302_/X sky130_fd_sc_hd__mux2_1
X_5282_ _5492_/A _5281_/B _5278_/Y vssd1 vssd1 vccd1 vccd1 _5498_/B sky130_fd_sc_hd__a21oi_4
XFILLER_99_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4233_ _4209_/X _4226_/X _4232_/Y vssd1 vssd1 vccd1 vccd1 _5990_/B sky130_fd_sc_hd__a21oi_4
X_7021_ _7021_/A _7021_/B vssd1 vssd1 vccd1 vccd1 _7022_/B sky130_fd_sc_hd__xnor2_2
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4164_ _4158_/X _4159_/Y _4230_/C vssd1 vssd1 vccd1 vccd1 _4164_/X sky130_fd_sc_hd__a21o_1
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4095_ _4095_/A _4095_/B vssd1 vssd1 vccd1 vccd1 _4103_/A sky130_fd_sc_hd__nand2_1
X_7923_ _7923_/A _7935_/B vssd1 vssd1 vccd1 vccd1 _7923_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7854_ _8037_/Q _7964_/C _7991_/D vssd1 vssd1 vccd1 vccd1 _7854_/X sky130_fd_sc_hd__a21bo_1
XFILLER_51_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7785_ _7833_/A _7833_/B _7908_/A vssd1 vssd1 vccd1 vccd1 _7785_/Y sky130_fd_sc_hd__o21bai_2
X_6805_ _7027_/A _6805_/B vssd1 vssd1 vccd1 vccd1 _6809_/A sky130_fd_sc_hd__nor2_1
X_6736_ _6701_/B _6735_/X _7583_/S vssd1 vssd1 vccd1 vccd1 _6757_/A sky130_fd_sc_hd__mux2_1
X_4997_ _4957_/B _5022_/A _4992_/A _4992_/B vssd1 vssd1 vccd1 vccd1 _4998_/C sky130_fd_sc_hd__o22ai_4
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6667_ _6666_/Y _6647_/A _6689_/S vssd1 vssd1 vccd1 vccd1 _6667_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6598_ _6617_/B _6617_/C _6617_/A vssd1 vssd1 vccd1 vccd1 _6626_/C sky130_fd_sc_hd__o21a_2
X_5618_ _5618_/A _5618_/B vssd1 vssd1 vccd1 vccd1 _5657_/A sky130_fd_sc_hd__xnor2_4
XFILLER_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5549_ _5549_/A _5549_/B vssd1 vssd1 vccd1 vccd1 _5560_/B sky130_fd_sc_hd__xor2_2
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7219_ _7219_/A _7219_/B vssd1 vssd1 vccd1 vccd1 _7242_/A sky130_fd_sc_hd__xor2_1
XFILLER_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout71 _7622_/A vssd1 vssd1 vccd1 vccd1 _7649_/A sky130_fd_sc_hd__buf_4
Xfanout60 _6364_/A vssd1 vssd1 vccd1 vccd1 _6443_/A sky130_fd_sc_hd__buf_6
Xfanout82 _5147_/X vssd1 vssd1 vccd1 vccd1 _7247_/C sky130_fd_sc_hd__buf_8
Xfanout93 _4446_/X vssd1 vssd1 vccd1 vccd1 _5014_/A sky130_fd_sc_hd__buf_8
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4920_ _4920_/A _5040_/B vssd1 vssd1 vccd1 vccd1 _4921_/C sky130_fd_sc_hd__and2_2
X_4851_ _4851_/A _4926_/A _4927_/A vssd1 vssd1 vccd1 vccd1 _4852_/B sky130_fd_sc_hd__or3_1
XFILLER_33_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7570_ _7639_/A _7570_/B vssd1 vssd1 vccd1 vccd1 _7570_/Y sky130_fd_sc_hd__nand2_1
X_4782_ _4782_/A _4782_/B vssd1 vssd1 vccd1 vccd1 _4783_/B sky130_fd_sc_hd__xnor2_1
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6521_ _6521_/A vssd1 vssd1 vccd1 vccd1 _6524_/A sky130_fd_sc_hd__inv_2
XFILLER_20_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6452_ _6451_/A _6450_/Y _6451_/Y vssd1 vssd1 vccd1 vccd1 _6452_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5403_ _5403_/A _5403_/B vssd1 vssd1 vccd1 vccd1 _5412_/A sky130_fd_sc_hd__xnor2_4
X_6383_ _6492_/A _6383_/B vssd1 vssd1 vccd1 vccd1 _6386_/B sky130_fd_sc_hd__nor2_2
XFILLER_88_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5334_ _5335_/A _5335_/B vssd1 vssd1 vccd1 vccd1 _5334_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8053_ _8077_/CLK _8053_/D vssd1 vssd1 vccd1 vccd1 _8053_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5265_ _5265_/A _5265_/B vssd1 vssd1 vccd1 vccd1 _5265_/Y sky130_fd_sc_hd__nand2_1
X_4216_ _8067_/Q _4216_/B _4216_/C _4221_/B vssd1 vssd1 vccd1 vccd1 _4216_/X sky130_fd_sc_hd__and4_1
XFILLER_68_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5196_ _5196_/A _5196_/B vssd1 vssd1 vccd1 vccd1 _5202_/A sky130_fd_sc_hd__xnor2_4
X_7004_ _7056_/A _7056_/B vssd1 vssd1 vccd1 vccd1 _7016_/B sky130_fd_sc_hd__nor2_1
X_4147_ _4147_/A _4147_/B _4147_/C _4147_/D vssd1 vssd1 vccd1 vccd1 _4352_/B sky130_fd_sc_hd__or4_4
XFILLER_95_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4078_ _4078_/A _4078_/B vssd1 vssd1 vccd1 vccd1 _4079_/B sky130_fd_sc_hd__nand2_2
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7906_ _7930_/A _7698_/X _7883_/A _7883_/B _7883_/C vssd1 vssd1 vccd1 vccd1 _7930_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_71_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7837_ _7837_/A _7837_/B vssd1 vssd1 vccd1 vccd1 _7839_/C sky130_fd_sc_hd__and2_1
XFILLER_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7768_ _7769_/A _7769_/B vssd1 vssd1 vccd1 vccd1 _7798_/A sky130_fd_sc_hd__or2_1
X_6719_ _6719_/A vssd1 vssd1 vccd1 vccd1 _6719_/Y sky130_fd_sc_hd__inv_2
X_7699_ _7639_/B _7571_/X _7639_/Y _7784_/A vssd1 vssd1 vccd1 vccd1 _7699_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5050_ _5050_/A _5054_/C vssd1 vssd1 vccd1 vccd1 _5378_/C sky130_fd_sc_hd__or2_1
XFILLER_85_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5952_ _5951_/A _5951_/B _5951_/C _6173_/A _6172_/A vssd1 vssd1 vccd1 vccd1 _6180_/A
+ sky130_fd_sc_hd__a311o_2
XFILLER_65_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4903_ _4903_/A _4903_/B vssd1 vssd1 vccd1 vccd1 _4938_/B sky130_fd_sc_hd__xnor2_1
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5883_ _7306_/B _5925_/B _5885_/B vssd1 vssd1 vccd1 vccd1 _5884_/C sky130_fd_sc_hd__a21oi_1
X_7622_ _7622_/A _7622_/B _7648_/C vssd1 vssd1 vccd1 vccd1 _7622_/X sky130_fd_sc_hd__or3_1
X_4834_ _4851_/A _4927_/A vssd1 vssd1 vccd1 vccd1 _4879_/A sky130_fd_sc_hd__xnor2_1
X_7553_ _7554_/C _7553_/B vssd1 vssd1 vccd1 vccd1 _7590_/A sky130_fd_sc_hd__and2b_1
X_4765_ _4832_/A _4766_/B vssd1 vssd1 vccd1 vccd1 _5095_/B sky130_fd_sc_hd__or2_1
XFILLER_119_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6504_ _6477_/Y _6503_/Y _6475_/X vssd1 vssd1 vccd1 vccd1 _6504_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_119_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7484_ _7463_/X _7483_/X _7624_/S vssd1 vssd1 vccd1 vccd1 _7484_/X sky130_fd_sc_hd__mux2_1
X_4696_ _4606_/Y _4693_/X _4650_/B _4648_/B vssd1 vssd1 vccd1 vccd1 _4697_/C sky130_fd_sc_hd__o211a_1
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6435_ _7306_/A _7281_/D _6456_/S vssd1 vssd1 vccd1 vccd1 _6478_/B sky130_fd_sc_hd__mux2_2
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6366_ _6468_/A _6468_/B vssd1 vssd1 vccd1 vccd1 _6366_/Y sky130_fd_sc_hd__nor2_2
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5317_ _5352_/A _5352_/B _5919_/A vssd1 vssd1 vccd1 vccd1 _5531_/A sky130_fd_sc_hd__and3_2
X_8036_ _8082_/CLK _8036_/D vssd1 vssd1 vccd1 vccd1 _8036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6297_ _6296_/X _6020_/A _6767_/S vssd1 vssd1 vccd1 vccd1 _6305_/A sky130_fd_sc_hd__mux2_8
XFILLER_88_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5248_ _5248_/A _5248_/B vssd1 vssd1 vccd1 vccd1 _5338_/B sky130_fd_sc_hd__nor2_8
XFILLER_68_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5179_ _5179_/A _5179_/B vssd1 vssd1 vccd1 vccd1 _5284_/A sky130_fd_sc_hd__xnor2_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4550_ _7285_/A _4920_/A _7281_/B _4456_/B vssd1 vssd1 vccd1 vccd1 _4551_/D sky130_fd_sc_hd__a22o_2
X_4481_ _4483_/A _6999_/A _4662_/A _4472_/A vssd1 vssd1 vccd1 vccd1 _4481_/X sky130_fd_sc_hd__a211o_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6220_ _7570_/B _6179_/X _6219_/X vssd1 vssd1 vccd1 vccd1 _6220_/Y sky130_fd_sc_hd__a21oi_1
X_6151_ _7319_/B _6139_/B _6127_/A _6146_/B _6150_/Y vssd1 vssd1 vccd1 vccd1 _6151_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5102_ _5198_/B _5530_/A vssd1 vssd1 vccd1 vccd1 _5187_/A sky130_fd_sc_hd__or2_4
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6081_/A _6081_/B _6088_/A vssd1 vssd1 vccd1 vccd1 _6110_/A sky130_fd_sc_hd__a21o_4
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5033_/A _5033_/B vssd1 vssd1 vccd1 vccd1 _5034_/C sky130_fd_sc_hd__nor2_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6984_ _6991_/B _6984_/B vssd1 vssd1 vccd1 vccd1 _6993_/B sky130_fd_sc_hd__or2_2
XFILLER_25_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5935_ _5876_/B _6241_/B _5874_/Y vssd1 vssd1 vccd1 vccd1 _6227_/B sky130_fd_sc_hd__a21o_4
XFILLER_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5866_ _5866_/A _5866_/B _5866_/C vssd1 vssd1 vccd1 vccd1 _5869_/A sky130_fd_sc_hd__or3_2
X_7605_ _7928_/A _7605_/B vssd1 vssd1 vccd1 vccd1 _8029_/D sky130_fd_sc_hd__nor2_1
X_4817_ _4854_/A _4817_/B vssd1 vssd1 vccd1 vccd1 _4826_/A sky130_fd_sc_hd__xnor2_1
XFILLER_21_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5797_ _5797_/A _5853_/B vssd1 vssd1 vccd1 vccd1 _5855_/C sky130_fd_sc_hd__or2_4
XFILLER_119_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7536_ _7889_/A _7542_/C _7543_/B _7543_/C vssd1 vssd1 vccd1 vccd1 _7536_/X sky130_fd_sc_hd__or4_1
X_4748_ _4832_/A _4748_/B vssd1 vssd1 vccd1 vccd1 _4850_/A sky130_fd_sc_hd__nor2_2
XFILLER_107_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7467_ _7403_/C _7403_/B _7502_/B vssd1 vssd1 vccd1 vccd1 _7467_/X sky130_fd_sc_hd__mux2_1
X_4679_ _4716_/A _4716_/B _4679_/C vssd1 vssd1 vccd1 vccd1 _4687_/A sky130_fd_sc_hd__and3_2
X_6418_ _6418_/A _6418_/B vssd1 vssd1 vccd1 vccd1 _6419_/B sky130_fd_sc_hd__nand2_1
X_7398_ _7398_/A _7398_/B vssd1 vssd1 vccd1 vccd1 _7403_/A sky130_fd_sc_hd__xnor2_4
XFILLER_102_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6349_ _6349_/A _6349_/B vssd1 vssd1 vccd1 vccd1 _6350_/B sky130_fd_sc_hd__and2_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8019_ _8075_/CLK _8019_/D vssd1 vssd1 vccd1 vccd1 _8019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5720_ _5720_/A _5720_/B vssd1 vssd1 vccd1 vccd1 _5763_/A sky130_fd_sc_hd__xnor2_4
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5651_ _5652_/B vssd1 vssd1 vccd1 vccd1 _5651_/Y sky130_fd_sc_hd__inv_2
X_5582_ _5582_/A _5683_/B vssd1 vssd1 vccd1 vccd1 _5639_/B sky130_fd_sc_hd__or2_4
X_4602_ _4602_/A _5013_/B vssd1 vssd1 vccd1 vccd1 _4604_/B sky130_fd_sc_hd__nor2_4
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7321_ _7326_/A _7326_/B vssd1 vssd1 vccd1 vccd1 _7321_/Y sky130_fd_sc_hd__nand2b_1
X_4533_ _6916_/A _7136_/A _4430_/A _5040_/A _4532_/X vssd1 vssd1 vccd1 vccd1 _4534_/B
+ sky130_fd_sc_hd__a41o_2
XFILLER_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7252_ _7252_/A _7252_/B vssd1 vssd1 vccd1 vccd1 _7256_/A sky130_fd_sc_hd__xnor2_4
XFILLER_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6203_ _7570_/B _6194_/X _6202_/X vssd1 vssd1 vccd1 vccd1 _6203_/Y sky130_fd_sc_hd__a21oi_1
X_4464_ _7165_/A _5020_/A _5040_/A _4430_/A vssd1 vssd1 vccd1 vccd1 _4465_/C sky130_fd_sc_hd__a22o_2
X_4395_ _4395_/A _4395_/B vssd1 vssd1 vccd1 vccd1 _4453_/A sky130_fd_sc_hd__xnor2_4
X_7183_ _7184_/A _7184_/B _7184_/C vssd1 vssd1 vccd1 vccd1 _7185_/A sky130_fd_sc_hd__a21oi_1
X_6134_ _6134_/A _6134_/B vssd1 vssd1 vccd1 vccd1 _6134_/X sky130_fd_sc_hd__or2_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _6065_/A _6065_/B vssd1 vssd1 vccd1 vccd1 _7426_/A sky130_fd_sc_hd__or2_2
XFILLER_97_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _5016_/A _5016_/B _5016_/C vssd1 vssd1 vccd1 vccd1 _5032_/A sky130_fd_sc_hd__and3_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6967_ _6967_/A _6967_/B vssd1 vssd1 vccd1 vccd1 _6977_/A sky130_fd_sc_hd__nor2_4
XFILLER_81_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5918_ _5918_/A _5918_/B vssd1 vssd1 vccd1 vccd1 _5919_/C sky130_fd_sc_hd__nor2_1
XFILLER_34_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6898_ _6999_/A _7195_/B vssd1 vssd1 vccd1 vccd1 _6943_/A sky130_fd_sc_hd__nand2_1
X_5849_ _5849_/A vssd1 vssd1 vccd1 vccd1 _6227_/A sky130_fd_sc_hd__inv_2
XFILLER_108_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7519_ _7366_/C _7365_/B _7367_/B _7367_/A vssd1 vssd1 vccd1 vccd1 _7519_/X sky130_fd_sc_hd__o211a_1
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4180_ _4228_/B vssd1 vssd1 vccd1 vccd1 _4180_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_95_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7870_ _7847_/A _7658_/Y _7766_/Y vssd1 vssd1 vccd1 vccd1 _7872_/B sky130_fd_sc_hd__o21bai_2
X_6821_ _6827_/B _6824_/A vssd1 vssd1 vccd1 vccd1 _6822_/B sky130_fd_sc_hd__nand2_2
XFILLER_35_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6752_ _6741_/X _6750_/X _6751_/X _6638_/A vssd1 vssd1 vccd1 vccd1 _6760_/A sky130_fd_sc_hd__o31a_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6683_ _6539_/A _6539_/B _6688_/S vssd1 vssd1 vccd1 vccd1 _6683_/X sky130_fd_sc_hd__mux2_1
X_5703_ _5703_/A _5703_/B vssd1 vssd1 vccd1 vccd1 _5908_/C sky130_fd_sc_hd__nand2_4
X_5634_ _5679_/A _5679_/B _5626_/X vssd1 vssd1 vccd1 vccd1 _5637_/A sky130_fd_sc_hd__a21o_4
XFILLER_117_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7304_ _7304_/A _7304_/B vssd1 vssd1 vccd1 vccd1 _7330_/A sky130_fd_sc_hd__or2_4
X_5565_ _5800_/A _5755_/A vssd1 vssd1 vccd1 vccd1 _5619_/A sky130_fd_sc_hd__nor2_4
XFILLER_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5496_ _5497_/A _5497_/B vssd1 vssd1 vccd1 vccd1 _5496_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4516_ _4516_/A _4516_/B _4795_/A vssd1 vssd1 vccd1 vccd1 _4517_/B sky130_fd_sc_hd__nand3_2
XFILLER_117_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7235_ _7294_/A _7235_/B vssd1 vssd1 vccd1 vccd1 _7239_/B sky130_fd_sc_hd__nor2_4
X_4447_ _6916_/A _4445_/X _4440_/X vssd1 vssd1 vccd1 vccd1 _4447_/Y sky130_fd_sc_hd__o21ai_4
X_7166_ _7205_/A _7205_/B vssd1 vssd1 vccd1 vccd1 _7177_/B sky130_fd_sc_hd__or2_4
XFILLER_98_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4378_ _7165_/A _4412_/B _4396_/B _4455_/A _4377_/A vssd1 vssd1 vccd1 vccd1 _4378_/X
+ sky130_fd_sc_hd__o2111a_1
X_6117_ _6118_/A _6118_/B vssd1 vssd1 vccd1 vccd1 _6117_/X sky130_fd_sc_hd__or2_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _7097_/A _7097_/B vssd1 vssd1 vccd1 vccd1 _7108_/B sky130_fd_sc_hd__xnor2_4
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6048_ _4548_/C _6047_/X _6048_/S vssd1 vssd1 vccd1 vccd1 _6054_/A sky130_fd_sc_hd__mux2_2
XFILLER_100_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7999_ _8074_/Q _8018_/Q _8004_/S vssd1 vssd1 vccd1 vccd1 _8074_/D sky130_fd_sc_hd__mux2_1
XFILLER_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5350_ _5530_/A _6971_/B vssd1 vssd1 vccd1 vccd1 _5354_/A sky130_fd_sc_hd__nor2_4
X_4301_ _4301_/A _4301_/B vssd1 vssd1 vccd1 vccd1 _4301_/Y sky130_fd_sc_hd__nand2_1
X_5281_ _5278_/Y _5281_/B vssd1 vssd1 vccd1 vccd1 _5492_/B sky130_fd_sc_hd__and2b_2
X_4232_ _4164_/X _4229_/X _4230_/X vssd1 vssd1 vccd1 vccd1 _4232_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_4_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7020_ _7015_/A _7015_/B _7007_/X vssd1 vssd1 vccd1 vccd1 _7022_/A sky130_fd_sc_hd__a21o_1
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4163_ _4158_/X _4159_/Y _4230_/C vssd1 vssd1 vccd1 vccd1 _4210_/A sky130_fd_sc_hd__a21oi_4
XFILLER_67_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4094_ _6326_/A _4094_/B vssd1 vssd1 vccd1 vccd1 _4095_/B sky130_fd_sc_hd__xor2_2
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7922_ _7935_/A _7900_/X _7921_/Y vssd1 vssd1 vccd1 vccd1 _7935_/B sky130_fd_sc_hd__a21o_1
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7853_ _6268_/X _7838_/Y _7839_/X _7852_/X vssd1 vssd1 vccd1 vccd1 _7853_/X sky130_fd_sc_hd__a31o_2
XFILLER_82_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7784_ _7784_/A _7784_/B vssd1 vssd1 vccd1 vccd1 _7833_/B sky130_fd_sc_hd__or2_4
X_6804_ _6804_/A _6804_/B vssd1 vssd1 vccd1 vccd1 _6815_/A sky130_fd_sc_hd__nand2_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4996_ _5001_/A _5001_/B vssd1 vssd1 vccd1 vccd1 _4996_/Y sky130_fd_sc_hd__nand2_1
X_6735_ _6728_/X _6734_/A _7581_/S vssd1 vssd1 vccd1 vccd1 _6735_/X sky130_fd_sc_hd__mux2_1
X_6666_ _6666_/A vssd1 vssd1 vccd1 vccd1 _6666_/Y sky130_fd_sc_hd__inv_2
X_6597_ _6605_/B _6612_/A _6605_/A vssd1 vssd1 vccd1 vccd1 _6617_/C sky130_fd_sc_hd__o21a_1
X_5617_ _5617_/A _5617_/B vssd1 vssd1 vccd1 vccd1 _5943_/A sky130_fd_sc_hd__nor2_4
X_5548_ _5548_/A _5548_/B vssd1 vssd1 vccd1 vccd1 _5560_/A sky130_fd_sc_hd__xor2_2
XFILLER_105_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5479_ _5613_/A _5480_/B vssd1 vssd1 vccd1 vccd1 _6147_/A sky130_fd_sc_hd__and2b_1
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7218_ _7219_/A _7219_/B vssd1 vssd1 vccd1 vccd1 _7218_/X sky130_fd_sc_hd__and2b_1
X_7149_ _7151_/B _7151_/A vssd1 vssd1 vccd1 vccd1 _7149_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_48_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout61 _6483_/A vssd1 vssd1 vccd1 vccd1 _6431_/S sky130_fd_sc_hd__clkbuf_8
Xfanout72 _5923_/A vssd1 vssd1 vccd1 vccd1 _7285_/B sky130_fd_sc_hd__buf_12
Xfanout50 _5364_/Y vssd1 vssd1 vccd1 vccd1 _5647_/B sky130_fd_sc_hd__buf_4
Xfanout83 _6873_/B vssd1 vssd1 vccd1 vccd1 _7269_/B sky130_fd_sc_hd__buf_12
Xfanout94 _4446_/X vssd1 vssd1 vccd1 vccd1 _4630_/B sky130_fd_sc_hd__buf_4
XFILLER_10_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_7__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _8082_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4850_ _4850_/A _4868_/D vssd1 vssd1 vccd1 vccd1 _4866_/A sky130_fd_sc_hd__xor2_2
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6520_ _6520_/A _6520_/B vssd1 vssd1 vccd1 vccd1 _6521_/A sky130_fd_sc_hd__xnor2_2
X_4781_ _4782_/B _4782_/A vssd1 vssd1 vccd1 vccd1 _4785_/B sky130_fd_sc_hd__and2b_1
XFILLER_119_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6451_ _6451_/A _6451_/B vssd1 vssd1 vccd1 vccd1 _6451_/Y sky130_fd_sc_hd__nand2_1
X_6382_ _6484_/S _6363_/C _6381_/X vssd1 vssd1 vccd1 vccd1 _6383_/B sky130_fd_sc_hd__o21ai_2
X_5402_ _5432_/A _5432_/B vssd1 vssd1 vccd1 vccd1 _5403_/B sky130_fd_sc_hd__xor2_4
X_5333_ _5335_/A _5335_/B vssd1 vssd1 vccd1 vccd1 _5333_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8052_ _8079_/CLK _8052_/D vssd1 vssd1 vccd1 vccd1 _8052_/Q sky130_fd_sc_hd__dfxtp_4
X_5264_ _5264_/A _5275_/A _5464_/B vssd1 vssd1 vccd1 vccd1 _5265_/B sky130_fd_sc_hd__or3_1
XFILLER_102_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4215_ _4221_/B _4215_/B vssd1 vssd1 vccd1 vccd1 _4215_/Y sky130_fd_sc_hd__nor2_1
X_5195_ _5196_/A _5196_/B vssd1 vssd1 vccd1 vccd1 _5195_/Y sky130_fd_sc_hd__nand2_1
X_7003_ _7306_/A _7007_/B _7000_/X vssd1 vssd1 vccd1 vccd1 _7056_/B sky130_fd_sc_hd__a21o_2
X_4146_ _8080_/Q _8079_/Q vssd1 vssd1 vccd1 vccd1 _4147_/D sky130_fd_sc_hd__or2_1
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4077_ _4087_/A _4077_/B vssd1 vssd1 vccd1 vccd1 _4078_/B sky130_fd_sc_hd__xor2_4
XFILLER_83_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7905_ _7903_/Y _7904_/X _7928_/A vssd1 vssd1 vccd1 vccd1 _8040_/D sky130_fd_sc_hd__o21ba_1
XFILLER_70_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7836_ _7883_/A _7836_/B vssd1 vssd1 vccd1 vccd1 _7839_/B sky130_fd_sc_hd__and2b_1
XFILLER_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7767_ _7766_/B _7551_/X _7766_/Y vssd1 vssd1 vccd1 vccd1 _7769_/B sky130_fd_sc_hd__a21o_1
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4979_ _4979_/A _4979_/B _4979_/C vssd1 vssd1 vccd1 vccd1 _5054_/C sky130_fd_sc_hd__and3_2
X_6718_ _6515_/B _6709_/A _6737_/B vssd1 vssd1 vccd1 vccd1 _6719_/A sky130_fd_sc_hd__mux2_1
X_7698_ _7639_/B _7571_/X _7639_/Y vssd1 vssd1 vccd1 vccd1 _7698_/X sky130_fd_sc_hd__o21a_1
X_6649_ _6647_/Y _6663_/B _6695_/S vssd1 vssd1 vccd1 vccd1 _6650_/B sky130_fd_sc_hd__mux2_1
XFILLER_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout240 _7952_/B1 vssd1 vssd1 vccd1 vccd1 _7903_/B1 sky130_fd_sc_hd__buf_6
XFILLER_78_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5951_ _5951_/A _5951_/B _5951_/C vssd1 vssd1 vccd1 vccd1 _6173_/B sky130_fd_sc_hd__and3_1
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4902_ _5040_/B _4902_/B vssd1 vssd1 vccd1 vccd1 _4938_/A sky130_fd_sc_hd__xor2_2
XFILLER_45_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5882_ _7306_/B _5858_/B _5859_/A vssd1 vssd1 vccd1 vccd1 _5884_/B sky130_fd_sc_hd__a21boi_1
X_7621_ _7622_/A _7622_/B _7648_/C vssd1 vssd1 vccd1 vccd1 _7621_/Y sky130_fd_sc_hd__o21ai_1
X_4833_ _4833_/A _4833_/B vssd1 vssd1 vccd1 vccd1 _4860_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7552_ _7495_/Y _7551_/X _7889_/A vssd1 vssd1 vccd1 vccd1 _7554_/C sky130_fd_sc_hd__mux2_2
XFILLER_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4764_ _5095_/A _4764_/B vssd1 vssd1 vccd1 vccd1 _4766_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6503_ _6543_/A _6502_/Y _6478_/X vssd1 vssd1 vccd1 vccd1 _6503_/Y sky130_fd_sc_hd__a21oi_4
X_7483_ _7479_/X _7441_/X _7483_/S vssd1 vssd1 vccd1 vccd1 _7483_/X sky130_fd_sc_hd__mux2_1
X_6434_ _6374_/A _6441_/S _6354_/X _6433_/X vssd1 vssd1 vccd1 vccd1 _6437_/A sky130_fd_sc_hd__a31o_1
X_4695_ _4648_/B _4650_/B _4693_/X _4606_/Y vssd1 vssd1 vccd1 vccd1 _4695_/X sky130_fd_sc_hd__a211o_2
X_6365_ _6969_/A _6806_/A _6456_/S vssd1 vssd1 vccd1 vccd1 _6468_/B sky130_fd_sc_hd__mux2_4
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6296_ _6296_/A _6296_/B vssd1 vssd1 vccd1 vccd1 _6296_/X sky130_fd_sc_hd__and2_2
X_5316_ _7213_/A _5977_/B _5977_/C _5977_/D vssd1 vssd1 vccd1 vccd1 _5316_/Y sky130_fd_sc_hd__nand4_4
XFILLER_114_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8035_ _8082_/CLK _8035_/D vssd1 vssd1 vccd1 vccd1 _8035_/Q sky130_fd_sc_hd__dfxtp_1
X_5247_ _5247_/A _5247_/B _5247_/C vssd1 vssd1 vccd1 vccd1 _5248_/B sky130_fd_sc_hd__and3_2
XFILLER_102_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5178_ _5181_/A _5178_/B vssd1 vssd1 vccd1 vccd1 _5179_/B sky130_fd_sc_hd__xnor2_2
XFILLER_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4129_ _5977_/B _4124_/X _4125_/X _4128_/X vssd1 vssd1 vccd1 vccd1 _7170_/B sky130_fd_sc_hd__a31o_4
XFILLER_56_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7819_ _7814_/X _7874_/C _7818_/Y vssd1 vssd1 vccd1 vccd1 _7819_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4480_ _4413_/X _4475_/X _4436_/A vssd1 vssd1 vccd1 vccd1 _4480_/X sky130_fd_sc_hd__a21o_1
X_6150_ _6242_/S _6150_/B vssd1 vssd1 vccd1 vccd1 _6150_/Y sky130_fd_sc_hd__nand2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5530_/A vssd1 vssd1 vccd1 vccd1 _5174_/B sky130_fd_sc_hd__inv_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6081_/A _6081_/B vssd1 vssd1 vccd1 vccd1 _6081_/Y sky130_fd_sc_hd__nand2_4
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5032_ _5032_/A _5032_/B vssd1 vssd1 vccd1 vccd1 _5038_/A sky130_fd_sc_hd__nor2_1
XFILLER_38_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6983_ _6983_/A _6983_/B _6995_/A vssd1 vssd1 vccd1 vccd1 _6984_/B sky130_fd_sc_hd__and3_1
XFILLER_15_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5934_ _5897_/Y _5932_/X _5933_/B vssd1 vssd1 vccd1 vccd1 _6241_/B sky130_fd_sc_hd__a21bo_1
XFILLER_80_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5865_ _5885_/A _5862_/A _5864_/Y _5863_/Y vssd1 vssd1 vccd1 vccd1 _5866_/C sky130_fd_sc_hd__o31a_1
X_7604_ _8029_/Q _7857_/B _7603_/X vssd1 vssd1 vccd1 vccd1 _7605_/B sky130_fd_sc_hd__a21oi_1
X_4816_ _4816_/A _4816_/B vssd1 vssd1 vccd1 vccd1 _4829_/A sky130_fd_sc_hd__nor2_2
XFILLER_119_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5796_ _6971_/B _5796_/B vssd1 vssd1 vccd1 vccd1 _5798_/C sky130_fd_sc_hd__nor2_1
X_7535_ _7535_/A _7535_/B vssd1 vssd1 vccd1 vccd1 _7543_/C sky130_fd_sc_hd__and2_1
X_4747_ _4868_/B _4775_/A _4746_/A vssd1 vssd1 vccd1 vccd1 _4748_/B sky130_fd_sc_hd__a21oi_2
XFILLER_119_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7466_ _7455_/X _7403_/D _7502_/B vssd1 vssd1 vccd1 vccd1 _7466_/X sky130_fd_sc_hd__mux2_1
X_4678_ _4716_/A _4716_/B vssd1 vssd1 vccd1 vccd1 _4717_/A sky130_fd_sc_hd__nand2_1
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7397_ _6005_/Y _7400_/B _6006_/X vssd1 vssd1 vccd1 vccd1 _7398_/B sky130_fd_sc_hd__a21o_4
X_6417_ _6418_/A _6418_/B vssd1 vssd1 vccd1 vccd1 _6417_/X sky130_fd_sc_hd__and2_1
XFILLER_115_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6348_ _7401_/A _6348_/B vssd1 vssd1 vccd1 vccd1 _6492_/B sky130_fd_sc_hd__xor2_4
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6279_ _4098_/B _4200_/B _6276_/X _6277_/X _6278_/X vssd1 vssd1 vccd1 vccd1 _6279_/X
+ sky130_fd_sc_hd__o221a_1
X_8018_ _8057_/CLK _8018_/D vssd1 vssd1 vccd1 vccd1 _8018_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_56_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
X_5650_ _5650_/A _5650_/B vssd1 vssd1 vccd1 vccd1 _5652_/B sky130_fd_sc_hd__and2_4
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4601_ _4594_/A _4594_/B _4594_/C vssd1 vssd1 vccd1 vccd1 _4604_/A sky130_fd_sc_hd__a21bo_4
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5581_ _5683_/A _5683_/B vssd1 vssd1 vccd1 vccd1 _5684_/A sky130_fd_sc_hd__nor2_2
XFILLER_30_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7320_ _7320_/A _7328_/A vssd1 vssd1 vccd1 vccd1 _7326_/B sky130_fd_sc_hd__xnor2_4
X_4532_ _4602_/A _4558_/B _4440_/X vssd1 vssd1 vccd1 vccd1 _4532_/X sky130_fd_sc_hd__o21a_1
X_7251_ _7251_/A _7251_/B vssd1 vssd1 vccd1 vccd1 _7252_/B sky130_fd_sc_hd__xnor2_4
X_4463_ _4602_/A _7116_/A _4988_/A _4630_/B vssd1 vssd1 vccd1 vccd1 _4516_/A sky130_fd_sc_hd__or4_4
X_6202_ _6199_/S _6149_/X _6189_/X _6219_/A vssd1 vssd1 vccd1 vccd1 _6202_/X sky130_fd_sc_hd__o211a_1
XFILLER_98_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4394_ _4395_/B _4395_/A vssd1 vssd1 vccd1 vccd1 _4394_/Y sky130_fd_sc_hd__nand2b_2
X_7182_ _7182_/A _7182_/B vssd1 vssd1 vccd1 vccd1 _7184_/C sky130_fd_sc_hd__xnor2_2
XFILLER_112_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6133_ _6134_/A _6134_/B vssd1 vssd1 vccd1 vccd1 _6225_/S sky130_fd_sc_hd__nor2_8
XFILLER_58_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6064_ _6065_/A _6065_/B vssd1 vssd1 vccd1 vccd1 _6064_/Y sky130_fd_sc_hd__nor2_2
XFILLER_97_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5013_/B _5013_/C _5040_/B _4947_/A vssd1 vssd1 vccd1 vccd1 _5016_/C sky130_fd_sc_hd__a2bb2o_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6966_ _6966_/A _6966_/B vssd1 vssd1 vccd1 vccd1 _6967_/B sky130_fd_sc_hd__and2_1
XFILLER_53_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5917_ _5917_/A _5922_/A vssd1 vssd1 vccd1 vccd1 _5918_/B sky130_fd_sc_hd__nor2_1
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6897_ _6947_/C _6897_/B vssd1 vssd1 vccd1 vccd1 _6909_/B sky130_fd_sc_hd__xor2_1
XFILLER_22_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5848_ _5848_/A _5848_/B vssd1 vssd1 vccd1 vccd1 _5849_/A sky130_fd_sc_hd__xnor2_1
X_5779_ _5779_/A _5779_/B vssd1 vssd1 vccd1 vccd1 _5781_/B sky130_fd_sc_hd__xor2_4
X_7518_ _7371_/A _7371_/B _7371_/C vssd1 vssd1 vccd1 vccd1 _7518_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7449_ _7445_/Y _7448_/Y _7479_/S vssd1 vssd1 vccd1 vccd1 _7449_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6820_ _6820_/A _6820_/B vssd1 vssd1 vccd1 vccd1 _6824_/B sky130_fd_sc_hd__xnor2_4
XFILLER_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6751_ _6740_/X _6656_/X _6751_/S vssd1 vssd1 vccd1 vccd1 _6751_/X sky130_fd_sc_hd__mux2_1
X_6682_ _6739_/S _6662_/X _6681_/Y vssd1 vssd1 vccd1 vccd1 _6704_/B sky130_fd_sc_hd__o21ai_1
X_5702_ _5706_/A _5706_/B vssd1 vssd1 vccd1 vccd1 _5702_/Y sky130_fd_sc_hd__nor2_1
X_5633_ _5633_/A _5633_/B vssd1 vssd1 vccd1 vccd1 _5679_/B sky130_fd_sc_hd__xnor2_4
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5564_ _7150_/B _5880_/A vssd1 vssd1 vccd1 vccd1 _5566_/B sky130_fd_sc_hd__nor2_8
XFILLER_117_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7303_ _7334_/B _7294_/B _7344_/B _4354_/X vssd1 vssd1 vccd1 vccd1 _7304_/B sky130_fd_sc_hd__o22a_1
X_4515_ _4516_/A _4516_/B _4795_/A vssd1 vssd1 vccd1 vccd1 _4517_/A sky130_fd_sc_hd__a21o_2
X_5495_ _5495_/A _5495_/B vssd1 vssd1 vccd1 vccd1 _5497_/B sky130_fd_sc_hd__xor2_4
XFILLER_104_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7234_ _7234_/A _7234_/B vssd1 vssd1 vccd1 vccd1 _7239_/A sky130_fd_sc_hd__xor2_4
X_4446_ _6916_/A _4445_/X _4440_/X vssd1 vssd1 vccd1 vccd1 _4446_/X sky130_fd_sc_hd__o21a_2
X_7165_ _7165_/A _7281_/D vssd1 vssd1 vccd1 vccd1 _7205_/B sky130_fd_sc_hd__nand2_2
X_4377_ _4377_/A _4455_/A _4396_/B vssd1 vssd1 vccd1 vccd1 _4377_/X sky130_fd_sc_hd__and3_1
XFILLER_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _5940_/X _5944_/Y _5710_/X vssd1 vssd1 vccd1 vccd1 _6118_/B sky130_fd_sc_hd__a21oi_2
XFILLER_112_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _7090_/A _7090_/B _7082_/A vssd1 vssd1 vccd1 vccd1 _7108_/A sky130_fd_sc_hd__o21ba_4
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6047_ _6272_/B _6274_/B _4547_/C vssd1 vssd1 vccd1 vccd1 _6047_/X sky130_fd_sc_hd__a21o_2
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7998_ _8073_/Q _8017_/Q _8007_/S vssd1 vssd1 vccd1 vccd1 _8073_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6949_ _6903_/A _7067_/A _6948_/X vssd1 vssd1 vccd1 vccd1 _6957_/A sky130_fd_sc_hd__o21ba_1
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4300_ _4062_/B _5993_/B _4297_/X _4303_/B vssd1 vssd1 vccd1 vccd1 _4301_/B sky130_fd_sc_hd__a211o_1
X_5280_ _5280_/A _5280_/B vssd1 vssd1 vccd1 vccd1 _5281_/B sky130_fd_sc_hd__nand2_2
XFILLER_5_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4231_ _4164_/X _4229_/X _4230_/X vssd1 vssd1 vccd1 vccd1 _4231_/X sky130_fd_sc_hd__o21a_2
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4162_ _4216_/B _6273_/B vssd1 vssd1 vccd1 vccd1 _4230_/C sky130_fd_sc_hd__xor2_4
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4093_ _8056_/Q _4093_/B vssd1 vssd1 vccd1 vccd1 _4094_/B sky130_fd_sc_hd__xnor2_4
X_7921_ _7921_/A _7921_/B vssd1 vssd1 vccd1 vccd1 _7921_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_95_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7852_ _7844_/Y _7845_/X _7851_/X _7952_/B1 vssd1 vssd1 vccd1 vccd1 _7852_/X sky130_fd_sc_hd__a211o_1
XFILLER_51_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7783_ _7759_/Y _7760_/X _6522_/S vssd1 vssd1 vccd1 vccd1 _7787_/A sky130_fd_sc_hd__o21a_1
XFILLER_91_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6803_ _6834_/A _6834_/B _6834_/C vssd1 vssd1 vccd1 vccd1 _6835_/A sky130_fd_sc_hd__o21a_1
X_4995_ _4995_/A _4995_/B vssd1 vssd1 vccd1 vccd1 _5001_/B sky130_fd_sc_hd__xor2_4
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6734_ _6734_/A vssd1 vssd1 vccd1 vccd1 _6734_/Y sky130_fd_sc_hd__inv_2
X_6665_ _6537_/Y _6547_/A _6688_/S vssd1 vssd1 vccd1 vccd1 _6666_/A sky130_fd_sc_hd__mux2_1
X_6596_ _6611_/A _6611_/B vssd1 vssd1 vccd1 vccd1 _6612_/A sky130_fd_sc_hd__nor2_1
X_5616_ _5616_/A _5616_/B _5616_/C vssd1 vssd1 vccd1 vccd1 _5617_/B sky130_fd_sc_hd__and3_1
X_5547_ _5547_/A _5547_/B vssd1 vssd1 vccd1 vccd1 _5548_/B sky130_fd_sc_hd__xnor2_4
XFILLER_117_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5478_ _5491_/A _5478_/B vssd1 vssd1 vccd1 vccd1 _5480_/B sky130_fd_sc_hd__and2_1
X_4429_ _4362_/X _4429_/B vssd1 vssd1 vccd1 vccd1 _4429_/X sky130_fd_sc_hd__and2b_1
X_7217_ _7251_/A _7251_/B _7214_/X vssd1 vssd1 vccd1 vccd1 _7219_/B sky130_fd_sc_hd__a21bo_1
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7148_ _7094_/B _7109_/X _7146_/B _7147_/Y vssd1 vssd1 vccd1 vccd1 _7151_/B sky130_fd_sc_hd__o31a_4
XFILLER_100_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7079_ _7079_/A _7079_/B vssd1 vssd1 vccd1 vccd1 _7081_/C sky130_fd_sc_hd__xnor2_2
XFILLER_100_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout40 _5273_/A vssd1 vssd1 vccd1 vccd1 _5386_/A sky130_fd_sc_hd__buf_8
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout62 _6347_/Y vssd1 vssd1 vccd1 vccd1 _6492_/A sky130_fd_sc_hd__buf_4
Xfanout51 _5344_/B vssd1 vssd1 vccd1 vccd1 _5755_/A sky130_fd_sc_hd__buf_12
Xfanout73 _7247_/D vssd1 vssd1 vccd1 vccd1 _6971_/B sky130_fd_sc_hd__buf_6
XFILLER_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout95 _4426_/X vssd1 vssd1 vccd1 vccd1 _5013_/A sky130_fd_sc_hd__buf_6
Xfanout84 _5137_/X vssd1 vssd1 vccd1 vccd1 _7235_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4780_ _4854_/A _4779_/B _4779_/A vssd1 vssd1 vccd1 vccd1 _4782_/B sky130_fd_sc_hd__o21ba_1
XFILLER_21_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6450_ _6483_/A _6438_/X _6449_/Y vssd1 vssd1 vccd1 vccd1 _6450_/Y sky130_fd_sc_hd__o21ai_1
X_6381_ _6451_/A _6381_/B vssd1 vssd1 vccd1 vccd1 _6381_/X sky130_fd_sc_hd__or2_1
X_5401_ _5401_/A _5401_/B vssd1 vssd1 vccd1 vccd1 _5432_/B sky130_fd_sc_hd__xnor2_4
X_5332_ _5332_/A _5332_/B vssd1 vssd1 vccd1 vccd1 _5335_/B sky130_fd_sc_hd__xor2_4
XFILLER_114_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8051_ _8075_/CLK _8051_/D vssd1 vssd1 vccd1 vccd1 _8051_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5263_ _5258_/A _5258_/B _5256_/Y vssd1 vssd1 vccd1 vccd1 _5267_/A sky130_fd_sc_hd__a21boi_4
X_4214_ _4228_/A _4216_/C vssd1 vssd1 vccd1 vccd1 _4215_/B sky130_fd_sc_hd__or2_1
X_7002_ _7306_/A _7007_/B vssd1 vssd1 vccd1 vccd1 _7008_/A sky130_fd_sc_hd__nand2_2
X_5194_ _5259_/A _5259_/B vssd1 vssd1 vccd1 vccd1 _5196_/B sky130_fd_sc_hd__and2b_4
X_4145_ _8078_/Q _8076_/Q _8075_/Q _8077_/Q vssd1 vssd1 vccd1 vccd1 _4147_/C sky130_fd_sc_hd__or4_4
XFILLER_68_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4076_ _8062_/Q _4076_/B vssd1 vssd1 vccd1 vccd1 _4077_/B sky130_fd_sc_hd__xnor2_4
XFILLER_83_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7904_ _8039_/Q _4018_/X _7857_/B _8040_/Q vssd1 vssd1 vccd1 vccd1 _7904_/X sky130_fd_sc_hd__a22o_1
XFILLER_71_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7835_ _7833_/A _7833_/B _7833_/C _7834_/Y vssd1 vssd1 vccd1 vccd1 _7836_/B sky130_fd_sc_hd__a31o_1
XFILLER_24_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7766_ _7766_/A _7766_/B vssd1 vssd1 vccd1 vccd1 _7766_/Y sky130_fd_sc_hd__nor2_4
XFILLER_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4978_ _4979_/A _4979_/B _4979_/C vssd1 vssd1 vccd1 vccd1 _4978_/X sky130_fd_sc_hd__a21o_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6717_ _6638_/Y _6703_/X _6707_/X _7616_/S _6716_/X vssd1 vssd1 vccd1 vccd1 _6732_/B
+ sky130_fd_sc_hd__a221o_1
X_7697_ _7760_/A _7697_/B vssd1 vssd1 vccd1 vccd1 _7697_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6648_ _6581_/A _6570_/Y _6737_/B vssd1 vssd1 vccd1 vccd1 _6663_/B sky130_fd_sc_hd__mux2_1
XFILLER_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6579_ _6594_/A _6594_/B vssd1 vssd1 vccd1 vccd1 _6605_/B sky130_fd_sc_hd__nor2_1
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout230 _8082_/Q vssd1 vssd1 vccd1 vccd1 _6770_/A sky130_fd_sc_hd__buf_8
Xfanout241 input1/X vssd1 vssd1 vccd1 vccd1 _7952_/B1 sky130_fd_sc_hd__buf_4
XFILLER_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5950_ _5502_/A _5948_/Y _5949_/X vssd1 vssd1 vccd1 vccd1 _5951_/C sky130_fd_sc_hd__o21a_1
XFILLER_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4901_ _5040_/B _4902_/B vssd1 vssd1 vccd1 vccd1 _4901_/Y sky130_fd_sc_hd__nand2_1
X_7620_ _7620_/A _7620_/B vssd1 vssd1 vccd1 vccd1 _7648_/C sky130_fd_sc_hd__xor2_2
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5881_ _5881_/A _5919_/A _5925_/A _5881_/D vssd1 vssd1 vccd1 vccd1 _5927_/C sky130_fd_sc_hd__or4_2
X_4832_ _4832_/A _4832_/B vssd1 vssd1 vccd1 vccd1 _4833_/B sky130_fd_sc_hd__and2_1
XFILLER_33_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7551_ _7500_/Y _7550_/X _7657_/B vssd1 vssd1 vccd1 vccd1 _7551_/X sky130_fd_sc_hd__mux2_1
X_4763_ _4763_/A _4763_/B vssd1 vssd1 vccd1 vccd1 _4764_/B sky130_fd_sc_hd__nand2_1
X_6502_ _6545_/A _6500_/Y _6501_/X vssd1 vssd1 vccd1 vccd1 _6502_/Y sky130_fd_sc_hd__o21ai_4
X_7482_ _7451_/X _7481_/X _7538_/S vssd1 vssd1 vccd1 vccd1 _7544_/A sky130_fd_sc_hd__mux2_1
X_4694_ _4648_/B _4650_/B _4693_/X _4606_/Y vssd1 vssd1 vccd1 vccd1 _4697_/B sky130_fd_sc_hd__a211oi_2
X_6433_ _6488_/A _6391_/Y _6432_/X _6492_/A _6443_/A vssd1 vssd1 vccd1 vccd1 _6433_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6364_ _6364_/A _6443_/B vssd1 vssd1 vccd1 vccd1 _6468_/A sky130_fd_sc_hd__nand2_1
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6295_ _6272_/B _4259_/B _6017_/A vssd1 vssd1 vccd1 vccd1 _6296_/B sky130_fd_sc_hd__a21o_1
X_5315_ _7213_/A _5977_/B _5977_/C _5977_/D vssd1 vssd1 vccd1 vccd1 _5315_/X sky130_fd_sc_hd__and4_1
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8034_ _8082_/CLK _8034_/D vssd1 vssd1 vccd1 vccd1 _8034_/Q sky130_fd_sc_hd__dfxtp_1
X_5246_ _5245_/A _5245_/B _5437_/A _5437_/B vssd1 vssd1 vccd1 vccd1 _5258_/A sky130_fd_sc_hd__a22o_4
XFILLER_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5177_ _5180_/A _5180_/B _5178_/B vssd1 vssd1 vccd1 vccd1 _5177_/X sky130_fd_sc_hd__and3_1
XFILLER_110_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4128_ _4088_/A _4303_/C _4126_/X _5268_/A _5135_/C1 vssd1 vssd1 vccd1 vccd1 _4128_/X
+ sky130_fd_sc_hd__o2111a_1
X_4059_ _6272_/A _4059_/B vssd1 vssd1 vccd1 vccd1 _4063_/A sky130_fd_sc_hd__xnor2_4
XFILLER_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7818_ _7814_/X _7874_/C _7802_/B2 vssd1 vssd1 vccd1 vccd1 _7818_/Y sky130_fd_sc_hd__o21bai_1
X_7749_ _7749_/A _7749_/B vssd1 vssd1 vccd1 vccd1 _7764_/B sky130_fd_sc_hd__xnor2_2
XFILLER_12_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6080_ _6081_/A _6081_/B vssd1 vssd1 vccd1 vccd1 _6259_/A sky130_fd_sc_hd__and2_1
X_5100_ _5100_/A _5100_/B vssd1 vssd1 vccd1 vccd1 _5244_/A sky130_fd_sc_hd__xor2_4
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5031_ _5016_/A _5016_/C _5016_/B vssd1 vssd1 vccd1 vccd1 _5032_/B sky130_fd_sc_hd__a21oi_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6982_ _6977_/A _6977_/B _6967_/A vssd1 vssd1 vccd1 vccd1 _6993_/A sky130_fd_sc_hd__a21o_2
XFILLER_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5933_ _5932_/X _5933_/B vssd1 vssd1 vccd1 vccd1 _6239_/B sky130_fd_sc_hd__and2b_1
XFILLER_80_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5864_ _6971_/B _5925_/B vssd1 vssd1 vccd1 vccd1 _5864_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7603_ _7578_/X _7600_/Y _7601_/X _7602_/X vssd1 vssd1 vccd1 vccd1 _7603_/X sky130_fd_sc_hd__o31a_1
X_4815_ _4832_/A _4815_/B vssd1 vssd1 vccd1 vccd1 _4816_/B sky130_fd_sc_hd__and2_1
XFILLER_21_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7534_ _7538_/S _7534_/B vssd1 vssd1 vccd1 vccd1 _7543_/B sky130_fd_sc_hd__and2_1
X_5795_ _5795_/A _5826_/A vssd1 vssd1 vccd1 vccd1 _5836_/A sky130_fd_sc_hd__xor2_2
X_4746_ _4746_/A _4868_/B _4775_/A vssd1 vssd1 vccd1 vccd1 _4832_/A sky130_fd_sc_hd__and3_4
XFILLER_119_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7465_ _7464_/X _7463_/X _7624_/S vssd1 vssd1 vccd1 vccd1 _7465_/X sky130_fd_sc_hd__mux2_1
X_4677_ _7214_/A _5013_/B vssd1 vssd1 vccd1 vccd1 _4679_/C sky130_fd_sc_hd__nor2_1
X_7396_ _7401_/A _7401_/B _6309_/Y vssd1 vssd1 vccd1 vccd1 _7400_/B sky130_fd_sc_hd__a21o_2
X_6416_ _6418_/A _6418_/B vssd1 vssd1 vccd1 vccd1 _6419_/A sky130_fd_sc_hd__or2_2
X_6347_ _6488_/A _6359_/A vssd1 vssd1 vccd1 vccd1 _6347_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6278_ _6278_/A _6278_/B vssd1 vssd1 vccd1 vccd1 _6278_/X sky130_fd_sc_hd__or2_1
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8017_ _8080_/CLK _8017_/D vssd1 vssd1 vccd1 vccd1 _8017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5229_ _5230_/A _5957_/A _5229_/C vssd1 vssd1 vccd1 vccd1 _5959_/A sky130_fd_sc_hd__or3_1
XFILLER_69_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4600_ _4599_/A _4599_/C _4599_/B vssd1 vssd1 vccd1 vccd1 _4606_/B sky130_fd_sc_hd__a21oi_4
X_5580_ _5580_/A _5580_/B vssd1 vssd1 vccd1 vccd1 _5643_/A sky130_fd_sc_hd__nor2_4
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4531_ _4773_/A _5033_/A vssd1 vssd1 vccd1 vccd1 _4795_/B sky130_fd_sc_hd__or2_4
X_7250_ _7257_/A _7257_/B vssd1 vssd1 vccd1 vccd1 _7250_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4462_ _7136_/A _5033_/A vssd1 vssd1 vccd1 vccd1 _4465_/A sky130_fd_sc_hd__nor2_2
X_6201_ _6193_/A _6199_/X _6200_/X vssd1 vssd1 vccd1 vccd1 _6250_/A sky130_fd_sc_hd__a21oi_2
X_7181_ _7181_/A _7181_/B vssd1 vssd1 vccd1 vccd1 _7203_/A sky130_fd_sc_hd__xor2_4
X_4393_ _4393_/A _4393_/B vssd1 vssd1 vccd1 vccd1 _4395_/B sky130_fd_sc_hd__xnor2_4
X_6132_ _6132_/A _6132_/B vssd1 vssd1 vccd1 vccd1 _6134_/B sky130_fd_sc_hd__xnor2_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6063_ _6326_/A _6951_/D _6015_/C vssd1 vssd1 vccd1 vccd1 _6065_/B sky130_fd_sc_hd__a21oi_4
XFILLER_58_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5014_ _5014_/A _5033_/B vssd1 vssd1 vccd1 vccd1 _5016_/B sky130_fd_sc_hd__nor2_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _6966_/A _6966_/B vssd1 vssd1 vccd1 vccd1 _6967_/A sky130_fd_sc_hd__nor2_2
X_5916_ _5916_/A _5916_/B vssd1 vssd1 vccd1 vccd1 _6236_/A sky130_fd_sc_hd__nand2_1
X_6896_ _6896_/A _6896_/B vssd1 vssd1 vccd1 vccd1 _6931_/A sky130_fd_sc_hd__xnor2_1
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5847_ _5847_/A _5847_/B vssd1 vssd1 vccd1 vccd1 _5847_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5778_ _5777_/A _5777_/B _5808_/B _5808_/A vssd1 vssd1 vccd1 vccd1 _5781_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7517_ _7517_/A _7517_/B vssd1 vssd1 vccd1 vccd1 _7517_/Y sky130_fd_sc_hd__nor2_1
X_4729_ _4728_/B _4728_/C _4720_/X vssd1 vssd1 vccd1 vccd1 _4730_/B sky130_fd_sc_hd__a21o_1
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7448_ _7448_/A _7448_/B vssd1 vssd1 vccd1 vccd1 _7448_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7379_ _7471_/A _7471_/B _7273_/A vssd1 vssd1 vccd1 vccd1 _7472_/B sky130_fd_sc_hd__o21ai_4
XFILLER_107_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6750_ _6657_/X _6675_/X _6703_/X _6707_/X _6749_/S vssd1 vssd1 vccd1 vccd1 _6750_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5701_ _5743_/A _5743_/B _5698_/Y vssd1 vssd1 vccd1 vccd1 _5706_/B sky130_fd_sc_hd__a21boi_4
X_6681_ _6713_/S _6681_/B vssd1 vssd1 vccd1 vccd1 _6681_/Y sky130_fd_sc_hd__nand2_1
X_5632_ _5632_/A _5632_/B vssd1 vssd1 vccd1 vccd1 _5633_/B sky130_fd_sc_hd__xnor2_4
XFILLER_31_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5563_ _5563_/A _5563_/B vssd1 vssd1 vccd1 vccd1 _5569_/B sky130_fd_sc_hd__xnor2_1
X_7302_ _7302_/A _7302_/B vssd1 vssd1 vccd1 vccd1 _7316_/A sky130_fd_sc_hd__xor2_4
X_4514_ _5445_/A _4642_/B vssd1 vssd1 vccd1 vccd1 _4795_/A sky130_fd_sc_hd__or2_4
X_5494_ _5495_/A _5495_/B vssd1 vssd1 vccd1 vccd1 _5499_/A sky130_fd_sc_hd__or2_4
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4445_ _4360_/A _4443_/Y _4444_/X _4404_/Y vssd1 vssd1 vccd1 vccd1 _4445_/X sky130_fd_sc_hd__o22a_2
X_7233_ _7240_/A _7240_/B _7231_/Y vssd1 vssd1 vccd1 vccd1 _7234_/B sky130_fd_sc_hd__a21boi_4
X_4376_ _4376_/A _4376_/B _4376_/C vssd1 vssd1 vccd1 vccd1 _4396_/B sky130_fd_sc_hd__or3_4
X_7164_ _7072_/B _7162_/Y _7169_/A vssd1 vssd1 vccd1 vccd1 _7205_/A sky130_fd_sc_hd__a21o_1
XFILLER_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6115_ _6115_/A _6115_/B vssd1 vssd1 vccd1 vccd1 _6115_/X sky130_fd_sc_hd__xor2_4
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7097_/B _7097_/A vssd1 vssd1 vccd1 vccd1 _7099_/A sky130_fd_sc_hd__nand2b_1
X_6046_ _6034_/A _6017_/A _4260_/C _6272_/B vssd1 vssd1 vccd1 vccd1 _6048_/S sky130_fd_sc_hd__a31o_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7997_ _8072_/Q _8016_/Q _8007_/S vssd1 vssd1 vccd1 vccd1 _8072_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6948_ _7101_/A _6902_/A _5137_/X _7012_/A vssd1 vssd1 vccd1 vccd1 _6948_/X sky130_fd_sc_hd__o22a_1
X_6879_ _6877_/A _6877_/B _6912_/A vssd1 vssd1 vccd1 vccd1 _6881_/B sky130_fd_sc_hd__o21ba_1
XFILLER_6_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4230_ _4230_/A _4230_/B _4230_/C vssd1 vssd1 vccd1 vccd1 _4230_/X sky130_fd_sc_hd__or3_4
X_4161_ _8080_/Q _4161_/B vssd1 vssd1 vccd1 vccd1 _6273_/B sky130_fd_sc_hd__xnor2_4
XFILLER_95_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4092_ _8055_/Q _4096_/B _4096_/A vssd1 vssd1 vccd1 vccd1 _4093_/B sky130_fd_sc_hd__o21ai_4
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7920_ _7920_/A _7921_/B vssd1 vssd1 vccd1 vccd1 _7920_/X sky130_fd_sc_hd__or2_1
X_7851_ _7846_/X _7874_/D _7850_/Y vssd1 vssd1 vccd1 vccd1 _7851_/X sky130_fd_sc_hd__o21a_1
XFILLER_82_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6802_ _6804_/B _6802_/B vssd1 vssd1 vccd1 vccd1 _6834_/C sky130_fd_sc_hd__and2_1
X_7782_ _7780_/X _7781_/Y _7856_/A vssd1 vssd1 vccd1 vccd1 _8035_/D sky130_fd_sc_hd__a21oi_1
XFILLER_51_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4994_ _5011_/A _5011_/B _4987_/Y vssd1 vssd1 vccd1 vccd1 _5001_/A sky130_fd_sc_hd__o21ai_4
X_6733_ _6616_/D _6616_/C _6733_/S vssd1 vssd1 vccd1 vccd1 _6734_/A sky130_fd_sc_hd__mux2_1
X_6664_ _6691_/B vssd1 vssd1 vccd1 vccd1 _6664_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5615_ _6118_/A _6123_/A vssd1 vssd1 vccd1 vccd1 _5615_/Y sky130_fd_sc_hd__nor2_2
X_6595_ _6605_/B _6595_/B vssd1 vssd1 vccd1 vccd1 _6611_/B sky130_fd_sc_hd__or2_1
X_5546_ _5547_/A _5547_/B vssd1 vssd1 vccd1 vccd1 _5546_/Y sky130_fd_sc_hd__nand2_1
X_5477_ _5477_/A _5477_/B _5477_/C vssd1 vssd1 vccd1 vccd1 _5478_/B sky130_fd_sc_hd__nand3_1
X_7216_ _7216_/A _7285_/C vssd1 vssd1 vccd1 vccd1 _7251_/B sky130_fd_sc_hd__xnor2_4
X_4428_ _4602_/A _5033_/A vssd1 vssd1 vccd1 vccd1 _4451_/A sky130_fd_sc_hd__nor2_2
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7147_ _7157_/A _7157_/B vssd1 vssd1 vccd1 vccd1 _7147_/Y sky130_fd_sc_hd__nand2_1
X_4359_ _7165_/A _4412_/B vssd1 vssd1 vccd1 vccd1 _4359_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7078_ _7091_/B _7091_/C _7091_/A vssd1 vssd1 vccd1 vccd1 _7094_/A sky130_fd_sc_hd__a21oi_4
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6029_ _6018_/A _4303_/C _6060_/A vssd1 vssd1 vccd1 vccd1 _6031_/A sky130_fd_sc_hd__a21o_2
XFILLER_100_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout30 _7430_/X vssd1 vssd1 vccd1 vccd1 _7889_/A sky130_fd_sc_hd__buf_6
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout74 _6871_/C vssd1 vssd1 vccd1 vccd1 _7247_/D sky130_fd_sc_hd__clkbuf_16
Xfanout41 _5244_/A vssd1 vssd1 vccd1 vccd1 _5530_/A sky130_fd_sc_hd__buf_12
Xfanout52 _5881_/A vssd1 vssd1 vccd1 vccd1 _5880_/A sky130_fd_sc_hd__buf_8
Xfanout63 _5070_/Y vssd1 vssd1 vccd1 vccd1 _7114_/B sky130_fd_sc_hd__clkbuf_16
Xfanout85 _5137_/X vssd1 vssd1 vccd1 vccd1 _6842_/B sky130_fd_sc_hd__buf_12
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout96 _4426_/X vssd1 vssd1 vccd1 vccd1 _5033_/A sky130_fd_sc_hd__buf_4
XFILLER_13_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6380_ _6368_/B _6379_/X _6431_/S vssd1 vssd1 vccd1 vccd1 _6381_/B sky130_fd_sc_hd__mux2_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5400_ _5621_/A _5672_/A vssd1 vssd1 vccd1 vccd1 _5401_/B sky130_fd_sc_hd__or2_4
X_5331_ _5530_/A _5797_/A vssd1 vssd1 vccd1 vccd1 _5332_/B sky130_fd_sc_hd__nor2_4
X_8050_ _8057_/CLK _8050_/D vssd1 vssd1 vccd1 vccd1 _8050_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_5_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5262_ _5262_/A _5262_/B vssd1 vssd1 vccd1 vccd1 _5482_/A sky130_fd_sc_hd__xnor2_4
X_7001_ _7001_/A _7150_/B vssd1 vssd1 vccd1 vccd1 _7007_/B sky130_fd_sc_hd__nor2_4
X_4213_ _8068_/Q _4213_/B vssd1 vssd1 vccd1 vccd1 _4221_/B sky130_fd_sc_hd__xor2_4
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5193_ _5541_/A _5342_/B vssd1 vssd1 vccd1 vccd1 _5259_/B sky130_fd_sc_hd__nor2_4
XFILLER_110_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4144_ _8076_/Q _8075_/Q _8077_/Q vssd1 vssd1 vccd1 vccd1 _4144_/X sky130_fd_sc_hd__or3_1
XFILLER_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4075_ _8061_/Q _4057_/B _4096_/A vssd1 vssd1 vccd1 vccd1 _4076_/B sky130_fd_sc_hd__o21ai_4
X_7903_ _7893_/X _7902_/X _7903_/B1 vssd1 vssd1 vccd1 vccd1 _7903_/Y sky130_fd_sc_hd__a21oi_2
X_7834_ _7908_/A _7834_/B vssd1 vssd1 vccd1 vccd1 _7834_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7765_ _7929_/A _7795_/A vssd1 vssd1 vccd1 vccd1 _7765_/X sky130_fd_sc_hd__or2_1
XFILLER_51_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6716_ _6749_/S _6716_/B vssd1 vssd1 vccd1 vccd1 _6716_/X sky130_fd_sc_hd__and2_1
X_4977_ _4979_/A _4979_/B _4979_/C vssd1 vssd1 vccd1 vccd1 _5050_/A sky130_fd_sc_hd__a21oi_1
X_7696_ _7928_/A _7696_/B vssd1 vssd1 vccd1 vccd1 _8032_/D sky130_fd_sc_hd__nor2_1
X_6647_ _6647_/A vssd1 vssd1 vccd1 vccd1 _6647_/Y sky130_fd_sc_hd__inv_2
X_6578_ _6578_/A _6578_/B vssd1 vssd1 vccd1 vccd1 _6594_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5529_ _5530_/A _5683_/B vssd1 vssd1 vccd1 vccd1 _5529_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout220 _7837_/A vssd1 vssd1 vccd1 vccd1 _7939_/A sky130_fd_sc_hd__clkbuf_4
Xfanout231 _4066_/A vssd1 vssd1 vccd1 vccd1 _4096_/A sky130_fd_sc_hd__buf_8
XFILLER_115_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4900_ _4900_/A _4900_/B vssd1 vssd1 vccd1 vccd1 _4902_/B sky130_fd_sc_hd__xnor2_4
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5880_ _5880_/A _5925_/A vssd1 vssd1 vccd1 vccd1 _5880_/Y sky130_fd_sc_hd__nor2_1
X_4831_ _5074_/A _5184_/A vssd1 vssd1 vccd1 vccd1 _4831_/X sky130_fd_sc_hd__or2_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7550_ _7549_/Y _7459_/A _7624_/S vssd1 vssd1 vccd1 vccd1 _7550_/X sky130_fd_sc_hd__mux2_1
X_4762_ _4763_/A _4763_/B vssd1 vssd1 vccd1 vccd1 _5095_/A sky130_fd_sc_hd__or2_2
X_6501_ _6444_/A _6444_/B _6447_/B vssd1 vssd1 vccd1 vccd1 _6501_/X sky130_fd_sc_hd__a21o_1
X_7481_ _7480_/X _7476_/X _7515_/S vssd1 vssd1 vccd1 vccd1 _7481_/X sky130_fd_sc_hd__mux2_1
X_4693_ _4606_/A _4606_/B _4606_/C vssd1 vssd1 vccd1 vccd1 _4693_/X sky130_fd_sc_hd__o21a_1
X_6432_ _6410_/B _6451_/B _6484_/S vssd1 vssd1 vccd1 vccd1 _6432_/X sky130_fd_sc_hd__mux2_1
X_6363_ _6488_/A _6484_/S _6363_/C vssd1 vssd1 vccd1 vccd1 _6443_/B sky130_fd_sc_hd__and3_1
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6294_ _6017_/B _6027_/A _6767_/S vssd1 vssd1 vccd1 vccd1 _6564_/A sky130_fd_sc_hd__mux2_4
X_5314_ _5314_/A _5314_/B vssd1 vssd1 vccd1 vccd1 _5503_/A sky130_fd_sc_hd__xor2_4
X_8033_ _8065_/CLK _8033_/D vssd1 vssd1 vccd1 vccd1 _8033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5245_ _5245_/A _5245_/B vssd1 vssd1 vccd1 vccd1 _5437_/B sky130_fd_sc_hd__xor2_4
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5176_ _5176_/A _5176_/B vssd1 vssd1 vccd1 vccd1 _5178_/B sky130_fd_sc_hd__xnor2_2
XFILLER_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4127_ _4074_/Y _4118_/X _4087_/B _4071_/Y vssd1 vssd1 vccd1 vccd1 _4127_/X sky130_fd_sc_hd__o211a_1
X_4058_ _8061_/Q _4058_/B vssd1 vssd1 vccd1 vccd1 _4059_/B sky130_fd_sc_hd__xnor2_4
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7817_ _7817_/A _7817_/B vssd1 vssd1 vccd1 vccd1 _7874_/C sky130_fd_sc_hd__xnor2_2
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7748_ _7748_/A _7748_/B _7749_/B vssd1 vssd1 vccd1 vccd1 _7769_/A sky130_fd_sc_hd__or3_1
X_7679_ _7720_/A _7679_/B vssd1 vssd1 vccd1 vccd1 _7682_/A sky130_fd_sc_hd__and2_1
XFILLER_118_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5030_ _5030_/A _5030_/B vssd1 vssd1 vccd1 vccd1 _5047_/A sky130_fd_sc_hd__xnor2_4
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6981_ _6983_/B _6995_/A _6983_/A vssd1 vssd1 vccd1 vccd1 _6991_/B sky130_fd_sc_hd__a21oi_4
XFILLER_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5932_ _6237_/S _5931_/Y _5914_/A vssd1 vssd1 vccd1 vccd1 _5932_/X sky130_fd_sc_hd__a21o_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5863_ _5879_/A _5879_/B vssd1 vssd1 vccd1 vccd1 _5863_/Y sky130_fd_sc_hd__nand2b_1
X_7602_ _8028_/Q _7879_/B _7562_/B vssd1 vssd1 vccd1 vccd1 _7602_/X sky130_fd_sc_hd__a21bo_1
XFILLER_61_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4814_ _4814_/A _4814_/B vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__or2_4
X_5794_ _5794_/A _5794_/B _5794_/C vssd1 vssd1 vccd1 vccd1 _5826_/A sky130_fd_sc_hd__nand3_4
X_7533_ _7481_/X _7515_/X _7538_/S vssd1 vssd1 vccd1 vccd1 _7542_/C sky130_fd_sc_hd__mux2_1
X_4745_ _4991_/A _5090_/B _4868_/B _4868_/C vssd1 vssd1 vccd1 vccd1 _4775_/A sky130_fd_sc_hd__nand4_4
X_7464_ _7449_/X _7453_/X _7483_/S vssd1 vssd1 vccd1 vccd1 _7464_/X sky130_fd_sc_hd__mux2_1
X_4676_ _4676_/A _4676_/B vssd1 vssd1 vccd1 vccd1 _4714_/A sky130_fd_sc_hd__nor2_1
X_7395_ _6368_/A _7513_/S _6350_/B vssd1 vssd1 vccd1 vccd1 _7401_/B sky130_fd_sc_hd__a21o_1
X_6415_ _6418_/A _6418_/B vssd1 vssd1 vccd1 vccd1 _6415_/X sky130_fd_sc_hd__and2b_1
Xposit_unit_242 vssd1 vssd1 vccd1 vccd1 posit_unit_242/HI io_out[0] sky130_fd_sc_hd__conb_1
X_6346_ _6488_/A _6359_/A vssd1 vssd1 vccd1 vccd1 _6441_/S sky130_fd_sc_hd__and2_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8016_ _8080_/CLK _8016_/D vssd1 vssd1 vccd1 vccd1 _8016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6277_ _6278_/A _6278_/B _4216_/C _4084_/B vssd1 vssd1 vccd1 vccd1 _6277_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5228_ _5957_/A _5229_/C vssd1 vssd1 vccd1 vccd1 _5230_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5159_ _5155_/A _5155_/B _5160_/B vssd1 vssd1 vccd1 vccd1 _5169_/A sky130_fd_sc_hd__a21bo_1
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4530_ _4530_/A _4530_/B vssd1 vssd1 vccd1 vccd1 _4537_/A sky130_fd_sc_hd__xnor2_4
X_4461_ _4461_/A _4461_/B vssd1 vssd1 vccd1 vccd1 _4467_/A sky130_fd_sc_hd__xor2_4
X_6200_ _6254_/S _6200_/B _6200_/C vssd1 vssd1 vccd1 vccd1 _6200_/X sky130_fd_sc_hd__and3_1
X_7180_ _7181_/A _7181_/B vssd1 vssd1 vccd1 vccd1 _7180_/X sky130_fd_sc_hd__and2b_1
XFILLER_98_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6131_ _6199_/S _6121_/Y _6129_/X vssd1 vssd1 vccd1 vccd1 _6131_/X sky130_fd_sc_hd__o21a_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4392_ _4392_/A _4392_/B vssd1 vssd1 vccd1 vccd1 _4393_/B sky130_fd_sc_hd__nand2_4
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6062_ _7558_/A _6304_/A vssd1 vssd1 vccd1 vccd1 _6065_/A sky130_fd_sc_hd__nor2_1
XFILLER_97_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5013_ _5013_/A _5013_/B _5013_/C _5040_/B vssd1 vssd1 vccd1 vccd1 _5016_/A sky130_fd_sc_hd__or4b_2
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6964_ _6964_/A _6964_/B vssd1 vssd1 vccd1 vccd1 _6966_/B sky130_fd_sc_hd__xnor2_2
X_6895_ _6895_/A _6895_/B vssd1 vssd1 vccd1 vccd1 _6987_/A sky130_fd_sc_hd__and2_1
X_5915_ _5915_/A _5915_/B vssd1 vssd1 vccd1 vccd1 _5916_/B sky130_fd_sc_hd__or2_1
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5846_ _5847_/A _6228_/A _5816_/A vssd1 vssd1 vccd1 vccd1 _5846_/Y sky130_fd_sc_hd__a21oi_1
X_5777_ _5777_/A _5777_/B vssd1 vssd1 vccd1 vccd1 _5808_/B sky130_fd_sc_hd__xor2_4
X_7516_ _7516_/A _7516_/B _7516_/C vssd1 vssd1 vccd1 vccd1 _7517_/B sky130_fd_sc_hd__and3_1
X_4728_ _4720_/X _4728_/B _4728_/C vssd1 vssd1 vccd1 vccd1 _4728_/X sky130_fd_sc_hd__and3b_1
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7447_ _7387_/B _7447_/B vssd1 vssd1 vccd1 vccd1 _7448_/B sky130_fd_sc_hd__and2b_1
X_4659_ _4625_/A _4625_/C _4625_/B vssd1 vssd1 vccd1 vccd1 _4660_/B sky130_fd_sc_hd__a21oi_2
XFILLER_89_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7378_ _7488_/A _7488_/B _7296_/X vssd1 vssd1 vccd1 vccd1 _7471_/B sky130_fd_sc_hd__a21oi_4
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6329_ _6330_/B vssd1 vssd1 vccd1 vccd1 _6329_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5700_ _5700_/A _5700_/B vssd1 vssd1 vccd1 vccd1 _5743_/B sky130_fd_sc_hd__xnor2_4
X_6680_ _6641_/B _6650_/B _6679_/X vssd1 vssd1 vccd1 vccd1 _6681_/B sky130_fd_sc_hd__a21oi_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5631_ _5723_/A _5919_/A _5631_/C vssd1 vssd1 vccd1 vccd1 _5631_/X sky130_fd_sc_hd__and3_1
X_5562_ _5562_/A _5562_/B vssd1 vssd1 vccd1 vccd1 _5579_/A sky130_fd_sc_hd__xnor2_2
X_7301_ _7301_/A _7301_/B vssd1 vssd1 vccd1 vccd1 _7327_/A sky130_fd_sc_hd__xnor2_4
X_4513_ _4513_/A _4513_/B vssd1 vssd1 vccd1 vccd1 _4519_/A sky130_fd_sc_hd__xnor2_4
X_5493_ _5487_/A _5486_/B _5484_/Y vssd1 vssd1 vccd1 vccd1 _5495_/B sky130_fd_sc_hd__a21oi_4
X_7232_ _7232_/A _7232_/B vssd1 vssd1 vccd1 vccd1 _7240_/B sky130_fd_sc_hd__xnor2_4
X_4444_ _4369_/Y _4424_/A _4424_/B _4413_/X _4377_/X vssd1 vssd1 vccd1 vccd1 _4444_/X
+ sky130_fd_sc_hd__a32o_1
X_7163_ _7281_/A _7281_/B _7195_/B _7269_/B vssd1 vssd1 vccd1 vccd1 _7169_/A sky130_fd_sc_hd__and4_4
X_4375_ _4501_/A _4455_/A vssd1 vssd1 vccd1 vccd1 _4424_/A sky130_fd_sc_hd__nor2_4
XFILLER_98_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7094_ _7094_/A _7094_/B vssd1 vssd1 vccd1 vccd1 _7097_/B sky130_fd_sc_hd__nor2_4
X_6114_ _6135_/A _6135_/B _5942_/A vssd1 vssd1 vccd1 vccd1 _6115_/B sky130_fd_sc_hd__o21bai_4
XFILLER_112_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6045_ _6088_/B _6091_/A vssd1 vssd1 vccd1 vccd1 _6045_/X sky130_fd_sc_hd__and2_4
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7996_ _8071_/Q _8015_/Q _8004_/S vssd1 vssd1 vccd1 vccd1 _8071_/D sky130_fd_sc_hd__mux2_1
X_6947_ _7334_/A _7235_/B _6947_/C _6943_/X vssd1 vssd1 vccd1 vccd1 _6978_/B sky130_fd_sc_hd__or4b_2
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6878_ _6877_/Y _6878_/B _6878_/C vssd1 vssd1 vccd1 vccd1 _6912_/A sky130_fd_sc_hd__and3b_1
XFILLER_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5829_ _7319_/B _5855_/A _5855_/B _5855_/C vssd1 vssd1 vccd1 vccd1 _5829_/Y sky130_fd_sc_hd__nor4_1
XFILLER_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4160_ _8079_/Q _4175_/B _4147_/B _4147_/C _4168_/B1 vssd1 vssd1 vccd1 vccd1 _4161_/B
+ sky130_fd_sc_hd__o41a_4
XFILLER_95_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4091_ _6326_/A _6274_/A vssd1 vssd1 vccd1 vccd1 _4095_/A sky130_fd_sc_hd__xor2_4
XFILLER_67_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7850_ _7846_/X _7874_/D _7918_/B vssd1 vssd1 vccd1 vccd1 _7850_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6801_ _7030_/A _6805_/B _6800_/C vssd1 vssd1 vccd1 vccd1 _6802_/B sky130_fd_sc_hd__o21ai_1
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7781_ _8034_/Q _4018_/X _7944_/B _8035_/Q vssd1 vssd1 vccd1 vccd1 _7781_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_51_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4993_ _4993_/A _4993_/B vssd1 vssd1 vccd1 vccd1 _5011_/B sky130_fd_sc_hd__xor2_4
X_6732_ _6732_/A _6732_/B _6732_/C _6732_/D vssd1 vssd1 vccd1 vccd1 _6732_/X sky130_fd_sc_hd__or4_1
XFILLER_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6663_ _6695_/S _6663_/B vssd1 vssd1 vccd1 vccd1 _6691_/B sky130_fd_sc_hd__or2_2
XFILLER_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5614_ _5614_/A _5614_/B vssd1 vssd1 vccd1 vccd1 _6123_/A sky130_fd_sc_hd__xnor2_2
X_6594_ _6594_/A _6594_/B vssd1 vssd1 vccd1 vccd1 _6595_/B sky130_fd_sc_hd__and2_1
X_5545_ _5545_/A _5545_/B vssd1 vssd1 vccd1 vccd1 _5547_/B sky130_fd_sc_hd__xor2_4
XFILLER_117_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5476_ _5491_/A vssd1 vssd1 vccd1 vccd1 _5476_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4427_ _5013_/A vssd1 vssd1 vccd1 vccd1 _4947_/A sky130_fd_sc_hd__inv_2
X_7215_ _7215_/A _7371_/B vssd1 vssd1 vccd1 vccd1 _7251_/A sky130_fd_sc_hd__nor2_4
XFILLER_59_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7146_ _7146_/A _7146_/B vssd1 vssd1 vccd1 vccd1 _7157_/B sky130_fd_sc_hd__xnor2_4
XFILLER_113_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4358_ _4356_/A _4406_/A _4551_/A vssd1 vssd1 vccd1 vccd1 _4412_/B sky130_fd_sc_hd__a21o_4
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4289_ _4287_/X _4288_/X _4341_/A1 vssd1 vssd1 vccd1 vccd1 _4354_/B sky130_fd_sc_hd__o21ai_4
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7077_ _7111_/A _7111_/B vssd1 vssd1 vccd1 vccd1 _7091_/C sky130_fd_sc_hd__or2_2
XFILLER_104_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6028_ _6017_/B _6027_/Y _6026_/X vssd1 vssd1 vccd1 vccd1 _6088_/B sky130_fd_sc_hd__o21a_4
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7979_ _8015_/Q _8055_/Q _7986_/S vssd1 vssd1 vccd1 vccd1 _8055_/D sky130_fd_sc_hd__mux2_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout20 _6733_/S vssd1 vssd1 vccd1 vccd1 _6751_/S sky130_fd_sc_hd__buf_4
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout31 _7430_/X vssd1 vssd1 vccd1 vccd1 _7847_/A sky130_fd_sc_hd__buf_4
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout42 _6739_/S vssd1 vssd1 vccd1 vccd1 _6713_/S sky130_fd_sc_hd__buf_4
Xfanout64 _5070_/Y vssd1 vssd1 vccd1 vccd1 _5782_/A sky130_fd_sc_hd__buf_4
Xfanout53 _5034_/B vssd1 vssd1 vccd1 vccd1 _5040_/B sky130_fd_sc_hd__buf_6
Xfanout97 _6448_/S vssd1 vssd1 vccd1 vccd1 _6766_/S sky130_fd_sc_hd__buf_8
Xfanout86 _5137_/X vssd1 vssd1 vccd1 vccd1 _6778_/B sky130_fd_sc_hd__buf_6
XFILLER_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout75 _7319_/B vssd1 vssd1 vccd1 vccd1 _7306_/B sky130_fd_sc_hd__buf_8
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5330_ _5330_/A _5330_/B vssd1 vssd1 vccd1 vccd1 _5332_/A sky130_fd_sc_hd__xnor2_4
X_5261_ _5262_/A _5262_/B vssd1 vssd1 vccd1 vccd1 _5261_/X sky130_fd_sc_hd__and2b_1
X_4212_ _8068_/Q _4213_/B vssd1 vssd1 vccd1 vccd1 _4212_/Y sky130_fd_sc_hd__xnor2_4
X_7000_ _7334_/A _7150_/B _7046_/B _7366_/A vssd1 vssd1 vccd1 vccd1 _7000_/X sky130_fd_sc_hd__o22a_1
X_5192_ _7046_/B _5516_/A vssd1 vssd1 vccd1 vccd1 _5259_/A sky130_fd_sc_hd__or2_4
X_4143_ _4175_/B _4147_/B vssd1 vssd1 vccd1 vccd1 _4241_/A sky130_fd_sc_hd__nor2_1
XFILLER_110_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4074_ _6272_/A _6289_/A vssd1 vssd1 vccd1 vccd1 _4074_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7902_ _7900_/X _7901_/Y _6269_/X _7888_/Y vssd1 vssd1 vccd1 vccd1 _7902_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_83_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7833_ _7833_/A _7833_/B _7833_/C _7833_/D vssd1 vssd1 vccd1 vccd1 _7883_/A sky130_fd_sc_hd__and4_4
XFILLER_91_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7764_ _7764_/A _7764_/B vssd1 vssd1 vccd1 vccd1 _7795_/A sky130_fd_sc_hd__nor2_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6715_ _6708_/X _6714_/X _6753_/S vssd1 vssd1 vccd1 vccd1 _6716_/B sky130_fd_sc_hd__mux2_1
XFILLER_11_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4976_ _4976_/A _4976_/B vssd1 vssd1 vccd1 vccd1 _4979_/C sky130_fd_sc_hd__xnor2_4
X_7695_ _8032_/Q _7857_/B _7693_/Y _7694_/Y vssd1 vssd1 vccd1 vccd1 _7696_/B sky130_fd_sc_hd__o2bb2a_1
X_6646_ _6546_/A _6581_/B _6688_/S vssd1 vssd1 vccd1 vccd1 _6647_/A sky130_fd_sc_hd__mux2_1
X_6577_ _6577_/A _6641_/B vssd1 vssd1 vccd1 vccd1 _6578_/B sky130_fd_sc_hd__nand2_1
X_5528_ _5582_/A _5855_/A vssd1 vssd1 vccd1 vccd1 _5531_/B sky130_fd_sc_hd__or2_4
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5459_ _5459_/A _5459_/B vssd1 vssd1 vccd1 vccd1 _5462_/A sky130_fd_sc_hd__xnor2_4
Xfanout232 _6188_/A vssd1 vssd1 vccd1 vccd1 _4066_/A sky130_fd_sc_hd__buf_4
Xfanout221 _6187_/X vssd1 vssd1 vccd1 vccd1 _7837_/A sky130_fd_sc_hd__buf_4
Xfanout210 _7949_/B vssd1 vssd1 vccd1 vccd1 _5207_/A sky130_fd_sc_hd__buf_6
XFILLER_101_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7129_ _7130_/B _7130_/A vssd1 vssd1 vccd1 vccd1 _7129_/X sky130_fd_sc_hd__and2b_1
XFILLER_115_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4830_ _5074_/B _4830_/B vssd1 vssd1 vccd1 vccd1 _5184_/A sky130_fd_sc_hd__nand2_4
XFILLER_60_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ _4761_/A _4761_/B vssd1 vssd1 vccd1 vccd1 _4763_/B sky130_fd_sc_hd__xor2_1
X_6500_ _6550_/B _6550_/D _6550_/C vssd1 vssd1 vccd1 vccd1 _6500_/Y sky130_fd_sc_hd__o21bai_4
X_7480_ _7478_/X _7479_/X _7527_/S vssd1 vssd1 vccd1 vccd1 _7480_/X sky130_fd_sc_hd__mux2_1
X_4692_ _4691_/A _4712_/A _4690_/A vssd1 vssd1 vccd1 vccd1 _4692_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6431_ _6420_/X _6430_/X _6431_/S vssd1 vssd1 vccd1 vccd1 _6451_/B sky130_fd_sc_hd__mux2_1
X_6362_ _6484_/S _6363_/C vssd1 vssd1 vccd1 vccd1 _6362_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5313_ _5314_/A _5314_/B vssd1 vssd1 vccd1 vccd1 _5313_/Y sky130_fd_sc_hd__nor2_1
X_6293_ _6034_/Y _6031_/B _6766_/S vssd1 vssd1 vccd1 vccd1 _6299_/A sky130_fd_sc_hd__mux2_4
XFILLER_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8032_ _8065_/CLK _8032_/D vssd1 vssd1 vccd1 vccd1 _8032_/Q sky130_fd_sc_hd__dfxtp_1
X_5244_ _5244_/A _5715_/A vssd1 vssd1 vccd1 vccd1 _5437_/A sky130_fd_sc_hd__nor2_4
X_5175_ _5232_/B _5175_/B _5176_/B vssd1 vssd1 vccd1 vccd1 _5230_/A sky130_fd_sc_hd__or3b_2
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4126_ _4078_/A _4119_/Y _4087_/B _4111_/A vssd1 vssd1 vccd1 vccd1 _4126_/X sky130_fd_sc_hd__a211o_1
XFILLER_56_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4057_ _4066_/A _4057_/B vssd1 vssd1 vccd1 vccd1 _4058_/B sky130_fd_sc_hd__nand2_2
XFILLER_83_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7816_ _7817_/A _7817_/B vssd1 vssd1 vccd1 vccd1 _7848_/A sky130_fd_sc_hd__and2b_1
XFILLER_64_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7747_ _7470_/Y _7746_/Y _7847_/A vssd1 vssd1 vccd1 vccd1 _7749_/B sky130_fd_sc_hd__mux2_2
XFILLER_51_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4959_ _4959_/A _4959_/B vssd1 vssd1 vccd1 vccd1 _4995_/A sky130_fd_sc_hd__xor2_4
X_7678_ _7677_/A _7677_/B _7677_/C vssd1 vssd1 vccd1 vccd1 _7679_/B sky130_fd_sc_hd__a21o_1
X_6629_ _6629_/A _6629_/B vssd1 vssd1 vccd1 vccd1 _6629_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_118_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6980_ _6994_/A _6994_/B vssd1 vssd1 vccd1 vccd1 _6995_/A sky130_fd_sc_hd__nand2_4
XFILLER_65_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5931_ _6236_/A _5931_/B vssd1 vssd1 vccd1 vccd1 _5931_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5862_ _5862_/A _5886_/A vssd1 vssd1 vccd1 vccd1 _5879_/B sky130_fd_sc_hd__xnor2_2
XFILLER_33_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7601_ _7923_/A _7588_/X _7589_/Y _7903_/B1 vssd1 vssd1 vccd1 vccd1 _7601_/X sky130_fd_sc_hd__a31o_1
X_4813_ _4813_/A _4813_/B _4816_/A vssd1 vssd1 vccd1 vccd1 _4814_/B sky130_fd_sc_hd__nor3_1
X_5793_ _5824_/A _5824_/B vssd1 vssd1 vccd1 vccd1 _5794_/C sky130_fd_sc_hd__and2_2
X_7532_ _7525_/Y _7527_/X _7530_/X _7531_/X vssd1 vssd1 vccd1 vccd1 _7537_/D sky130_fd_sc_hd__a22o_1
X_4744_ _4989_/A _4988_/A _4751_/C _4773_/A vssd1 vssd1 vccd1 vccd1 _4868_/C sky130_fd_sc_hd__a211oi_4
X_7463_ _7443_/X _7446_/X _7502_/B vssd1 vssd1 vccd1 vccd1 _7463_/X sky130_fd_sc_hd__mux2_1
X_4675_ _4675_/A _4675_/B vssd1 vssd1 vccd1 vccd1 _4676_/B sky130_fd_sc_hd__and2_1
X_6414_ _4343_/Y _7281_/C _6445_/S vssd1 vssd1 vccd1 vccd1 _6418_/B sky130_fd_sc_hd__mux2_1
X_7394_ _7454_/A _7454_/B _7455_/S vssd1 vssd1 vccd1 vccd1 _7394_/X sky130_fd_sc_hd__a21o_1
Xposit_unit_243 vssd1 vssd1 vccd1 vccd1 posit_unit_243/HI io_out[1] sky130_fd_sc_hd__conb_1
X_6345_ _6064_/Y _6340_/X _6341_/Y _6344_/X vssd1 vssd1 vccd1 vccd1 _6359_/A sky130_fd_sc_hd__a211oi_4
X_6276_ _4084_/B _4216_/C _4221_/B _4087_/B _6275_/X vssd1 vssd1 vccd1 vccd1 _6276_/X
+ sky130_fd_sc_hd__o221a_1
X_8015_ _8079_/CLK _8015_/D vssd1 vssd1 vccd1 vccd1 _8015_/Q sky130_fd_sc_hd__dfxtp_1
X_5227_ _5227_/A _5227_/B vssd1 vssd1 vccd1 vccd1 _5229_/C sky130_fd_sc_hd__and2_1
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5158_ _5227_/A _5158_/B vssd1 vssd1 vccd1 vccd1 _5160_/B sky130_fd_sc_hd__and2_1
XFILLER_56_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4109_ _4064_/B _4108_/Y _4079_/B vssd1 vssd1 vccd1 vccd1 _6018_/A sky130_fd_sc_hd__a21oi_4
X_5089_ _7213_/A _5082_/X _5085_/X _5087_/X vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__a31o_2
XFILLER_71_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4460_ _4460_/A _4460_/B vssd1 vssd1 vccd1 vccd1 _4461_/B sky130_fd_sc_hd__xor2_4
X_4391_ _4456_/B _7306_/A _4585_/B _4551_/A vssd1 vssd1 vccd1 vccd1 _4392_/B sky130_fd_sc_hd__a22o_1
X_6130_ _6199_/S _6121_/Y _6129_/X vssd1 vssd1 vccd1 vccd1 _6130_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_98_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6061_ _6326_/A _6326_/B vssd1 vssd1 vccd1 vccd1 _6304_/A sky130_fd_sc_hd__nand2_4
XFILLER_85_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _4984_/A _4984_/C _4984_/B vssd1 vssd1 vccd1 vccd1 _5018_/B sky130_fd_sc_hd__a21o_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6963_ _6978_/B _6978_/C _6978_/A vssd1 vssd1 vccd1 vccd1 _6983_/B sky130_fd_sc_hd__a21o_2
X_6894_ _6894_/A _6894_/B vssd1 vssd1 vccd1 vccd1 _6895_/B sky130_fd_sc_hd__nand2_1
X_5914_ _5914_/A _5914_/B vssd1 vssd1 vccd1 vccd1 _6237_/S sky130_fd_sc_hd__nor2_1
XFILLER_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5845_ _5848_/A _5848_/B vssd1 vssd1 vccd1 vccd1 _6228_/A sky130_fd_sc_hd__or2_1
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5776_ _5776_/A _5776_/B vssd1 vssd1 vccd1 vccd1 _5777_/B sky130_fd_sc_hd__xnor2_4
X_7515_ _7491_/X _7514_/X _7515_/S vssd1 vssd1 vccd1 vccd1 _7515_/X sky130_fd_sc_hd__mux2_1
X_4727_ _4727_/A _4727_/B _4837_/A _4837_/B vssd1 vssd1 vccd1 vccd1 _4728_/C sky130_fd_sc_hd__nor4_1
X_7446_ _7442_/X _7445_/Y _7479_/S vssd1 vssd1 vccd1 vccd1 _7446_/X sky130_fd_sc_hd__mux2_1
X_4658_ _4675_/A _4675_/B vssd1 vssd1 vccd1 vccd1 _4676_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7377_ _7325_/B _7487_/B _7323_/Y vssd1 vssd1 vccd1 vccd1 _7488_/B sky130_fd_sc_hd__a21o_4
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4589_ _4627_/A _4589_/B vssd1 vssd1 vccd1 vccd1 _4596_/A sky130_fd_sc_hd__xor2_4
XFILLER_103_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6328_ _6020_/A _6296_/X _6767_/S vssd1 vssd1 vccd1 vccd1 _6330_/B sky130_fd_sc_hd__mux2_2
XFILLER_103_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6259_ _6259_/A _6259_/B _6259_/C vssd1 vssd1 vccd1 vccd1 _6259_/X sky130_fd_sc_hd__and3_1
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5630_ _5723_/A _5919_/A vssd1 vssd1 vccd1 vccd1 _5676_/A sky130_fd_sc_hd__nand2_4
XFILLER_31_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5561_ _5561_/A _5561_/B vssd1 vssd1 vccd1 vccd1 _5600_/A sky130_fd_sc_hd__xnor2_4
X_5492_ _5492_/A _5492_/B vssd1 vssd1 vccd1 vccd1 _5495_/A sky130_fd_sc_hd__xnor2_4
X_7300_ _7300_/A _7300_/B vssd1 vssd1 vccd1 vccd1 _7320_/A sky130_fd_sc_hd__xor2_4
XFILLER_8_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4512_ _4513_/A _4513_/B vssd1 vssd1 vccd1 vccd1 _4512_/Y sky130_fd_sc_hd__nand2_1
XFILLER_105_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7231_ _7232_/A _7232_/B vssd1 vssd1 vccd1 vccd1 _7231_/Y sky130_fd_sc_hd__nand2b_1
X_4443_ _4424_/A _4413_/B _4442_/X vssd1 vssd1 vccd1 vccd1 _4443_/Y sky130_fd_sc_hd__a21oi_1
X_4374_ _7215_/A _4371_/X _4372_/X _4373_/Y _4361_/X vssd1 vssd1 vccd1 vccd1 _4374_/X
+ sky130_fd_sc_hd__a32o_1
X_7162_ _7281_/A _7269_/B vssd1 vssd1 vccd1 vccd1 _7162_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6113_ _6259_/A _6192_/B _6192_/C vssd1 vssd1 vccd1 vccd1 _6113_/X sky130_fd_sc_hd__or3_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7093_ _7110_/A _7110_/B vssd1 vssd1 vccd1 vccd1 _7094_/B sky130_fd_sc_hd__and2b_2
XFILLER_100_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6044_ _6044_/A _6044_/B vssd1 vssd1 vccd1 vccd1 _6091_/A sky130_fd_sc_hd__nor2_4
XFILLER_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7995_ _8070_/Q _8014_/Q _8004_/S vssd1 vssd1 vccd1 vccd1 _8070_/D sky130_fd_sc_hd__mux2_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6946_ _7334_/A _7235_/B _6947_/C vssd1 vssd1 vccd1 vccd1 _6998_/A sky130_fd_sc_hd__or3_1
XFILLER_22_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6877_ _6877_/A _6877_/B vssd1 vssd1 vccd1 vccd1 _6877_/Y sky130_fd_sc_hd__xnor2_1
X_5828_ _5855_/A _5853_/B vssd1 vssd1 vccd1 vccd1 _5889_/B sky130_fd_sc_hd__nor2_4
XFILLER_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5759_ _5759_/A _5759_/B _5759_/C vssd1 vssd1 vccd1 vccd1 _5762_/A sky130_fd_sc_hd__nand3_4
XFILLER_108_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7429_ _7430_/A _7430_/B vssd1 vssd1 vccd1 vccd1 _7766_/B sky130_fd_sc_hd__nor2_8
XFILLER_118_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4090_ _8057_/Q _4090_/B vssd1 vssd1 vccd1 vccd1 _6274_/A sky130_fd_sc_hd__xor2_4
XFILLER_95_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6800_ _7030_/A _6800_/B _6800_/C vssd1 vssd1 vccd1 vccd1 _6804_/B sky130_fd_sc_hd__or3_2
XFILLER_36_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7780_ _7763_/X _7772_/Y _7779_/X _7903_/B1 vssd1 vssd1 vccd1 vccd1 _7780_/X sky130_fd_sc_hd__a31o_2
XFILLER_91_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4992_ _4992_/A _4992_/B vssd1 vssd1 vccd1 vccd1 _5011_/A sky130_fd_sc_hd__xnor2_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6731_ _6727_/X _6730_/A _6749_/S vssd1 vssd1 vccd1 vccd1 _6732_/D sky130_fd_sc_hd__mux2_1
X_6662_ _6661_/Y _6655_/B _6691_/A vssd1 vssd1 vccd1 vccd1 _6662_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_2__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _8077_/CLK sky130_fd_sc_hd__clkbuf_16
X_5613_ _5613_/A _5613_/B vssd1 vssd1 vccd1 vccd1 _5614_/B sky130_fd_sc_hd__nand2_2
X_6593_ _6592_/A _6592_/B _6615_/A _6613_/B vssd1 vssd1 vccd1 vccd1 _6611_/A sky130_fd_sc_hd__o22a_1
XFILLER_117_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5544_ _5538_/A _5536_/Y _5535_/Y vssd1 vssd1 vccd1 vccd1 _5547_/A sky130_fd_sc_hd__o21ai_4
X_5475_ _5477_/A _5477_/B _5477_/C vssd1 vssd1 vccd1 vccd1 _5491_/A sky130_fd_sc_hd__a21o_4
X_4426_ _4411_/B _4425_/X _4494_/A vssd1 vssd1 vccd1 vccd1 _4426_/X sky130_fd_sc_hd__mux2_4
X_7214_ _7214_/A _7247_/D _7216_/A vssd1 vssd1 vccd1 vccd1 _7214_/X sky130_fd_sc_hd__or3_1
X_7145_ _7182_/A _7182_/B _7143_/B _7142_/B _7142_/A vssd1 vssd1 vccd1 vccd1 _7157_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4357_ _4547_/C _4406_/A _7213_/B vssd1 vssd1 vccd1 vccd1 _4407_/A sky130_fd_sc_hd__a21oi_4
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4288_ _4199_/X _5989_/B _4250_/X _4315_/B vssd1 vssd1 vccd1 vccd1 _4288_/X sky130_fd_sc_hd__o211a_2
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7076_ _7076_/A _7076_/B vssd1 vssd1 vccd1 vccd1 _7111_/B sky130_fd_sc_hd__xnor2_4
X_6027_ _6027_/A _7413_/A vssd1 vssd1 vccd1 vccd1 _6027_/Y sky130_fd_sc_hd__nand2_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7978_ _8014_/Q _8054_/Q _7986_/S vssd1 vssd1 vccd1 vccd1 _8054_/D sky130_fd_sc_hd__mux2_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout21 _6610_/Y vssd1 vssd1 vccd1 vccd1 _6733_/S sky130_fd_sc_hd__buf_6
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout10 _6113_/X vssd1 vssd1 vccd1 vccd1 _6262_/S sky130_fd_sc_hd__buf_4
X_6929_ _6931_/B _6931_/C _6931_/A vssd1 vssd1 vccd1 vccd1 _6987_/B sky130_fd_sc_hd__o21a_1
Xfanout32 _6590_/B vssd1 vssd1 vccd1 vccd1 _6737_/B sky130_fd_sc_hd__buf_4
Xfanout43 _6614_/A vssd1 vssd1 vccd1 vccd1 _6739_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_80_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout65 _7150_/B vssd1 vssd1 vccd1 vccd1 _5367_/A sky130_fd_sc_hd__clkbuf_16
Xfanout54 _4878_/A vssd1 vssd1 vccd1 vccd1 _5013_/C sky130_fd_sc_hd__buf_4
Xfanout98 _6448_/S vssd1 vssd1 vccd1 vccd1 _6767_/S sky130_fd_sc_hd__buf_6
Xfanout76 _5271_/Y vssd1 vssd1 vccd1 vccd1 _7319_/B sky130_fd_sc_hd__clkbuf_16
Xfanout87 _7195_/B vssd1 vssd1 vccd1 vccd1 _6878_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_22_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5260_ _5459_/A _5459_/B vssd1 vssd1 vccd1 vccd1 _5262_/B sky130_fd_sc_hd__and2_2
X_4211_ _8067_/Q _4211_/B vssd1 vssd1 vccd1 vccd1 _4213_/B sky130_fd_sc_hd__nand2_8
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5191_ _5541_/A _5516_/A vssd1 vssd1 vccd1 vccd1 _5191_/X sky130_fd_sc_hd__or2_1
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4142_ _8074_/Q _8072_/Q _8071_/Q _8073_/Q vssd1 vssd1 vccd1 vccd1 _4147_/B sky130_fd_sc_hd__or4_4
XFILLER_68_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4073_ _6060_/A _6289_/A vssd1 vssd1 vccd1 vccd1 _4078_/A sky130_fd_sc_hd__xnor2_4
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7901_ _7900_/A _7900_/B _6774_/X vssd1 vssd1 vccd1 vccd1 _7901_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_64_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7832_ _7834_/B vssd1 vssd1 vccd1 vccd1 _7833_/D sky130_fd_sc_hd__inv_2
X_7763_ _7763_/A _7763_/B vssd1 vssd1 vccd1 vccd1 _7763_/X sky130_fd_sc_hd__or2_1
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4975_ _4980_/B _4980_/A vssd1 vssd1 vccd1 vccd1 _4979_/B sky130_fd_sc_hd__nand2b_1
X_6714_ _6698_/X _6713_/X _6751_/S vssd1 vssd1 vccd1 vccd1 _6714_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7694_ _8031_/Q _7964_/C _7562_/B vssd1 vssd1 vccd1 vccd1 _7694_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_20_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6645_ _6645_/A _6645_/B vssd1 vssd1 vccd1 vccd1 _6645_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6576_ _6580_/A _6580_/B vssd1 vssd1 vccd1 vccd1 _6594_/A sky130_fd_sc_hd__nand2b_1
X_5527_ _5683_/A _5855_/A vssd1 vssd1 vccd1 vccd1 _5639_/A sky130_fd_sc_hd__or2_4
XFILLER_105_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5458_ _5451_/A _5451_/B _5442_/Y vssd1 vssd1 vccd1 vccd1 _5473_/A sky130_fd_sc_hd__a21o_2
XFILLER_115_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout222 _6522_/S vssd1 vssd1 vccd1 vccd1 _7728_/A sky130_fd_sc_hd__buf_6
Xfanout200 _5106_/Y vssd1 vssd1 vccd1 vccd1 _6800_/B sky130_fd_sc_hd__buf_12
Xfanout211 _4352_/Y vssd1 vssd1 vccd1 vccd1 _7949_/B sky130_fd_sc_hd__clkbuf_16
X_4409_ _4436_/A _4402_/X _4406_/X _4408_/Y vssd1 vssd1 vccd1 vccd1 _4409_/X sky130_fd_sc_hd__o211a_1
X_5389_ _5389_/A _5389_/B vssd1 vssd1 vccd1 vccd1 _5391_/B sky130_fd_sc_hd__xnor2_4
Xfanout233 _8066_/Q vssd1 vssd1 vccd1 vccd1 _6188_/A sky130_fd_sc_hd__buf_8
X_7128_ _7128_/A _7128_/B vssd1 vssd1 vccd1 vccd1 _7130_/B sky130_fd_sc_hd__xnor2_2
XFILLER_115_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7059_ _7101_/A _7001_/A _7124_/A2 _7334_/A vssd1 vssd1 vccd1 vccd1 _7059_/X sky130_fd_sc_hd__o22a_1
XFILLER_47_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4760_ _4761_/B _4761_/A vssd1 vssd1 vccd1 vccd1 _5093_/A sky130_fd_sc_hd__nand2b_1
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4691_ _4691_/A _4712_/A vssd1 vssd1 vccd1 vccd1 _4691_/X sky130_fd_sc_hd__and2_1
X_6430_ _7281_/D _7306_/A _6456_/S vssd1 vssd1 vccd1 vccd1 _6430_/X sky130_fd_sc_hd__mux2_1
X_6361_ _6354_/A _6360_/X _6431_/S vssd1 vssd1 vccd1 vccd1 _6363_/C sky130_fd_sc_hd__mux2_2
XFILLER_115_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5312_ _5504_/A _5504_/B _5621_/A _5306_/S vssd1 vssd1 vccd1 vccd1 _5314_/B sky130_fd_sc_hd__o2bb2a_4
XFILLER_114_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6292_ _6271_/Y _6273_/X _6291_/X _6272_/Y vssd1 vssd1 vccd1 vccd1 _6448_/S sky130_fd_sc_hd__a31o_4
XFILLER_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8031_ _8065_/CLK _8031_/D vssd1 vssd1 vccd1 vccd1 _8031_/Q sky130_fd_sc_hd__dfxtp_1
X_5243_ _5243_/A _6778_/B vssd1 vssd1 vccd1 vccd1 _5245_/B sky130_fd_sc_hd__nor2_4
X_5174_ _5174_/A _5174_/B _6951_/D vssd1 vssd1 vccd1 vccd1 _5176_/B sky130_fd_sc_hd__and3_2
XFILLER_96_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4125_ _4084_/B _5134_/A2 _4122_/X _5135_/C1 vssd1 vssd1 vccd1 vccd1 _4125_/X sky130_fd_sc_hd__a211o_2
X_4056_ _4117_/A _4117_/B _4056_/S vssd1 vssd1 vccd1 vccd1 _4064_/A sky130_fd_sc_hd__mux2_4
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7815_ _7766_/B _7594_/A _7766_/Y vssd1 vssd1 vccd1 vccd1 _7817_/B sky130_fd_sc_hd__a21oi_2
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7746_ _7657_/B _7624_/X _7657_/Y vssd1 vssd1 vccd1 vccd1 _7746_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_61_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4958_ _5033_/B _4991_/A vssd1 vssd1 vccd1 vccd1 _4959_/B sky130_fd_sc_hd__nand2b_4
X_7677_ _7677_/A _7677_/B _7677_/C vssd1 vssd1 vccd1 vccd1 _7720_/A sky130_fd_sc_hd__nand3_4
X_4889_ _4847_/X _4848_/Y _4773_/A _4988_/A vssd1 vssd1 vccd1 vccd1 _4919_/C sky130_fd_sc_hd__a211o_4
X_6628_ _6628_/A _6628_/B vssd1 vssd1 vccd1 vccd1 _6629_/B sky130_fd_sc_hd__xnor2_1
X_6559_ _6559_/A _6565_/A vssd1 vssd1 vccd1 vccd1 _6560_/B sky130_fd_sc_hd__and2_1
XFILLER_106_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5930_ _6236_/B _5929_/X _5919_/X vssd1 vssd1 vccd1 vccd1 _5931_/B sky130_fd_sc_hd__o21ba_1
XFILLER_46_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7600_ _7918_/B _7600_/B _7600_/C vssd1 vssd1 vccd1 vccd1 _7600_/Y sky130_fd_sc_hd__nor3_1
X_5861_ _5885_/A _5885_/B vssd1 vssd1 vccd1 vccd1 _5886_/A sky130_fd_sc_hd__nor2_2
XFILLER_34_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4812_ _4814_/A vssd1 vssd1 vccd1 vccd1 _4812_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5792_ _5822_/A _5822_/B vssd1 vssd1 vccd1 vccd1 _5824_/B sky130_fd_sc_hd__nor2_4
XFILLER_33_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7531_ _7538_/S _7531_/B _7531_/C _7534_/B vssd1 vssd1 vccd1 vccd1 _7531_/X sky130_fd_sc_hd__or4_1
X_4743_ _4773_/A _4989_/A _4988_/A _4751_/C vssd1 vssd1 vccd1 vccd1 _4868_/B sky130_fd_sc_hd__or4_4
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7462_ _7537_/B vssd1 vssd1 vccd1 vccd1 _7462_/Y sky130_fd_sc_hd__inv_2
X_6413_ _6488_/B _6413_/B vssd1 vssd1 vccd1 vccd1 _6418_/A sky130_fd_sc_hd__or2_2
X_4674_ _4670_/B _4670_/C _4670_/A vssd1 vssd1 vccd1 vccd1 _4689_/B sky130_fd_sc_hd__a21o_1
Xposit_unit_244 vssd1 vssd1 vccd1 vccd1 posit_unit_244/HI io_out[2] sky130_fd_sc_hd__conb_1
X_7393_ _6831_/A _6831_/B _7392_/X vssd1 vssd1 vccd1 vccd1 _7455_/S sky130_fd_sc_hd__a21o_1
XFILLER_115_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6344_ _6325_/Y _6342_/X _6343_/Y vssd1 vssd1 vccd1 vccd1 _6344_/X sky130_fd_sc_hd__a21o_1
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6275_ _8052_/Q _4221_/B _4315_/A _4088_/A vssd1 vssd1 vccd1 vccd1 _6275_/X sky130_fd_sc_hd__a211o_1
X_8014_ _8079_/CLK _8014_/D vssd1 vssd1 vccd1 vccd1 _8014_/Q sky130_fd_sc_hd__dfxtp_2
X_5226_ _5957_/A vssd1 vssd1 vccd1 vccd1 _5226_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5157_ _6806_/A _5244_/A _5156_/C vssd1 vssd1 vccd1 vccd1 _5158_/B sky130_fd_sc_hd__o21ai_1
XFILLER_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4108_ _4103_/A _4107_/Y _4064_/A vssd1 vssd1 vccd1 vccd1 _4108_/Y sky130_fd_sc_hd__o21ai_2
X_5088_ _7213_/A _5082_/X _5085_/X _5087_/X vssd1 vssd1 vccd1 vccd1 _5088_/Y sky130_fd_sc_hd__a31oi_4
X_4039_ _4088_/A _8054_/Q _8053_/Q _8052_/Q vssd1 vssd1 vccd1 vccd1 _4096_/B sky130_fd_sc_hd__or4_4
XFILLER_72_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7729_ _6225_/S _7608_/Y _7639_/Y vssd1 vssd1 vccd1 vccd1 _7729_/X sky130_fd_sc_hd__a21bo_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4390_ _7214_/A _5090_/A _7247_/A _4585_/B vssd1 vssd1 vccd1 vccd1 _4392_/A sky130_fd_sc_hd__or4b_4
XFILLER_97_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _6060_/A _6272_/B vssd1 vssd1 vccd1 vccd1 _6060_/Y sky130_fd_sc_hd__nor2_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _5011_/A _5011_/B vssd1 vssd1 vccd1 vccd1 _5027_/A sky130_fd_sc_hd__xor2_4
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6962_ _6996_/A _6996_/B vssd1 vssd1 vccd1 vccd1 _6978_/C sky130_fd_sc_hd__nand2_1
XFILLER_81_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6893_ _6893_/A _6893_/B vssd1 vssd1 vccd1 vccd1 _6936_/A sky130_fd_sc_hd__xor2_1
X_5913_ _5912_/A _5912_/B _5912_/C vssd1 vssd1 vccd1 vccd1 _5914_/B sky130_fd_sc_hd__a21oi_1
X_5844_ _5850_/A _5850_/B _5841_/X vssd1 vssd1 vccd1 vccd1 _5848_/B sky130_fd_sc_hd__a21oi_2
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7514_ _7513_/X _7509_/X _7527_/S vssd1 vssd1 vccd1 vccd1 _7514_/X sky130_fd_sc_hd__mux2_1
X_5775_ _5804_/A _5804_/B _5766_/Y vssd1 vssd1 vccd1 vccd1 _5777_/A sky130_fd_sc_hd__o21a_4
X_4726_ _4726_/A _4726_/B vssd1 vssd1 vccd1 vccd1 _4726_/Y sky130_fd_sc_hd__nor2_1
X_7445_ _7445_/A _7445_/B vssd1 vssd1 vccd1 vccd1 _7445_/Y sky130_fd_sc_hd__xnor2_1
X_4657_ _4663_/A _4663_/B vssd1 vssd1 vccd1 vccd1 _4675_/B sky130_fd_sc_hd__xnor2_1
X_7376_ _7508_/A _7508_/B _7347_/X vssd1 vssd1 vccd1 vccd1 _7487_/B sky130_fd_sc_hd__a21o_1
XFILLER_107_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6327_ _6336_/A _6327_/B vssd1 vssd1 vccd1 vccd1 _6330_/A sky130_fd_sc_hd__nand2b_1
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4588_ _4627_/A _4589_/B vssd1 vssd1 vccd1 vccd1 _4588_/X sky130_fd_sc_hd__and2_1
XFILLER_115_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6258_ _7611_/D _6258_/B _6258_/C _6258_/D vssd1 vssd1 vccd1 vccd1 _6258_/X sky130_fd_sc_hd__or4_1
XFILLER_67_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6189_ _6081_/Y _6111_/B _6111_/C _6163_/D vssd1 vssd1 vccd1 vccd1 _6189_/X sky130_fd_sc_hd__a31o_1
XFILLER_69_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5209_ _5202_/A _5202_/B _5195_/Y vssd1 vssd1 vccd1 vccd1 _5212_/A sky130_fd_sc_hd__o21ai_4
XFILLER_29_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5560_ _5560_/A _5560_/B vssd1 vssd1 vccd1 vccd1 _5604_/A sky130_fd_sc_hd__xnor2_1
X_5491_ _5491_/A _5491_/B vssd1 vssd1 vccd1 vccd1 _6148_/A sky130_fd_sc_hd__xnor2_4
X_4511_ _4511_/A _4511_/B vssd1 vssd1 vccd1 vccd1 _4513_/B sky130_fd_sc_hd__xor2_4
XFILLER_117_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4442_ _4430_/A _4430_/B _7214_/A _4396_/B _4430_/C vssd1 vssd1 vccd1 vccd1 _4442_/X
+ sky130_fd_sc_hd__o221a_1
X_7230_ _7241_/A _7241_/B _7223_/Y vssd1 vssd1 vccd1 vccd1 _7232_/B sky130_fd_sc_hd__a21bo_4
XFILLER_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4373_ _4430_/A _4407_/B vssd1 vssd1 vccd1 vccd1 _4373_/Y sky130_fd_sc_hd__nor2_1
X_7161_ _7161_/A _7161_/B vssd1 vssd1 vccd1 vccd1 _7177_/A sky130_fd_sc_hd__xnor2_4
XFILLER_112_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6112_ _6192_/B _6192_/C _6112_/C vssd1 vssd1 vccd1 vccd1 _6112_/X sky130_fd_sc_hd__or3_2
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7092_ _7094_/A _7092_/B vssd1 vssd1 vccd1 vccd1 _7110_/B sky130_fd_sc_hd__nor2_4
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6043_ _6043_/A _6343_/A vssd1 vssd1 vccd1 vccd1 _6044_/B sky130_fd_sc_hd__nor2_4
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7994_ _8069_/Q _8013_/Q _8004_/S vssd1 vssd1 vccd1 vccd1 _8069_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _7101_/A _7334_/A vssd1 vssd1 vccd1 vccd1 _7072_/A sky130_fd_sc_hd__or2_2
XFILLER_22_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6876_ _6914_/A _6875_/B _6872_/A vssd1 vssd1 vccd1 vccd1 _6877_/B sky130_fd_sc_hd__o21a_1
XFILLER_22_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5827_ _5826_/A _5826_/B _5826_/C vssd1 vssd1 vccd1 vccd1 _5834_/B sky130_fd_sc_hd__a21o_1
X_5758_ _5755_/A _5925_/A _5756_/X _5754_/X vssd1 vssd1 vccd1 vccd1 _5759_/C sky130_fd_sc_hd__o31ai_4
X_4709_ _4708_/B _4709_/B vssd1 vssd1 vccd1 vccd1 _4709_/Y sky130_fd_sc_hd__nand2b_1
X_7428_ _7428_/A _7428_/B vssd1 vssd1 vccd1 vccd1 _7430_/B sky130_fd_sc_hd__nand2_4
X_5689_ _5715_/A _5689_/B vssd1 vssd1 vccd1 vccd1 _5691_/B sky130_fd_sc_hd__nor2_4
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7359_ _7359_/A _7359_/B vssd1 vssd1 vccd1 vccd1 _7363_/B sky130_fd_sc_hd__xor2_1
XFILLER_103_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6730_ _6730_/A vssd1 vssd1 vccd1 vccd1 _6730_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4991_ _4991_/A _5020_/B vssd1 vssd1 vccd1 vccd1 _4992_/B sky130_fd_sc_hd__nand2_4
X_6661_ _6661_/A vssd1 vssd1 vccd1 vccd1 _6661_/Y sky130_fd_sc_hd__inv_2
X_6592_ _6592_/A _6592_/B vssd1 vssd1 vccd1 vccd1 _6613_/B sky130_fd_sc_hd__xnor2_4
X_5612_ _5612_/A _5612_/B _5612_/C vssd1 vssd1 vccd1 vccd1 _5613_/B sky130_fd_sc_hd__nand3_1
X_5543_ _5596_/A _5596_/B vssd1 vssd1 vccd1 vccd1 _5548_/A sky130_fd_sc_hd__nand2b_2
X_5474_ _5474_/A _5474_/B vssd1 vssd1 vccd1 vccd1 _5477_/C sky130_fd_sc_hd__xnor2_2
X_7213_ _7213_/A _7213_/B _7213_/C vssd1 vssd1 vccd1 vccd1 _7285_/C sky130_fd_sc_hd__and3_4
X_4425_ _4360_/A _4423_/X _4424_/Y _4416_/Y _4421_/X vssd1 vssd1 vccd1 vccd1 _4425_/X
+ sky130_fd_sc_hd__o32a_1
X_4356_ _4356_/A _4356_/B vssd1 vssd1 vccd1 vccd1 _4356_/Y sky130_fd_sc_hd__nand2_1
X_7144_ _7134_/X _7158_/B _7133_/X vssd1 vssd1 vccd1 vccd1 _7146_/B sky130_fd_sc_hd__o21ba_4
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4287_ _4212_/Y _5989_/B _4246_/X _4548_/B vssd1 vssd1 vccd1 vccd1 _4287_/X sky130_fd_sc_hd__o211a_2
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7075_ _7076_/A _7076_/B vssd1 vssd1 vccd1 vccd1 _7081_/B sky130_fd_sc_hd__nand2_1
X_6026_ _5996_/A _6027_/A _7413_/A vssd1 vssd1 vccd1 vccd1 _6026_/X sky130_fd_sc_hd__a21o_2
XFILLER_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7977_ _8013_/Q _8053_/Q _7986_/S vssd1 vssd1 vccd1 vccd1 _8053_/D sky130_fd_sc_hd__mux2_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout22 _7581_/S vssd1 vssd1 vccd1 vccd1 _6753_/S sky130_fd_sc_hd__buf_4
Xfanout11 _6254_/S vssd1 vssd1 vccd1 vccd1 _7570_/B sky130_fd_sc_hd__buf_4
X_6928_ _6940_/A _6940_/B vssd1 vssd1 vccd1 vccd1 _6931_/C sky130_fd_sc_hd__nor2_1
Xfanout33 _6590_/B vssd1 vssd1 vccd1 vccd1 _6688_/S sky130_fd_sc_hd__clkbuf_4
X_6859_ _6862_/A _6862_/B _6858_/A vssd1 vssd1 vccd1 vccd1 _6861_/B sky130_fd_sc_hd__a21o_2
Xfanout55 _4868_/D vssd1 vssd1 vccd1 vccd1 _4947_/C sky130_fd_sc_hd__buf_4
Xfanout44 _5342_/B vssd1 vssd1 vccd1 vccd1 _5672_/A sky130_fd_sc_hd__buf_8
Xfanout99 _6445_/S vssd1 vssd1 vccd1 vccd1 _6456_/S sky130_fd_sc_hd__buf_6
Xfanout77 _7294_/B vssd1 vssd1 vccd1 vccd1 _5800_/A sky130_fd_sc_hd__buf_6
Xfanout88 _5089_/X vssd1 vssd1 vccd1 vccd1 _7195_/B sky130_fd_sc_hd__buf_8
Xfanout66 _6791_/A vssd1 vssd1 vccd1 vccd1 _7150_/B sky130_fd_sc_hd__buf_12
XFILLER_13_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4210_ _4210_/A _4210_/B _4210_/C vssd1 vssd1 vccd1 vccd1 _4241_/B sky130_fd_sc_hd__nand3_4
XFILLER_79_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5190_ _5722_/A _5722_/B vssd1 vssd1 vccd1 vccd1 _5516_/A sky130_fd_sc_hd__nand2_4
XFILLER_95_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4141_ _8067_/Q _8068_/Q _8070_/Q _8069_/Q vssd1 vssd1 vccd1 vccd1 _4147_/A sky130_fd_sc_hd__or4_4
XFILLER_110_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4072_ _8063_/Q _4072_/B vssd1 vssd1 vccd1 vccd1 _6289_/A sky130_fd_sc_hd__xnor2_4
XFILLER_95_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7900_ _7900_/A _7900_/B vssd1 vssd1 vccd1 vccd1 _7900_/X sky130_fd_sc_hd__or2_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7831_ _7831_/A _7831_/B vssd1 vssd1 vccd1 vccd1 _7834_/B sky130_fd_sc_hd__and2_1
XFILLER_51_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7762_ _7728_/A _7759_/Y _7760_/X _6269_/X vssd1 vssd1 vccd1 vccd1 _7763_/B sky130_fd_sc_hd__a31o_1
XFILLER_63_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4974_ _4974_/A _4974_/B vssd1 vssd1 vccd1 vccd1 _4980_/B sky130_fd_sc_hd__xnor2_4
XFILLER_17_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6713_ _6697_/X _6712_/X _6713_/S vssd1 vssd1 vccd1 vccd1 _6713_/X sky130_fd_sc_hd__mux2_1
X_7693_ _6268_/X _7674_/Y _7683_/X _7692_/X _7903_/B1 vssd1 vssd1 vccd1 vccd1 _7693_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_6644_ _6642_/X _6654_/B _6695_/S vssd1 vssd1 vccd1 vccd1 _6645_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6575_ _6310_/A _5985_/X _6766_/S vssd1 vssd1 vccd1 vccd1 _6580_/B sky130_fd_sc_hd__mux2_8
XFILLER_117_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5526_ _5526_/A _5526_/B vssd1 vssd1 vccd1 vccd1 _5561_/A sky130_fd_sc_hd__xor2_4
X_5457_ _5450_/A _5450_/B _5448_/Y vssd1 vssd1 vccd1 vccd1 _5474_/A sky130_fd_sc_hd__a21bo_4
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4408_ _4407_/A _4407_/B _4430_/A vssd1 vssd1 vccd1 vccd1 _4408_/Y sky130_fd_sc_hd__a21oi_1
Xfanout223 _6522_/S vssd1 vssd1 vccd1 vccd1 _6544_/S sky130_fd_sc_hd__buf_8
Xfanout201 _4087_/A vssd1 vssd1 vccd1 vccd1 _6272_/A sky130_fd_sc_hd__buf_12
XFILLER_87_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout212 _4228_/A vssd1 vssd1 vccd1 vccd1 _4216_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_59_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5388_ _6970_/A _5388_/B vssd1 vssd1 vccd1 vccd1 _5389_/B sky130_fd_sc_hd__xor2_4
XFILLER_115_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout234 _8051_/Q vssd1 vssd1 vccd1 vccd1 _4088_/A sky130_fd_sc_hd__buf_6
XFILLER_59_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4339_ _4376_/B _4376_/C vssd1 vssd1 vccd1 vccd1 _4339_/Y sky130_fd_sc_hd__nor2_1
X_7127_ _7127_/A _7127_/B vssd1 vssd1 vccd1 vccd1 _7128_/B sky130_fd_sc_hd__xnor2_4
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7058_ _7281_/B _7195_/B vssd1 vssd1 vccd1 vccd1 _7072_/B sky130_fd_sc_hd__nand2_2
X_6009_ _6009_/A _7400_/A vssd1 vssd1 vccd1 vccd1 _6009_/X sky130_fd_sc_hd__xor2_4
XFILLER_74_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4690_ _4690_/A _4712_/A vssd1 vssd1 vccd1 vccd1 _4690_/Y sky130_fd_sc_hd__nor2_1
X_6360_ _5745_/A _6916_/A _6445_/S vssd1 vssd1 vccd1 vccd1 _6360_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5311_ _5311_/A _5311_/B vssd1 vssd1 vccd1 vccd1 _5504_/B sky130_fd_sc_hd__xnor2_4
XFILLER_115_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8030_ _8063_/CLK _8030_/D vssd1 vssd1 vccd1 vccd1 _8030_/Q sky130_fd_sc_hd__dfxtp_1
X_6291_ _6289_/A _6289_/B _6273_/B _6273_/A _6290_/X vssd1 vssd1 vccd1 vccd1 _6291_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5242_ _5352_/A _5352_/B _5842_/B vssd1 vssd1 vccd1 vccd1 _5407_/A sky130_fd_sc_hd__and3_4
XFILLER_69_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5173_ _5232_/B _5175_/B vssd1 vssd1 vccd1 vccd1 _5176_/A sky130_fd_sc_hd__or2_2
XFILLER_110_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4124_ _4098_/B _5134_/A2 _4123_/X _4303_/B vssd1 vssd1 vccd1 vccd1 _4124_/X sky130_fd_sc_hd__a211o_2
XFILLER_110_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput1 io_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_4
X_4055_ _6272_/A _4055_/B vssd1 vssd1 vccd1 vccd1 _4117_/B sky130_fd_sc_hd__nor2_2
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7814_ _7874_/A _7874_/B _7837_/A vssd1 vssd1 vccd1 vccd1 _7814_/X sky130_fd_sc_hd__o21a_1
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7745_ _7837_/A _7764_/A vssd1 vssd1 vccd1 vccd1 _7750_/A sky130_fd_sc_hd__nand2_1
XFILLER_61_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4957_ _4957_/A _4957_/B vssd1 vssd1 vccd1 vccd1 _4959_/A sky130_fd_sc_hd__xnor2_4
X_7676_ _6757_/C _7894_/B _7718_/S vssd1 vssd1 vccd1 vccd1 _7677_/C sky130_fd_sc_hd__mux2_2
X_4888_ _5189_/B _4888_/B vssd1 vssd1 vccd1 vccd1 _5247_/A sky130_fd_sc_hd__or2_4
X_6627_ _6627_/A _6627_/B vssd1 vssd1 vccd1 vccd1 _6628_/B sky130_fd_sc_hd__and2_1
X_6558_ _6559_/A _6565_/A vssd1 vssd1 vccd1 vccd1 _6626_/B sky130_fd_sc_hd__nor2_2
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6489_ _6452_/Y _6488_/Y _6364_/A _6413_/B vssd1 vssd1 vccd1 vccd1 _6584_/A sky130_fd_sc_hd__o2bb2a_2
XFILLER_3_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5509_ _5745_/A _5714_/A _5714_/C vssd1 vssd1 vccd1 vccd1 _5566_/A sky130_fd_sc_hd__and3_4
XFILLER_105_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5860_ _5859_/A _5881_/D _5825_/A vssd1 vssd1 vccd1 vccd1 _5885_/B sky130_fd_sc_hd__o21a_1
XFILLER_34_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4811_ _4813_/B _4816_/A _4813_/A vssd1 vssd1 vccd1 vccd1 _4814_/A sky130_fd_sc_hd__o21a_1
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5791_ _6971_/B _5880_/A vssd1 vssd1 vccd1 vccd1 _5822_/B sky130_fd_sc_hd__or2_2
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7530_ _7525_/A _7529_/X _7526_/X vssd1 vssd1 vccd1 vccd1 _7530_/X sky130_fd_sc_hd__a21o_1
X_4742_ _5019_/A _5020_/A _5090_/B vssd1 vssd1 vccd1 vccd1 _4874_/A sky130_fd_sc_hd__and3_1
XFILLER_119_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7461_ _7451_/X _7460_/X _7535_/A vssd1 vssd1 vccd1 vccd1 _7537_/B sky130_fd_sc_hd__mux2_1
X_4673_ _4673_/A _4673_/B _4673_/C vssd1 vssd1 vccd1 vccd1 _4690_/A sky130_fd_sc_hd__and3_2
X_6412_ _6371_/B _6453_/B _6441_/S vssd1 vssd1 vccd1 vccd1 _6413_/B sky130_fd_sc_hd__mux2_1
X_7392_ _7392_/A _7392_/B _7392_/C vssd1 vssd1 vccd1 vccd1 _7392_/X sky130_fd_sc_hd__or3_1
XFILLER_115_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6343_ _6343_/A _6343_/B vssd1 vssd1 vccd1 vccd1 _6343_/Y sky130_fd_sc_hd__xnor2_1
X_6274_ _6274_/A _6274_/B vssd1 vssd1 vccd1 vccd1 _6274_/Y sky130_fd_sc_hd__nor2_1
X_8013_ _8079_/CLK _8013_/D vssd1 vssd1 vccd1 vccd1 _8013_/Q sky130_fd_sc_hd__dfxtp_2
X_5225_ _5227_/A _5227_/B _5166_/X vssd1 vssd1 vccd1 vccd1 _5957_/A sky130_fd_sc_hd__o21bai_4
XFILLER_102_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5156_ _6806_/A _5244_/A _5156_/C vssd1 vssd1 vccd1 vccd1 _5227_/A sky130_fd_sc_hd__or3_4
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4107_ _4107_/A _4107_/B vssd1 vssd1 vccd1 vccd1 _4107_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5087_ _5322_/A _5087_/B _5268_/B vssd1 vssd1 vccd1 vccd1 _5087_/X sky130_fd_sc_hd__and3_2
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4038_ _7974_/A _4038_/B vssd1 vssd1 vccd1 vccd1 _8027_/D sky130_fd_sc_hd__and2b_1
XFILLER_72_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _6272_/B _5989_/B vssd1 vssd1 vccd1 vccd1 _6017_/B sky130_fd_sc_hd__xnor2_4
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7728_ _7728_/A _7728_/B vssd1 vssd1 vccd1 vccd1 _7728_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7659_ _7542_/B _7658_/Y _7847_/A vssd1 vssd1 vccd1 vccd1 _7687_/B sky130_fd_sc_hd__mux2_4
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5010_ _5010_/A _5010_/B vssd1 vssd1 vccd1 vccd1 _5030_/A sky130_fd_sc_hd__xnor2_4
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6961_ _6961_/A vssd1 vssd1 vccd1 vccd1 _6996_/B sky130_fd_sc_hd__inv_2
XFILLER_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6892_ _6892_/A _6892_/B vssd1 vssd1 vccd1 vccd1 _7387_/B sky130_fd_sc_hd__xor2_1
XFILLER_34_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5912_ _5912_/A _5912_/B _5912_/C vssd1 vssd1 vccd1 vccd1 _5914_/A sky130_fd_sc_hd__and3_1
XFILLER_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5843_ _5843_/A _5843_/B vssd1 vssd1 vccd1 vccd1 _5850_/B sky130_fd_sc_hd__xnor2_2
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7513_ _7512_/Y _7508_/X _7513_/S vssd1 vssd1 vccd1 vccd1 _7513_/X sky130_fd_sc_hd__mux2_1
X_5774_ _5774_/A vssd1 vssd1 vccd1 vccd1 _5804_/B sky130_fd_sc_hd__inv_2
X_4725_ _4726_/B _4725_/B vssd1 vssd1 vccd1 vccd1 _4837_/B sky130_fd_sc_hd__or2_1
XFILLER_107_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7444_ _7441_/X _7443_/X _7483_/S vssd1 vssd1 vccd1 vccd1 _7444_/X sky130_fd_sc_hd__mux2_1
X_4656_ _4663_/A _4663_/B vssd1 vssd1 vccd1 vccd1 _4664_/A sky130_fd_sc_hd__nand2_1
X_7375_ _7517_/A _7512_/B _7362_/X vssd1 vssd1 vccd1 vccd1 _7508_/B sky130_fd_sc_hd__a21o_1
X_4587_ _4587_/A _4587_/B vssd1 vssd1 vccd1 vccd1 _4589_/B sky130_fd_sc_hd__and2_2
X_6326_ _6326_/A _6326_/B vssd1 vssd1 vccd1 vccd1 _6336_/A sky130_fd_sc_hd__nor2_1
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6257_ _6166_/X _6226_/X _6255_/Y _6256_/X _7784_/A vssd1 vssd1 vccd1 vccd1 _6258_/D
+ sky130_fd_sc_hd__o41a_1
XFILLER_67_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6188_ _6188_/A _6770_/A vssd1 vssd1 vccd1 vccd1 _7886_/A sky130_fd_sc_hd__xnor2_4
X_5208_ _5208_/A _5465_/A _6871_/B vssd1 vssd1 vccd1 vccd1 _5265_/A sky130_fd_sc_hd__or3_4
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5139_ _5386_/A _6842_/B vssd1 vssd1 vccd1 vccd1 _5264_/A sky130_fd_sc_hd__or2_4
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5490_ _5490_/A _5490_/B vssd1 vssd1 vccd1 vccd1 _5491_/B sky130_fd_sc_hd__xor2_4
X_4510_ _4511_/A _4511_/B vssd1 vssd1 vccd1 vccd1 _4510_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4441_ _4441_/A _4441_/B vssd1 vssd1 vccd1 vccd1 _4441_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7160_ _7160_/A _7160_/B vssd1 vssd1 vccd1 vccd1 _7181_/A sky130_fd_sc_hd__nand2_4
X_6111_ _6112_/C _6111_/B _6111_/C vssd1 vssd1 vccd1 vccd1 _6219_/A sky130_fd_sc_hd__and3b_1
X_4372_ _4360_/A _7245_/A _4430_/A vssd1 vssd1 vccd1 vccd1 _4372_/X sky130_fd_sc_hd__a21o_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _7091_/A _7091_/B _7091_/C vssd1 vssd1 vccd1 vccd1 _7092_/B sky130_fd_sc_hd__and3_2
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6042_ _6042_/A vssd1 vssd1 vccd1 vccd1 _6044_/A sky130_fd_sc_hd__inv_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7993_ _8068_/Q _8012_/Q _8004_/S vssd1 vssd1 vccd1 vccd1 _8068_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6944_ _7334_/A _7235_/B vssd1 vssd1 vccd1 vccd1 _7114_/C sky130_fd_sc_hd__nor2_2
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6875_ _6875_/A _6875_/B vssd1 vssd1 vccd1 vccd1 _6914_/B sky130_fd_sc_hd__nor2_2
XFILLER_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5826_ _5826_/A _5826_/B _5826_/C vssd1 vssd1 vccd1 vccd1 _5834_/A sky130_fd_sc_hd__nand3_1
XFILLER_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5757_ _5754_/A _5822_/A _5756_/X vssd1 vssd1 vccd1 vccd1 _5790_/B sky130_fd_sc_hd__o21ba_2
X_4708_ _4708_/A _4708_/B vssd1 vssd1 vccd1 vccd1 _4708_/X sky130_fd_sc_hd__or2_2
X_7427_ _7423_/A _7422_/B _6064_/Y _7426_/B _7766_/A vssd1 vssd1 vccd1 vccd1 _7428_/B
+ sky130_fd_sc_hd__a2111o_2
X_5688_ _5688_/A _5688_/B vssd1 vssd1 vccd1 vccd1 _5740_/A sky130_fd_sc_hd__xor2_4
X_4639_ _4639_/A _4639_/B _4639_/C vssd1 vssd1 vccd1 vccd1 _4668_/A sky130_fd_sc_hd__nand3_2
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7358_ _7371_/A _7358_/B vssd1 vssd1 vccd1 vccd1 _7363_/A sky130_fd_sc_hd__or2_1
X_6309_ _6315_/A _6310_/B vssd1 vssd1 vccd1 vccd1 _6309_/Y sky130_fd_sc_hd__nor2_1
X_7289_ _7286_/A _7286_/B _7282_/Y vssd1 vssd1 vccd1 vccd1 _7301_/A sky130_fd_sc_hd__a21bo_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4990_ _4990_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _4992_/A sky130_fd_sc_hd__xor2_4
X_6660_ _6695_/S _6642_/X _6659_/X vssd1 vssd1 vccd1 vccd1 _6661_/A sky130_fd_sc_hd__a21oi_2
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6591_ _6614_/A _6614_/B vssd1 vssd1 vccd1 vccd1 _6615_/A sky130_fd_sc_hd__nand2_2
X_5611_ _5611_/A _5617_/A vssd1 vssd1 vccd1 vccd1 _6118_/A sky130_fd_sc_hd__xnor2_4
X_5542_ _5594_/A _5542_/B vssd1 vssd1 vccd1 vccd1 _5596_/B sky130_fd_sc_hd__xnor2_4
XFILLER_31_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5473_ _5473_/A _5473_/B vssd1 vssd1 vccd1 vccd1 _5474_/B sky130_fd_sc_hd__xnor2_4
X_4424_ _4424_/A _4424_/B vssd1 vssd1 vccd1 vccd1 _4424_/Y sky130_fd_sc_hd__nor2_1
X_7212_ _7212_/A _7212_/B vssd1 vssd1 vccd1 vccd1 _7219_/A sky130_fd_sc_hd__xnor2_2
X_4355_ _4548_/C _4355_/B vssd1 vssd1 vccd1 vccd1 _4355_/Y sky130_fd_sc_hd__nor2_4
X_7143_ _7143_/A _7143_/B vssd1 vssd1 vccd1 vccd1 _7158_/B sky130_fd_sc_hd__xnor2_4
XFILLER_101_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7074_ _7081_/A _7074_/B vssd1 vssd1 vccd1 vccd1 _7076_/B sky130_fd_sc_hd__and2_2
X_4286_ _6035_/A0 _4285_/X _4283_/X vssd1 vssd1 vccd1 vccd1 _4286_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _6043_/A _6025_/B vssd1 vssd1 vccd1 vccd1 _7413_/A sky130_fd_sc_hd__and2_4
XFILLER_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7976_ _8012_/Q _8052_/Q _7986_/S vssd1 vssd1 vccd1 vccd1 _8052_/D sky130_fd_sc_hd__mux2_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout12 _6112_/X vssd1 vssd1 vccd1 vccd1 _6254_/S sky130_fd_sc_hd__buf_4
X_6927_ _6931_/B _6927_/B vssd1 vssd1 vccd1 vccd1 _6940_/B sky130_fd_sc_hd__or2_1
Xfanout23 _6623_/Y vssd1 vssd1 vccd1 vccd1 _7581_/S sky130_fd_sc_hd__clkbuf_4
Xfanout34 _6689_/S vssd1 vssd1 vccd1 vccd1 _6695_/S sky130_fd_sc_hd__buf_4
X_6858_ _6858_/A _6858_/B vssd1 vssd1 vccd1 vccd1 _6862_/B sky130_fd_sc_hd__nor2_2
Xfanout56 _4738_/Y vssd1 vssd1 vccd1 vccd1 _4795_/C sky130_fd_sc_hd__buf_4
Xfanout45 _5243_/A vssd1 vssd1 vccd1 vccd1 _5582_/A sky130_fd_sc_hd__buf_8
Xfanout78 _6917_/B vssd1 vssd1 vccd1 vccd1 _7294_/B sky130_fd_sc_hd__clkbuf_16
Xfanout89 _7124_/A2 vssd1 vssd1 vccd1 vccd1 _5621_/A sky130_fd_sc_hd__buf_6
XFILLER_10_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout67 _4642_/B vssd1 vssd1 vccd1 vccd1 _5013_/B sky130_fd_sc_hd__buf_6
X_5809_ _5811_/A _5811_/B vssd1 vssd1 vccd1 vccd1 _5815_/A sky130_fd_sc_hd__or2_1
X_6789_ _6836_/A _6836_/B vssd1 vssd1 vccd1 vccd1 _6834_/B sky130_fd_sc_hd__and2_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4140_ _8067_/Q _8068_/Q vssd1 vssd1 vccd1 vccd1 _4196_/B sky130_fd_sc_hd__or2_4
XFILLER_68_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4071_ _4087_/A _4071_/B vssd1 vssd1 vccd1 vccd1 _4071_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7830_ _7856_/A _7830_/B vssd1 vssd1 vccd1 vccd1 _8037_/D sky130_fd_sc_hd__nor2_1
XFILLER_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7761_ _7728_/A _7760_/X _7759_/Y vssd1 vssd1 vccd1 vccd1 _7763_/A sky130_fd_sc_hd__a21oi_1
X_4973_ _4968_/A _4968_/B _4969_/B _5020_/B vssd1 vssd1 vccd1 vccd1 _4980_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_36_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6712_ _6697_/S _6651_/Y _6711_/X vssd1 vssd1 vccd1 vccd1 _6712_/X sky130_fd_sc_hd__a21bo_1
X_7692_ _7929_/A _7707_/A _7707_/B _7691_/Y vssd1 vssd1 vccd1 vccd1 _7692_/X sky130_fd_sc_hd__o31a_2
X_6643_ _6554_/B _6581_/A _6688_/S vssd1 vssd1 vccd1 vccd1 _6654_/B sky130_fd_sc_hd__mux2_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6574_ _6588_/S _6555_/A _6573_/Y _6568_/Y _6525_/A vssd1 vssd1 vccd1 vccd1 _6580_/A
+ sky130_fd_sc_hd__o32ai_4
X_5525_ _5526_/A _5526_/B vssd1 vssd1 vccd1 vccd1 _5525_/Y sky130_fd_sc_hd__nor2_2
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5456_ _5612_/A _5612_/B _5612_/C vssd1 vssd1 vccd1 vccd1 _5613_/A sky130_fd_sc_hd__a21o_2
X_4407_ _4407_/A _4407_/B vssd1 vssd1 vccd1 vccd1 _5969_/B sky130_fd_sc_hd__and2_2
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout202 _4087_/A vssd1 vssd1 vccd1 vccd1 _6326_/A sky130_fd_sc_hd__buf_12
XFILLER_87_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout213 _6326_/B vssd1 vssd1 vccd1 vccd1 _4228_/A sky130_fd_sc_hd__buf_6
X_5387_ _6970_/A _5388_/B vssd1 vssd1 vccd1 vccd1 _5387_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout235 _7974_/A vssd1 vssd1 vccd1 vccd1 _7928_/A sky130_fd_sc_hd__buf_4
XFILLER_101_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout224 _6522_/S vssd1 vssd1 vccd1 vccd1 _7607_/A sky130_fd_sc_hd__buf_2
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4338_ _4548_/A _4317_/A _4317_/B _4548_/C vssd1 vssd1 vccd1 vccd1 _4376_/C sky130_fd_sc_hd__a31o_2
X_7126_ _7167_/A _7124_/X _7122_/X vssd1 vssd1 vccd1 vccd1 _7130_/A sky130_fd_sc_hd__o21ai_2
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4269_ _4341_/A1 _4266_/X _4267_/X vssd1 vssd1 vccd1 vccd1 _4483_/A sky130_fd_sc_hd__a21oi_4
X_7057_ _7057_/A _7294_/B vssd1 vssd1 vccd1 vccd1 _7112_/A sky130_fd_sc_hd__nor2_1
XFILLER_101_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6008_ _6009_/A _7400_/A vssd1 vssd1 vccd1 vccd1 _6008_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7959_ _8012_/Q _7961_/A _8045_/Q vssd1 vssd1 vccd1 vccd1 _7960_/B sky130_fd_sc_hd__a21oi_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6290_ _4077_/B _4242_/A _6287_/Y _6288_/X _6289_/X vssd1 vssd1 vccd1 vccd1 _6290_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5310_ _5672_/A _5800_/A vssd1 vssd1 vccd1 vccd1 _5311_/B sky130_fd_sc_hd__or2_4
XFILLER_115_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5241_ _5241_/A _5241_/B vssd1 vssd1 vccd1 vccd1 _5262_/A sky130_fd_sc_hd__xnor2_4
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5172_ _5172_/A _5172_/B vssd1 vssd1 vccd1 vccd1 _5175_/B sky130_fd_sc_hd__nor2_1
XFILLER_68_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4123_ _4074_/Y _4118_/X _4094_/B _4071_/Y vssd1 vssd1 vccd1 vccd1 _4123_/X sky130_fd_sc_hd__o211a_1
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4054_ _8058_/Q _4054_/B vssd1 vssd1 vccd1 vccd1 _4056_/S sky130_fd_sc_hd__xor2_4
Xinput2 io_in[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_2
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7813_ _7887_/A _7837_/B vssd1 vssd1 vccd1 vccd1 _7813_/X sky130_fd_sc_hd__or2_1
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7744_ _7744_/A _7744_/B vssd1 vssd1 vccd1 vccd1 _7764_/A sky130_fd_sc_hd__or2_1
XFILLER_24_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4956_ _4957_/A _4957_/B vssd1 vssd1 vccd1 vccd1 _4956_/X sky130_fd_sc_hd__or2_1
X_7675_ _7583_/S _6748_/X _6631_/X vssd1 vssd1 vccd1 vccd1 _7894_/B sky130_fd_sc_hd__o21ba_1
X_4887_ _4887_/A _4887_/B vssd1 vssd1 vccd1 vccd1 _4888_/B sky130_fd_sc_hd__and2_1
XFILLER_32_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6626_ _6626_/A _6626_/B _6626_/C vssd1 vssd1 vccd1 vccd1 _6627_/B sky130_fd_sc_hd__or3_1
X_6557_ _6564_/A _6697_/S vssd1 vssd1 vccd1 vccd1 _6565_/A sky130_fd_sc_hd__or2_1
XFILLER_20_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5508_ _5714_/A _5714_/C vssd1 vssd1 vccd1 vccd1 _5858_/B sky130_fd_sc_hd__and2_4
XFILLER_105_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6488_ _6488_/A _6488_/B vssd1 vssd1 vccd1 vccd1 _6488_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5439_ _5439_/A _5439_/B vssd1 vssd1 vccd1 vccd1 _5440_/B sky130_fd_sc_hd__xnor2_4
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7109_ _7094_/A _7092_/B _7110_/A vssd1 vssd1 vccd1 vccd1 _7109_/X sky130_fd_sc_hd__o21a_1
XFILLER_59_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4810_ _4832_/A _4815_/B vssd1 vssd1 vccd1 vccd1 _4816_/A sky130_fd_sc_hd__nor2_2
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5790_ _5790_/A _5790_/B vssd1 vssd1 vccd1 vccd1 _5824_/A sky130_fd_sc_hd__xnor2_4
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4773_/A _4989_/A _4795_/C vssd1 vssd1 vccd1 vccd1 _4890_/A sky130_fd_sc_hd__or3_4
X_7460_ _7459_/Y _7456_/X _7624_/S vssd1 vssd1 vccd1 vccd1 _7460_/X sky130_fd_sc_hd__mux2_1
X_4672_ _4673_/A _4673_/B _4673_/C vssd1 vssd1 vccd1 vccd1 _4691_/A sky130_fd_sc_hd__a21o_2
XFILLER_119_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6411_ _6484_/S _6390_/B _6410_/X vssd1 vssd1 vccd1 vccd1 _6453_/B sky130_fd_sc_hd__o21ai_1
X_7391_ _6823_/B _6860_/Y _7452_/A _7452_/B vssd1 vssd1 vccd1 vccd1 _7454_/B sky130_fd_sc_hd__a2bb2o_1
X_6342_ _7413_/A _6342_/B vssd1 vssd1 vccd1 vccd1 _6342_/X sky130_fd_sc_hd__or2_1
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6273_ _6273_/A _6273_/B vssd1 vssd1 vccd1 vccd1 _6273_/X sky130_fd_sc_hd__or2_1
X_8012_ _8057_/CLK _8012_/D vssd1 vssd1 vccd1 vccd1 _8012_/Q sky130_fd_sc_hd__dfxtp_2
X_5224_ _5166_/C _5956_/A _5223_/Y vssd1 vssd1 vccd1 vccd1 _5227_/B sky130_fd_sc_hd__o21ai_4
X_5155_ _5155_/A _5155_/B vssd1 vssd1 vccd1 vccd1 _5160_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4106_ _4088_/A _6060_/A _4084_/X _4087_/X vssd1 vssd1 vccd1 vccd1 _4107_/B sky130_fd_sc_hd__o211a_1
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5086_ _4074_/Y _4118_/X _6018_/A _8051_/Q _4071_/Y vssd1 vssd1 vccd1 vccd1 _5268_/B
+ sky130_fd_sc_hd__o2111a_1
X_4037_ _8027_/Q input2/X _7991_/D vssd1 vssd1 vccd1 vccd1 _4038_/B sky130_fd_sc_hd__mux2_1
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _6310_/A _5987_/B _5985_/X _6011_/B vssd1 vssd1 vccd1 vccd1 _6009_/A sky130_fd_sc_hd__a2bb2o_4
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7727_ _7760_/A _7760_/B _7697_/B vssd1 vssd1 vccd1 vccd1 _7728_/B sky130_fd_sc_hd__or3b_1
X_4939_ _4939_/A _4939_/B vssd1 vssd1 vccd1 vccd1 _4942_/B sky130_fd_sc_hd__nand2_2
X_7658_ _7538_/S _7550_/X _7657_/Y vssd1 vssd1 vccd1 vccd1 _7658_/Y sky130_fd_sc_hd__a21boi_2
X_6609_ _7773_/A _6621_/A vssd1 vssd1 vccd1 vccd1 _6610_/B sky130_fd_sc_hd__nand2_1
X_7589_ _7649_/A _7648_/A _7648_/B vssd1 vssd1 vccd1 vccd1 _7589_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6960_ _6978_/B _6960_/B vssd1 vssd1 vccd1 vccd1 _6961_/A sky130_fd_sc_hd__nand2_1
XFILLER_93_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5911_ _5909_/A _5907_/Y _5916_/A vssd1 vssd1 vccd1 vccd1 _5912_/C sky130_fd_sc_hd__o21ai_1
X_6891_ _6893_/A _6893_/B vssd1 vssd1 vccd1 vccd1 _6892_/B sky130_fd_sc_hd__nand2b_2
XFILLER_46_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5842_ _5908_/A _5842_/B _5908_/C vssd1 vssd1 vccd1 vccd1 _5850_/A sky130_fd_sc_hd__and3_1
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5773_ _5798_/B _5772_/Y _5808_/A vssd1 vssd1 vccd1 vccd1 _5774_/A sky130_fd_sc_hd__a21oi_1
X_7512_ _7512_/A _7512_/B vssd1 vssd1 vccd1 vccd1 _7512_/Y sky130_fd_sc_hd__xnor2_1
X_4724_ _7281_/A _5034_/A _4718_/C vssd1 vssd1 vccd1 vccd1 _4725_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7443_ _7440_/X _7442_/X _7479_/S vssd1 vssd1 vccd1 vccd1 _7443_/X sky130_fd_sc_hd__mux2_1
X_4655_ _7247_/A _5013_/A vssd1 vssd1 vccd1 vccd1 _4663_/B sky130_fd_sc_hd__nor2_2
X_7374_ _7374_/A _7374_/B vssd1 vssd1 vccd1 vccd1 _7512_/B sky130_fd_sc_hd__xnor2_2
X_4586_ _4551_/A _4551_/B _4552_/A _4551_/D vssd1 vssd1 vccd1 vccd1 _4587_/B sky130_fd_sc_hd__a22o_1
X_6325_ _7413_/A _6342_/B vssd1 vssd1 vccd1 vccd1 _6325_/Y sky130_fd_sc_hd__nand2_1
X_6256_ _6211_/X _6212_/X _6225_/X vssd1 vssd1 vccd1 vccd1 _6256_/X sky130_fd_sc_hd__a21bo_1
X_6187_ _6188_/A _6770_/A vssd1 vssd1 vccd1 vccd1 _6187_/X sky130_fd_sc_hd__xor2_4
XFILLER_97_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5207_ _5207_/A _5800_/A vssd1 vssd1 vccd1 vccd1 _6871_/B sky130_fd_sc_hd__or2_4
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5138_ _6842_/B vssd1 vssd1 vccd1 vccd1 _5842_/B sky130_fd_sc_hd__clkinv_4
X_5069_ _5977_/A _5065_/Y _5066_/Y _5068_/Y vssd1 vssd1 vccd1 vccd1 _6791_/A sky130_fd_sc_hd__o31a_4
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4440_ _4360_/A _4439_/X _4438_/X _4494_/A vssd1 vssd1 vccd1 vccd1 _4440_/X sky130_fd_sc_hd__a211o_2
X_6110_ _6110_/A _6259_/B vssd1 vssd1 vccd1 vccd1 _6112_/C sky130_fd_sc_hd__xnor2_1
X_4371_ _7245_/A _4407_/A _4360_/A vssd1 vssd1 vccd1 vccd1 _4371_/X sky130_fd_sc_hd__a21o_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7090_ _7090_/A _7090_/B vssd1 vssd1 vccd1 vccd1 _7110_/A sky130_fd_sc_hd__xnor2_4
X_6041_ _6043_/A _6343_/A vssd1 vssd1 vccd1 vccd1 _6042_/A sky130_fd_sc_hd__nand2_2
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7992_ _8067_/Q _8011_/Q _8004_/S vssd1 vssd1 vccd1 vccd1 _8067_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6943_ _6943_/A _6943_/B vssd1 vssd1 vccd1 vccd1 _6943_/X sky130_fd_sc_hd__xor2_1
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6874_ _6916_/A _7281_/C _5275_/C vssd1 vssd1 vccd1 vccd1 _6875_/B sky130_fd_sc_hd__a21oi_2
X_5825_ _5825_/A _5885_/A _5862_/A vssd1 vssd1 vccd1 vccd1 _5826_/C sky130_fd_sc_hd__nor3_2
X_5756_ _5800_/A _5880_/A _5714_/X vssd1 vssd1 vccd1 vccd1 _5756_/X sky130_fd_sc_hd__o21ba_2
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5687_ _5688_/A _5688_/B vssd1 vssd1 vccd1 vccd1 _5687_/Y sky130_fd_sc_hd__nand2_1
X_4707_ _4708_/A _4708_/B vssd1 vssd1 vccd1 vccd1 _4707_/Y sky130_fd_sc_hd__nor2_1
X_7426_ _7426_/A _7426_/B _7426_/C vssd1 vssd1 vccd1 vccd1 _7428_/A sky130_fd_sc_hd__nand3_2
X_4638_ _4638_/A _4638_/B vssd1 vssd1 vccd1 vccd1 _4639_/C sky130_fd_sc_hd__xor2_4
XFILLER_118_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7357_ _7370_/A _7369_/A vssd1 vssd1 vccd1 vccd1 _7359_/B sky130_fd_sc_hd__nand2_1
X_4569_ _4570_/B _4570_/A vssd1 vssd1 vccd1 vccd1 _4569_/X sky130_fd_sc_hd__and2b_2
XFILLER_116_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6308_ _6308_/A _6308_/B vssd1 vssd1 vccd1 vccd1 _6626_/A sky130_fd_sc_hd__xnor2_2
XFILLER_103_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7288_ _7290_/A _7290_/B vssd1 vssd1 vccd1 vccd1 _7288_/Y sky130_fd_sc_hd__nor2_1
X_6239_ _6241_/A _6239_/B vssd1 vssd1 vccd1 vccd1 _6240_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6590_ _6590_/A _6590_/B vssd1 vssd1 vccd1 vccd1 _6614_/B sky130_fd_sc_hd__xor2_2
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5610_ _5611_/A _5617_/A vssd1 vssd1 vccd1 vccd1 _5610_/Y sky130_fd_sc_hd__nand2_1
X_5541_ _5541_/A _5853_/B vssd1 vssd1 vccd1 vccd1 _5596_/A sky130_fd_sc_hd__or2_4
X_7211_ _7211_/A _7211_/B vssd1 vssd1 vccd1 vccd1 _7212_/B sky130_fd_sc_hd__xnor2_4
X_5472_ _5473_/B _5473_/A vssd1 vssd1 vccd1 vccd1 _5472_/X sky130_fd_sc_hd__and2b_1
X_4423_ _4370_/Y _4422_/Y _4424_/A vssd1 vssd1 vccd1 vccd1 _4423_/X sky130_fd_sc_hd__o21a_1
X_4354_ _4354_/A _4354_/B vssd1 vssd1 vccd1 vccd1 _4354_/X sky130_fd_sc_hd__or2_2
X_7142_ _7142_/A _7142_/B vssd1 vssd1 vccd1 vccd1 _7143_/B sky130_fd_sc_hd__xor2_4
XFILLER_98_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7073_ _7072_/A _7072_/B _7072_/C vssd1 vssd1 vccd1 vccd1 _7074_/B sky130_fd_sc_hd__o21ai_1
X_6024_ _6024_/A _6024_/B vssd1 vssd1 vccd1 vccd1 _6025_/B sky130_fd_sc_hd__nand2_1
X_4285_ _4219_/Y _4244_/B _4284_/X vssd1 vssd1 vccd1 vccd1 _4285_/X sky130_fd_sc_hd__o21a_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7975_ _8011_/Q _4088_/A _7986_/S vssd1 vssd1 vccd1 vccd1 _8051_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6926_ _6909_/B _6926_/B vssd1 vssd1 vccd1 vccd1 _6927_/B sky130_fd_sc_hd__and2b_1
Xfanout13 _6219_/A vssd1 vssd1 vccd1 vccd1 _6193_/A sky130_fd_sc_hd__buf_4
Xfanout35 _6580_/A vssd1 vssd1 vccd1 vccd1 _6689_/S sky130_fd_sc_hd__buf_2
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout24 _7502_/B vssd1 vssd1 vccd1 vccd1 _7527_/S sky130_fd_sc_hd__buf_4
X_6857_ _6857_/A _6857_/B _6857_/C vssd1 vssd1 vccd1 vccd1 _6858_/B sky130_fd_sc_hd__and3_1
Xfanout46 _5338_/B vssd1 vssd1 vccd1 vccd1 _5723_/A sky130_fd_sc_hd__clkbuf_16
Xfanout68 _5541_/A vssd1 vssd1 vccd1 vccd1 _6806_/A sky130_fd_sc_hd__buf_8
X_6788_ _6788_/A _6788_/B vssd1 vssd1 vccd1 vccd1 _6836_/B sky130_fd_sc_hd__xnor2_2
Xfanout79 _5204_/X vssd1 vssd1 vccd1 vccd1 _7281_/C sky130_fd_sc_hd__buf_12
XFILLER_50_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout57 _4738_/Y vssd1 vssd1 vccd1 vccd1 _4751_/C sky130_fd_sc_hd__buf_8
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5808_ _5808_/A _5808_/B vssd1 vssd1 vccd1 vccd1 _5811_/B sky130_fd_sc_hd__xnor2_4
X_5739_ _5776_/A _5776_/B _5731_/Y vssd1 vssd1 vccd1 vccd1 _5741_/A sky130_fd_sc_hd__a21o_4
XFILLER_108_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7409_ _7949_/B _6805_/B _6304_/A _6065_/B _7426_/B vssd1 vssd1 vccd1 vccd1 _7766_/A
+ sky130_fd_sc_hd__o32a_4
XFILLER_116_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4070_ _6060_/A _4071_/B vssd1 vssd1 vccd1 vccd1 _4111_/A sky130_fd_sc_hd__xnor2_4
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7760_ _7760_/A _7760_/B _7733_/X _7697_/B vssd1 vssd1 vccd1 vccd1 _7760_/X sky130_fd_sc_hd__or4bb_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4972_ _4974_/A _4974_/B vssd1 vssd1 vccd1 vccd1 _4979_/A sky130_fd_sc_hd__nand2_1
XFILLER_17_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6711_ _6709_/Y _6710_/X _6691_/A _6679_/B vssd1 vssd1 vccd1 vccd1 _6711_/X sky130_fd_sc_hd__a2bb2o_1
X_7691_ _7918_/B _7691_/B vssd1 vssd1 vccd1 vccd1 _7691_/Y sky130_fd_sc_hd__nor2_1
X_6642_ _6547_/A _6547_/B _6737_/B vssd1 vssd1 vccd1 vccd1 _6642_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6573_ _6571_/B _6570_/Y _6572_/Y _6555_/B vssd1 vssd1 vccd1 vccd1 _6573_/Y sky130_fd_sc_hd__a31oi_4
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5524_ _5562_/A _5562_/B _5523_/A vssd1 vssd1 vccd1 vccd1 _5526_/B sky130_fd_sc_hd__a21oi_4
XFILLER_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5455_ _5455_/A _5455_/B vssd1 vssd1 vccd1 vccd1 _5612_/C sky130_fd_sc_hd__xor2_1
XFILLER_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4406_ _4406_/A _4472_/A _7245_/A vssd1 vssd1 vccd1 vccd1 _4406_/X sky130_fd_sc_hd__or3_1
Xfanout203 _4046_/Y vssd1 vssd1 vccd1 vccd1 _4087_/A sky130_fd_sc_hd__buf_8
Xfanout214 _4149_/Y vssd1 vssd1 vccd1 vccd1 _6326_/B sky130_fd_sc_hd__clkbuf_16
X_5386_ _5386_/A _5797_/A vssd1 vssd1 vccd1 vccd1 _5388_/B sky130_fd_sc_hd__nor2_4
X_7125_ _7122_/A _7216_/A _7124_/X vssd1 vssd1 vccd1 vccd1 _7167_/B sky130_fd_sc_hd__o21ba_2
XFILLER_115_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout236 _7974_/A vssd1 vssd1 vccd1 vccd1 _7856_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout225 _6187_/X vssd1 vssd1 vccd1 vccd1 _6522_/S sky130_fd_sc_hd__clkbuf_4
X_4337_ _4548_/A _4317_/A _4317_/B _4354_/A vssd1 vssd1 vccd1 vccd1 _4340_/B sky130_fd_sc_hd__a31oi_4
X_4268_ _4341_/A1 _4266_/A _4266_/B _4267_/X vssd1 vssd1 vccd1 vccd1 _4268_/X sky130_fd_sc_hd__a31o_1
X_7056_ _7056_/A _7056_/B vssd1 vssd1 vccd1 vccd1 _7063_/A sky130_fd_sc_hd__xor2_4
X_6007_ _6007_/A _6317_/A vssd1 vssd1 vccd1 vccd1 _7400_/A sky130_fd_sc_hd__xor2_4
XFILLER_67_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4199_ _8070_/Q _4199_/B vssd1 vssd1 vccd1 vccd1 _4199_/X sky130_fd_sc_hd__xor2_4
XFILLER_55_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7958_ _7974_/A _7991_/C _7991_/D vssd1 vssd1 vccd1 vccd1 _7961_/B sky130_fd_sc_hd__or3b_2
XFILLER_82_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7889_ _7889_/A _7889_/B vssd1 vssd1 vccd1 vccd1 _7913_/B sky130_fd_sc_hd__nor2_4
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6909_ _6926_/B _6909_/B vssd1 vssd1 vccd1 vccd1 _6931_/B sky130_fd_sc_hd__and2b_1
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5240_ _5240_/A _5240_/B vssd1 vssd1 vccd1 vccd1 _5280_/A sky130_fd_sc_hd__xnor2_2
XFILLER_114_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5171_ _5172_/A _5172_/B vssd1 vssd1 vccd1 vccd1 _5232_/B sky130_fd_sc_hd__and2_1
XFILLER_68_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4122_ _4074_/Y _4118_/X _6278_/A _4071_/Y vssd1 vssd1 vccd1 vccd1 _4122_/X sky130_fd_sc_hd__o211a_1
XFILLER_68_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4053_ _8058_/Q _4054_/B vssd1 vssd1 vccd1 vccd1 _4053_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_56_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput3 io_in[2] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
X_7812_ _7887_/A _7837_/B vssd1 vssd1 vccd1 vccd1 _7812_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7743_ _7743_/A _7743_/B vssd1 vssd1 vccd1 vccd1 _7743_/Y sky130_fd_sc_hd__nand2_1
X_4955_ _5019_/A _5040_/B vssd1 vssd1 vccd1 vccd1 _4990_/A sky130_fd_sc_hd__nand2_2
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7674_ _7760_/A _7674_/B vssd1 vssd1 vccd1 vccd1 _7674_/Y sky130_fd_sc_hd__xnor2_4
X_4886_ _4887_/A _4887_/B vssd1 vssd1 vccd1 vccd1 _5189_/B sky130_fd_sc_hd__nor2_4
X_6625_ _6616_/X _6619_/Y _7773_/A vssd1 vssd1 vccd1 vccd1 _6628_/A sky130_fd_sc_hd__o21ai_1
X_6556_ _6588_/S _6556_/B vssd1 vssd1 vccd1 vccd1 _6697_/S sky130_fd_sc_hd__nor2_8
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5507_ _5047_/B _5047_/C _5047_/A vssd1 vssd1 vccd1 vccd1 _5714_/C sky130_fd_sc_hd__o21ai_4
X_6487_ _6374_/A _6386_/B _6486_/Y _6443_/A vssd1 vssd1 vccd1 vccd1 _6549_/A sky130_fd_sc_hd__a22o_4
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5438_ _5439_/A _5439_/B vssd1 vssd1 vccd1 vccd1 _5438_/X sky130_fd_sc_hd__and2b_1
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5369_ _5369_/A _5369_/B vssd1 vssd1 vccd1 vccd1 _5377_/A sky130_fd_sc_hd__nand2_4
X_7108_ _7108_/A _7108_/B vssd1 vssd1 vccd1 vccd1 _7151_/A sky130_fd_sc_hd__xnor2_4
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7039_ _7039_/A _7054_/A vssd1 vssd1 vccd1 vccd1 _7041_/B sky130_fd_sc_hd__and2_2
XFILLER_90_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4998_/A _5090_/B vssd1 vssd1 vccd1 vccd1 _4746_/A sky130_fd_sc_hd__nand2_2
X_4671_ _4670_/A _4670_/C _4670_/B vssd1 vssd1 vccd1 vccd1 _4673_/C sky130_fd_sc_hd__a21bo_1
X_6410_ _6451_/A _6410_/B vssd1 vssd1 vccd1 vccd1 _6410_/X sky130_fd_sc_hd__or2_1
X_7390_ _6833_/A _6823_/B _6860_/Y _7389_/Y vssd1 vssd1 vccd1 vccd1 _7452_/B sky130_fd_sc_hd__a31oi_4
X_6341_ _7420_/A _6341_/B vssd1 vssd1 vccd1 vccd1 _6341_/Y sky130_fd_sc_hd__xnor2_2
X_6272_ _6272_/A _6272_/B vssd1 vssd1 vccd1 vccd1 _6272_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8011_ _8075_/CLK _8011_/D vssd1 vssd1 vccd1 vccd1 _8011_/Q sky130_fd_sc_hd__dfxtp_2
X_5223_ _6805_/B _5386_/A _5164_/X vssd1 vssd1 vccd1 vccd1 _5223_/Y sky130_fd_sc_hd__o21ai_2
X_5154_ _5154_/A _5154_/B vssd1 vssd1 vccd1 vccd1 _5180_/A sky130_fd_sc_hd__xor2_2
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4105_ _4080_/C _4103_/X _4081_/B vssd1 vssd1 vccd1 vccd1 _6030_/A sky130_fd_sc_hd__a21o_4
XFILLER_84_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5085_ _5083_/X _5084_/X _5087_/B vssd1 vssd1 vccd1 vccd1 _5085_/X sky130_fd_sc_hd__a21o_1
X_4036_ _8025_/Q _8026_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _8026_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5987_ _6315_/A _5987_/B vssd1 vssd1 vccd1 vccd1 _6011_/B sky130_fd_sc_hd__xnor2_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7726_ _7724_/X _7725_/Y _7928_/A vssd1 vssd1 vccd1 vccd1 _8033_/D sky130_fd_sc_hd__a21oi_1
X_4938_ _4938_/A _4938_/B vssd1 vssd1 vccd1 vccd1 _4939_/B sky130_fd_sc_hd__or2_1
X_7657_ _7657_/A _7657_/B vssd1 vssd1 vccd1 vccd1 _7657_/Y sky130_fd_sc_hd__nand2_1
X_4869_ _4868_/B _4868_/C _4868_/D _4991_/A vssd1 vssd1 vccd1 vccd1 _4870_/B sky130_fd_sc_hd__a22o_1
X_6608_ _7773_/A _6621_/A vssd1 vssd1 vccd1 vccd1 _6608_/X sky130_fd_sc_hd__and2_1
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7588_ _7649_/A _7648_/A _7648_/B vssd1 vssd1 vccd1 vccd1 _7588_/X sky130_fd_sc_hd__or3_1
X_6539_ _6539_/A _6539_/B _6539_/C vssd1 vssd1 vccd1 vccd1 _6540_/B sky130_fd_sc_hd__or3_1
XFILLER_106_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5910_ _5915_/A _5915_/B vssd1 vssd1 vccd1 vccd1 _5916_/A sky130_fd_sc_hd__nand2_1
X_6890_ _6888_/A _6888_/B _6895_/A vssd1 vssd1 vccd1 vccd1 _6893_/B sky130_fd_sc_hd__o21ai_4
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5841_ _5843_/B _5843_/A vssd1 vssd1 vccd1 vccd1 _5841_/X sky130_fd_sc_hd__and2b_1
X_5772_ _5691_/B _5768_/Y _5771_/B vssd1 vssd1 vccd1 vccd1 _5772_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7511_ _7506_/X _7510_/X _7515_/S vssd1 vssd1 vccd1 vccd1 _7534_/B sky130_fd_sc_hd__mux2_1
X_4723_ _5013_/B _7001_/A _4716_/B vssd1 vssd1 vccd1 vccd1 _4837_/A sky130_fd_sc_hd__or3b_1
XFILLER_21_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7442_ _7442_/A _7442_/B vssd1 vssd1 vccd1 vccd1 _7442_/X sky130_fd_sc_hd__xor2_1
X_4654_ _4654_/A _5013_/A vssd1 vssd1 vccd1 vccd1 _4716_/B sky130_fd_sc_hd__nor2_1
X_7373_ _7512_/A vssd1 vssd1 vccd1 vccd1 _7517_/A sky130_fd_sc_hd__inv_2
X_4585_ _7281_/A _4585_/B _5019_/A _7281_/B vssd1 vssd1 vccd1 vccd1 _4627_/A sky130_fd_sc_hd__and4_4
X_6324_ _6564_/A _6327_/B _6320_/B _7398_/A vssd1 vssd1 vccd1 vccd1 _6342_/B sky130_fd_sc_hd__a2bb2o_2
X_6255_ _6255_/A _6255_/B _6255_/C _6255_/D vssd1 vssd1 vccd1 vccd1 _6255_/Y sky130_fd_sc_hd__nand4_1
XFILLER_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5206_ _5386_/A _6917_/B vssd1 vssd1 vccd1 vccd1 _5464_/B sky130_fd_sc_hd__nor2_2
X_6186_ _6166_/X _7784_/B _7784_/A vssd1 vssd1 vccd1 vccd1 _7611_/D sky130_fd_sc_hd__mux2_8
XFILLER_69_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5137_ _5977_/B _5133_/Y _5136_/Y _5322_/A vssd1 vssd1 vccd1 vccd1 _5137_/X sky130_fd_sc_hd__a211o_4
XFILLER_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5068_ _5322_/A _5362_/B vssd1 vssd1 vccd1 vccd1 _5068_/Y sky130_fd_sc_hd__nand2_2
XFILLER_57_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4019_ _7562_/B _7879_/B vssd1 vssd1 vccd1 vccd1 _4020_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7709_ _7709_/A vssd1 vssd1 vccd1 vccd1 _7709_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ _7165_/A _4412_/B vssd1 vssd1 vccd1 vccd1 _4370_/Y sky130_fd_sc_hd__nor2_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6343_/A vssd1 vssd1 vccd1 vccd1 _7416_/A sky130_fd_sc_hd__inv_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7991_ _7974_/A _8008_/Q _7991_/C _7991_/D vssd1 vssd1 vccd1 vccd1 _7991_/X sky130_fd_sc_hd__and4b_1
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6942_ _6942_/A _6942_/B vssd1 vssd1 vccd1 vccd1 _6978_/A sky130_fd_sc_hd__xor2_2
XFILLER_81_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6873_ _6873_/A _6873_/B vssd1 vssd1 vccd1 vccd1 _6914_/A sky130_fd_sc_hd__nand2_4
XFILLER_62_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5824_ _5824_/A _5824_/B vssd1 vssd1 vccd1 vccd1 _5862_/A sky130_fd_sc_hd__xnor2_4
X_5755_ _5755_/A _5925_/A vssd1 vssd1 vccd1 vccd1 _5790_/A sky130_fd_sc_hd__or2_4
X_5686_ _5686_/A _5686_/B vssd1 vssd1 vccd1 vccd1 _5688_/B sky130_fd_sc_hd__xor2_4
X_4706_ _4611_/X _4704_/Y _4700_/A _4695_/X vssd1 vssd1 vccd1 vccd1 _4708_/B sky130_fd_sc_hd__o211a_1
XFILLER_108_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7425_ _7423_/A _7422_/B _6065_/A vssd1 vssd1 vccd1 vccd1 _7426_/C sky130_fd_sc_hd__a21bo_1
X_4637_ _4636_/B _4636_/C _4660_/A vssd1 vssd1 vccd1 vccd1 _4639_/B sky130_fd_sc_hd__a21o_1
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7356_ _7356_/A vssd1 vssd1 vccd1 vccd1 _7369_/A sky130_fd_sc_hd__inv_2
X_4568_ _4561_/A _4561_/C _4561_/B vssd1 vssd1 vccd1 vccd1 _4570_/B sky130_fd_sc_hd__a21boi_4
X_6307_ _6308_/A _6559_/A vssd1 vssd1 vccd1 vccd1 _6601_/B sky130_fd_sc_hd__nand2_2
XFILLER_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7287_ _7302_/A _7302_/B vssd1 vssd1 vccd1 vccd1 _7290_/B sky130_fd_sc_hd__or2_4
XFILLER_1_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4499_ _4461_/A _4461_/B _4467_/X vssd1 vssd1 vccd1 vccd1 _4513_/A sky130_fd_sc_hd__a21o_2
XFILLER_89_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6238_ _6238_/A _6238_/B _6237_/X vssd1 vssd1 vccd1 vccd1 _6238_/X sky130_fd_sc_hd__or3b_1
X_6169_ _6081_/B _6134_/A _6262_/S _7755_/A vssd1 vssd1 vccd1 vccd1 _6169_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5540_ _5549_/A _5549_/B vssd1 vssd1 vccd1 vccd1 _5540_/Y sky130_fd_sc_hd__nor2_1
X_5471_ _5471_/A _5471_/B vssd1 vssd1 vccd1 vccd1 _5473_/B sky130_fd_sc_hd__xnor2_4
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7210_ _7245_/A _7210_/B _7244_/A vssd1 vssd1 vccd1 vccd1 _7220_/B sky130_fd_sc_hd__or3_2
X_4422_ _4441_/A _7214_/A _4662_/A vssd1 vssd1 vccd1 vccd1 _4422_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_98_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4353_ _4354_/A _4354_/B vssd1 vssd1 vccd1 vccd1 _4353_/Y sky130_fd_sc_hd__nor2_2
X_7141_ _7141_/A _7141_/B vssd1 vssd1 vccd1 vccd1 _7142_/B sky130_fd_sc_hd__xnor2_4
XFILLER_101_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4284_ _4170_/X _4259_/B _4236_/X _4315_/B vssd1 vssd1 vccd1 vccd1 _4284_/X sky130_fd_sc_hd__a211o_1
X_7072_ _7072_/A _7072_/B _7072_/C vssd1 vssd1 vccd1 vccd1 _7081_/A sky130_fd_sc_hd__or3_1
X_6023_ _6024_/A _6024_/B vssd1 vssd1 vccd1 vccd1 _6043_/A sky130_fd_sc_hd__or2_4
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7974_ _7974_/A _8008_/Q _7974_/C _7991_/D vssd1 vssd1 vccd1 vccd1 _7974_/X sky130_fd_sc_hd__or4b_4
XFILLER_82_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6925_ _6925_/A _6925_/B vssd1 vssd1 vccd1 vccd1 _6940_/A sky130_fd_sc_hd__xnor2_1
XFILLER_22_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout36 _6641_/B vssd1 vssd1 vccd1 vccd1 _6691_/A sky130_fd_sc_hd__buf_4
Xfanout14 _7930_/A vssd1 vssd1 vccd1 vccd1 _7784_/A sky130_fd_sc_hd__clkbuf_16
Xfanout25 _7483_/S vssd1 vssd1 vccd1 vccd1 _7502_/B sky130_fd_sc_hd__buf_6
X_6856_ _6857_/B _6857_/C _6857_/A vssd1 vssd1 vccd1 vccd1 _6858_/A sky130_fd_sc_hd__a21oi_2
XFILLER_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout47 _5689_/B vssd1 vssd1 vccd1 vccd1 _5853_/B sky130_fd_sc_hd__buf_6
Xfanout69 _7101_/A vssd1 vssd1 vccd1 vccd1 _5541_/A sky130_fd_sc_hd__buf_12
X_6787_ _6806_/A _7030_/A vssd1 vssd1 vccd1 vccd1 _6836_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout58 _5041_/D1 vssd1 vssd1 vccd1 vccd1 _5020_/B sky130_fd_sc_hd__clkbuf_16
X_5807_ _5840_/A _5840_/B _5805_/Y vssd1 vssd1 vccd1 vccd1 _5811_/A sky130_fd_sc_hd__a21boi_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5738_ _5779_/A _5738_/B vssd1 vssd1 vccd1 vccd1 _5776_/B sky130_fd_sc_hd__nor2_4
XFILLER_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5669_ _5670_/B _5669_/B vssd1 vssd1 vccd1 vccd1 _5671_/A sky130_fd_sc_hd__and2b_2
X_7408_ _7420_/A _7420_/B _6055_/A vssd1 vssd1 vccd1 vccd1 _7426_/B sky130_fd_sc_hd__a21o_2
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7339_ _7352_/A _7352_/B vssd1 vssd1 vccd1 vccd1 _7340_/B sky130_fd_sc_hd__nand2_4
XFILLER_104_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4971_ _4971_/A _4971_/B vssd1 vssd1 vccd1 vccd1 _4974_/B sky130_fd_sc_hd__xor2_4
X_6710_ _6524_/B _6737_/B _6688_/X _6695_/S _6691_/A vssd1 vssd1 vccd1 vccd1 _6710_/X
+ sky130_fd_sc_hd__a221o_1
X_7690_ _7929_/A _7707_/A _7707_/B vssd1 vssd1 vccd1 vccd1 _7691_/B sky130_fd_sc_hd__o21a_1
XFILLER_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6641_ _6697_/S _6641_/B vssd1 vssd1 vccd1 vccd1 _6645_/A sky130_fd_sc_hd__or2_1
XFILLER_20_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6572_ _6572_/A _6572_/B vssd1 vssd1 vccd1 vccd1 _6572_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5523_ _5523_/A _5523_/B vssd1 vssd1 vccd1 vccd1 _5562_/B sky130_fd_sc_hd__nor2_4
X_5454_ _5455_/B _5455_/A vssd1 vssd1 vccd1 vccd1 _5477_/B sky130_fd_sc_hd__nand2b_1
X_5385_ _5445_/A _7344_/B vssd1 vssd1 vccd1 vccd1 _6916_/C sky130_fd_sc_hd__nor2_8
X_4405_ _4436_/A _7165_/A vssd1 vssd1 vccd1 vccd1 _4405_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout204 _8007_/S vssd1 vssd1 vccd1 vccd1 _8004_/S sky130_fd_sc_hd__buf_6
X_4336_ _4312_/B _4312_/C _4548_/A vssd1 vssd1 vccd1 vccd1 _4340_/A sky130_fd_sc_hd__a21o_1
X_7124_ _4654_/A _7124_/A2 _7247_/C _7214_/A vssd1 vssd1 vccd1 vccd1 _7124_/X sky130_fd_sc_hd__o22a_1
Xfanout215 _4020_/X vssd1 vssd1 vccd1 vccd1 _7955_/S sky130_fd_sc_hd__buf_6
Xfanout237 input4/X vssd1 vssd1 vccd1 vccd1 _7974_/A sky130_fd_sc_hd__clkbuf_4
Xfanout226 _4147_/A vssd1 vssd1 vccd1 vccd1 _4175_/B sky130_fd_sc_hd__buf_6
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4267_ _4315_/A _4548_/B _5989_/B _4548_/A vssd1 vssd1 vccd1 vccd1 _4267_/X sky130_fd_sc_hd__o31a_4
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7055_ _7055_/A _7055_/B vssd1 vssd1 vccd1 vccd1 _7091_/A sky130_fd_sc_hd__xnor2_4
XFILLER_101_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6006_ _6317_/A _6007_/A vssd1 vssd1 vccd1 vccd1 _6006_/X sky130_fd_sc_hd__and2b_2
X_4198_ _8070_/Q _4199_/B vssd1 vssd1 vccd1 vccd1 _6278_/B sky130_fd_sc_hd__xnor2_4
X_7957_ _7974_/C vssd1 vssd1 vccd1 vccd1 _7991_/C sky130_fd_sc_hd__inv_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7888_ _7888_/A _7888_/B vssd1 vssd1 vccd1 vccd1 _7888_/Y sky130_fd_sc_hd__xnor2_1
X_6908_ _7150_/B _6900_/X _6942_/A _6906_/X vssd1 vssd1 vccd1 vccd1 _6926_/B sky130_fd_sc_hd__o22a_1
X_6839_ _7025_/A _6839_/B _6871_/B vssd1 vssd1 vccd1 vccd1 _6843_/A sky130_fd_sc_hd__or3_2
XFILLER_24_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5170_ _5232_/A _5170_/B vssd1 vssd1 vccd1 vccd1 _5172_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4121_ _4078_/A _4119_/Y _4111_/A vssd1 vssd1 vccd1 vccd1 _4121_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4052_ _4096_/A _4052_/B vssd1 vssd1 vccd1 vccd1 _4054_/B sky130_fd_sc_hd__and2_2
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 rst vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7811_ _7833_/A _7833_/B _7833_/C _7810_/Y vssd1 vssd1 vccd1 vccd1 _7837_/B sky130_fd_sc_hd__a31oi_4
XFILLER_91_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7742_ _7741_/A _7741_/B _6774_/X vssd1 vssd1 vccd1 vccd1 _7743_/B sky130_fd_sc_hd__a21oi_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4954_ _5020_/A _5034_/B vssd1 vssd1 vccd1 vccd1 _4957_/B sky130_fd_sc_hd__nand2_4
X_7673_ _7929_/A _7697_/B vssd1 vssd1 vccd1 vccd1 _7674_/B sky130_fd_sc_hd__or2_4
XFILLER_60_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4885_ _4911_/A _4911_/B _4882_/Y vssd1 vssd1 vccd1 vccd1 _4887_/B sky130_fd_sc_hd__a21boi_4
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6624_ _6733_/S _7581_/S _6616_/X vssd1 vssd1 vccd1 vccd1 _6629_/A sky130_fd_sc_hd__or3b_1
XFILLER_20_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6555_ _6555_/A _6555_/B vssd1 vssd1 vccd1 vccd1 _6556_/B sky130_fd_sc_hd__nor2_4
X_5506_ _5666_/A _5432_/A _5505_/X vssd1 vssd1 vccd1 vccd1 _5522_/A sky130_fd_sc_hd__a21o_1
X_6486_ _6492_/A _6423_/Y _6485_/Y vssd1 vssd1 vccd1 vccd1 _6486_/Y sky130_fd_sc_hd__a21oi_1
X_5437_ _5437_/A _5437_/B vssd1 vssd1 vccd1 vccd1 _5439_/B sky130_fd_sc_hd__xor2_4
XFILLER_99_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5368_ _5386_/A _5683_/B vssd1 vssd1 vccd1 vccd1 _5542_/B sky130_fd_sc_hd__nor2_4
XFILLER_114_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4319_ _4548_/A _4319_/B vssd1 vssd1 vccd1 vccd1 _4355_/B sky130_fd_sc_hd__or2_2
X_5299_ _5299_/A _5714_/A vssd1 vssd1 vccd1 vccd1 _5299_/X sky130_fd_sc_hd__and2_1
X_7107_ _7107_/A _7107_/B vssd1 vssd1 vccd1 vccd1 _7154_/A sky130_fd_sc_hd__xnor2_1
XFILLER_101_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7038_ _7053_/A _7053_/B vssd1 vssd1 vccd1 vccd1 _7054_/A sky130_fd_sc_hd__or2_1
XFILLER_28_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4670_ _4670_/A _4670_/B _4670_/C vssd1 vssd1 vccd1 vccd1 _4689_/A sky130_fd_sc_hd__nand3_1
X_6340_ _6303_/B _6338_/X _6339_/Y _6341_/B _6058_/B vssd1 vssd1 vccd1 vccd1 _6340_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_6_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6271_ _6272_/A _6272_/B vssd1 vssd1 vccd1 vccd1 _6271_/Y sky130_fd_sc_hd__nand2_1
X_8010_ _8080_/CLK _8010_/D vssd1 vssd1 vccd1 vccd1 _8010_/Q sky130_fd_sc_hd__dfxtp_4
X_5222_ _5284_/A _5284_/B vssd1 vssd1 vccd1 vccd1 _5285_/A sky130_fd_sc_hd__or2_4
X_5153_ _5114_/X _5152_/B _5154_/A _5154_/B vssd1 vssd1 vccd1 vccd1 _5179_/A sky130_fd_sc_hd__a22o_1
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4104_ _4080_/C _4103_/X _4081_/B vssd1 vssd1 vccd1 vccd1 _5268_/A sky130_fd_sc_hd__a21oi_4
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5084_ _4087_/B _5993_/B _4305_/X _5135_/C1 vssd1 vssd1 vccd1 vccd1 _5084_/X sky130_fd_sc_hd__a211o_4
XFILLER_56_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4035_ _8024_/Q _8025_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _8025_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5986_ _5271_/B _5984_/B _5986_/S vssd1 vssd1 vccd1 vccd1 _6310_/B sky130_fd_sc_hd__mux2_8
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7725_ _8032_/Q _4018_/X _7857_/B _8033_/Q vssd1 vssd1 vccd1 vccd1 _7725_/Y sky130_fd_sc_hd__a22oi_1
X_4937_ _4971_/A _4971_/B _4928_/X vssd1 vssd1 vccd1 vccd1 _4942_/A sky130_fd_sc_hd__a21oi_4
X_7656_ _7656_/A _7656_/B vssd1 vssd1 vccd1 vccd1 _7684_/A sky130_fd_sc_hd__nand2_1
X_4868_ _4991_/A _4868_/B _4868_/C _4868_/D vssd1 vssd1 vccd1 vccd1 _4874_/B sky130_fd_sc_hd__and4_1
X_6607_ _7773_/A _6621_/A vssd1 vssd1 vccd1 vccd1 _6610_/A sky130_fd_sc_hd__or2_1
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7587_ _7620_/A _7587_/B vssd1 vssd1 vccd1 vccd1 _7648_/B sky130_fd_sc_hd__nand2_1
X_4799_ _4820_/S _4798_/A _4923_/B vssd1 vssd1 vccd1 vccd1 _4800_/B sky130_fd_sc_hd__o21ai_2
XFILLER_20_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6538_ _6538_/A _6538_/B vssd1 vssd1 vccd1 vccd1 _6539_/C sky130_fd_sc_hd__or2_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6469_ _6467_/Y _6472_/B _6366_/Y vssd1 vssd1 vccd1 vccd1 _6469_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5840_ _5840_/A _5840_/B vssd1 vssd1 vccd1 vccd1 _5843_/B sky130_fd_sc_hd__xnor2_2
X_5771_ _5798_/B _5771_/B vssd1 vssd1 vccd1 vccd1 _5808_/A sky130_fd_sc_hd__and2b_4
X_7510_ _7509_/X _7489_/X _7527_/S vssd1 vssd1 vccd1 vccd1 _7510_/X sky130_fd_sc_hd__mux2_1
X_4722_ _4720_/A _4720_/B _4720_/C vssd1 vssd1 vccd1 vccd1 _4728_/B sky130_fd_sc_hd__a21o_1
X_7441_ _7439_/X _7440_/X _7479_/S vssd1 vssd1 vccd1 vccd1 _7441_/X sky130_fd_sc_hd__mux2_1
X_4653_ _4652_/B _4652_/C _4652_/A vssd1 vssd1 vccd1 vccd1 _4673_/B sky130_fd_sc_hd__a21o_1
X_7372_ _7516_/B _7516_/C _7516_/A vssd1 vssd1 vccd1 vccd1 _7512_/A sky130_fd_sc_hd__a21o_1
X_4584_ _5019_/A _7281_/B vssd1 vssd1 vccd1 vccd1 _4675_/A sky130_fd_sc_hd__nand2_1
X_6323_ _5996_/B _5996_/A _6766_/S vssd1 vssd1 vccd1 vccd1 _6327_/B sky130_fd_sc_hd__mux2_2
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6254_ _6248_/X _6253_/X _6254_/S vssd1 vssd1 vccd1 vccd1 _6258_/C sky130_fd_sc_hd__mux2_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5205_ _7213_/A _7170_/B vssd1 vssd1 vccd1 vccd1 _6917_/B sky130_fd_sc_hd__nand2_8
XFILLER_97_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6185_ _6170_/X _6184_/X _6225_/S vssd1 vssd1 vccd1 vccd1 _7784_/B sky130_fd_sc_hd__mux2_1
XFILLER_97_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5136_ _5977_/C _5977_/D _5977_/B vssd1 vssd1 vccd1 vccd1 _5136_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_29_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5067_ _8051_/Q _4303_/C _4126_/X _5087_/B _5135_/C1 vssd1 vssd1 vccd1 vccd1 _5362_/B
+ sky130_fd_sc_hd__o2111a_2
X_4018_ _7562_/B _7964_/C vssd1 vssd1 vccd1 vccd1 _4018_/X sky130_fd_sc_hd__and2_4
XFILLER_65_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5969_ _4360_/Y _5969_/B _5969_/C vssd1 vssd1 vccd1 vccd1 _5969_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7708_ _7538_/S _7592_/B _7657_/Y vssd1 vssd1 vccd1 vccd1 _7709_/A sky130_fd_sc_hd__a21boi_1
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7639_ _7639_/A _7639_/B vssd1 vssd1 vccd1 vccd1 _7639_/Y sky130_fd_sc_hd__nand2_4
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7990_ _8026_/Q _4066_/A _7990_/S vssd1 vssd1 vccd1 vccd1 _8066_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6941_ _6931_/C _6941_/B vssd1 vssd1 vccd1 vccd1 _6983_/A sky130_fd_sc_hd__nand2b_2
XFILLER_81_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6872_ _6872_/A vssd1 vssd1 vccd1 vccd1 _6875_/A sky130_fd_sc_hd__inv_2
XFILLER_62_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5823_ _5824_/B _5823_/B vssd1 vssd1 vccd1 vccd1 _5885_/A sky130_fd_sc_hd__or2_2
X_5754_ _5754_/A _5822_/A vssd1 vssd1 vccd1 vccd1 _5754_/X sky130_fd_sc_hd__or2_2
X_5685_ _5730_/A _5730_/B _5680_/Y vssd1 vssd1 vccd1 vccd1 _5688_/A sky130_fd_sc_hd__a21o_4
X_4705_ _4695_/X _4700_/A _4704_/Y _4611_/X vssd1 vssd1 vccd1 vccd1 _4708_/A sky130_fd_sc_hd__a211oi_4
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7424_ _7424_/A _7424_/B vssd1 vssd1 vccd1 vccd1 _7430_/A sky130_fd_sc_hd__nand2_4
X_4636_ _4660_/A _4636_/B _4636_/C vssd1 vssd1 vccd1 vccd1 _4639_/A sky130_fd_sc_hd__nand3_2
XFILLER_116_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7355_ _7366_/C _7367_/A _7365_/B vssd1 vssd1 vccd1 vccd1 _7356_/A sky130_fd_sc_hd__or3_1
XFILLER_116_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6306_ _6308_/B vssd1 vssd1 vccd1 vccd1 _6559_/A sky130_fd_sc_hd__clkinv_2
X_4567_ _4566_/A _4566_/C _4566_/B vssd1 vssd1 vccd1 vccd1 _4574_/B sky130_fd_sc_hd__a21oi_4
XFILLER_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7286_ _7286_/A _7286_/B vssd1 vssd1 vccd1 vccd1 _7302_/B sky130_fd_sc_hd__xnor2_4
X_4498_ _4497_/A _4498_/B vssd1 vssd1 vccd1 vccd1 _4521_/A sky130_fd_sc_hd__and2b_2
XFILLER_89_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6237_ _6236_/X _5931_/Y _6237_/S vssd1 vssd1 vccd1 vccd1 _6237_/X sky130_fd_sc_hd__mux2_1
X_6168_ _6012_/B _6262_/S _6167_/X vssd1 vssd1 vccd1 vccd1 _6168_/X sky130_fd_sc_hd__o21a_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _5093_/A _5093_/B _5118_/X _4757_/B vssd1 vssd1 vccd1 vccd1 _5119_/X sky130_fd_sc_hd__o211a_1
X_6099_ _6099_/A _6099_/B vssd1 vssd1 vccd1 vccd1 _6259_/C sky130_fd_sc_hd__nand2_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5470_ _5470_/A _5470_/B vssd1 vssd1 vccd1 vccd1 _5471_/B sky130_fd_sc_hd__xnor2_4
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4421_ _4472_/A _4472_/B _4418_/X _4420_/X _7085_/A vssd1 vssd1 vccd1 vccd1 _4421_/X
+ sky130_fd_sc_hd__a311o_1
X_4352_ _8081_/Q _4352_/B vssd1 vssd1 vccd1 vccd1 _4352_/Y sky130_fd_sc_hd__nor2_8
X_7140_ _7128_/A _7128_/B _7129_/X vssd1 vssd1 vccd1 vccd1 _7142_/A sky130_fd_sc_hd__a21o_4
XFILLER_98_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4283_ _4281_/X _4282_/X _4341_/A1 vssd1 vssd1 vccd1 vccd1 _4283_/X sky130_fd_sc_hd__a21o_1
X_7071_ _7071_/A _7071_/B vssd1 vssd1 vccd1 vccd1 _7072_/C sky130_fd_sc_hd__or2_1
XFILLER_101_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6022_ _6024_/A _6024_/B vssd1 vssd1 vccd1 vccd1 _6022_/X sky130_fd_sc_hd__and2b_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7973_ _8050_/Q _7970_/X _7972_/X vssd1 vssd1 vccd1 vccd1 _8050_/D sky130_fd_sc_hd__o21ba_1
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6924_ _6964_/A _6964_/B _6921_/Y vssd1 vssd1 vccd1 vccd1 _6925_/B sky130_fd_sc_hd__a21bo_1
XFILLER_81_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout37 _6562_/Y vssd1 vssd1 vccd1 vccd1 _6641_/B sky130_fd_sc_hd__clkbuf_4
Xfanout15 _6107_/X vssd1 vssd1 vccd1 vccd1 _7930_/A sky130_fd_sc_hd__buf_6
Xfanout26 _7624_/S vssd1 vssd1 vccd1 vccd1 _7515_/S sky130_fd_sc_hd__buf_4
X_6855_ _7057_/A _7046_/B _6903_/A vssd1 vssd1 vccd1 vccd1 _6857_/C sky130_fd_sc_hd__or3_2
X_6786_ _6788_/B _6788_/A vssd1 vssd1 vccd1 vccd1 _6834_/A sky130_fd_sc_hd__and2b_1
Xfanout59 _4842_/X vssd1 vssd1 vccd1 vccd1 _5041_/D1 sky130_fd_sc_hd__buf_4
XFILLER_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout48 _5647_/B vssd1 vssd1 vccd1 vccd1 _5855_/B sky130_fd_sc_hd__buf_4
X_5806_ _5806_/A _5806_/B vssd1 vssd1 vccd1 vccd1 _5840_/B sky130_fd_sc_hd__xnor2_4
XFILLER_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5737_ _5695_/A _5733_/Y _5771_/B vssd1 vssd1 vccd1 vccd1 _5738_/B sky130_fd_sc_hd__a21boi_2
X_7407_ _6343_/A _7416_/B _6039_/A vssd1 vssd1 vccd1 vccd1 _7420_/B sky130_fd_sc_hd__a21o_2
X_5668_ _5666_/A _5666_/B _5713_/A _5713_/B vssd1 vssd1 vccd1 vccd1 _5669_/B sky130_fd_sc_hd__o2bb2ai_1
X_5599_ _5650_/A _5599_/B vssd1 vssd1 vccd1 vccd1 _5618_/A sky130_fd_sc_hd__xnor2_4
X_4619_ _4620_/A _4619_/B _4619_/C vssd1 vssd1 vccd1 vccd1 _4625_/A sky130_fd_sc_hd__nand3_4
X_7338_ _7354_/A _7338_/B vssd1 vssd1 vccd1 vccd1 _7352_/B sky130_fd_sc_hd__xnor2_4
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7269_ _7319_/A _7269_/B vssd1 vssd1 vccd1 vccd1 _7274_/B sky130_fd_sc_hd__nand2_2
XFILLER_92_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4970_ _5003_/A _5003_/B _4964_/X vssd1 vssd1 vccd1 vccd1 _4974_/A sky130_fd_sc_hd__a21o_2
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6640_ _6640_/A vssd1 vssd1 vccd1 vccd1 _7580_/B sky130_fd_sc_hd__inv_2
X_6571_ _7728_/A _6571_/B vssd1 vssd1 vccd1 vccd1 _6572_/B sky130_fd_sc_hd__nand2_2
X_5522_ _5522_/A _5522_/B vssd1 vssd1 vccd1 vccd1 _5523_/B sky130_fd_sc_hd__and2_1
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5453_ _5453_/A _5453_/B vssd1 vssd1 vccd1 vccd1 _5455_/B sky130_fd_sc_hd__xnor2_1
X_4404_ _4377_/A _4397_/Y _4403_/X _4360_/A vssd1 vssd1 vccd1 vccd1 _4404_/Y sky130_fd_sc_hd__o31ai_2
X_5384_ _6800_/B _5855_/B vssd1 vssd1 vccd1 vccd1 _5389_/A sky130_fd_sc_hd__or2_4
Xfanout205 _7991_/X vssd1 vssd1 vccd1 vccd1 _8007_/S sky130_fd_sc_hd__buf_4
X_4335_ _4312_/B _4312_/C _4548_/A vssd1 vssd1 vccd1 vccd1 _4376_/B sky130_fd_sc_hd__a21oi_2
X_7123_ _7123_/A _7281_/D vssd1 vssd1 vccd1 vccd1 _7167_/A sky130_fd_sc_hd__nand2_4
Xfanout227 _7879_/B vssd1 vssd1 vccd1 vccd1 _7964_/C sky130_fd_sc_hd__buf_4
XFILLER_115_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout216 _4020_/X vssd1 vssd1 vccd1 vccd1 _4036_/S sky130_fd_sc_hd__buf_4
Xfanout238 _7991_/D vssd1 vssd1 vccd1 vccd1 _7562_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4266_ _4266_/A _4266_/B vssd1 vssd1 vccd1 vccd1 _4266_/X sky130_fd_sc_hd__and2_2
X_7054_ _7054_/A _7054_/B vssd1 vssd1 vccd1 vccd1 _7097_/A sky130_fd_sc_hd__and2_2
X_4197_ _8069_/Q _4196_/B _4211_/B vssd1 vssd1 vccd1 vccd1 _4199_/B sky130_fd_sc_hd__o21a_4
X_6005_ _6007_/A _6317_/A vssd1 vssd1 vccd1 vccd1 _6005_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_27_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7956_ _8049_/Q _7956_/B _7956_/C _8050_/Q vssd1 vssd1 vccd1 vccd1 _7974_/C sky130_fd_sc_hd__or4b_2
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7887_ _7887_/A _7887_/B _7910_/C vssd1 vssd1 vccd1 vccd1 _7888_/B sky130_fd_sc_hd__or3b_1
XFILLER_70_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6907_ _7150_/B _6900_/X _6906_/X vssd1 vssd1 vccd1 vccd1 _6942_/B sky130_fd_sc_hd__o21ba_1
X_6838_ _6838_/A _6838_/B vssd1 vssd1 vccd1 vccd1 _6845_/A sky130_fd_sc_hd__nor2_4
XFILLER_50_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6769_ _7579_/A _7935_/A _7579_/B vssd1 vssd1 vccd1 vccd1 _6776_/A sky130_fd_sc_hd__o21ai_1
XFILLER_109_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4120_ _4078_/A _4119_/Y _4111_/A vssd1 vssd1 vccd1 vccd1 _4303_/C sky130_fd_sc_hd__a21oi_4
XFILLER_110_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4051_ _6272_/A _4055_/B vssd1 vssd1 vccd1 vccd1 _4117_/A sky130_fd_sc_hd__and2_2
XFILLER_110_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7810_ _7833_/A _7833_/B _7809_/X vssd1 vssd1 vccd1 vccd1 _7810_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_64_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7741_ _7741_/A _7741_/B vssd1 vssd1 vccd1 vccd1 _7743_/A sky130_fd_sc_hd__or2_1
XFILLER_101_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4953_ _4960_/A _4960_/B vssd1 vssd1 vccd1 vccd1 _4953_/X sky130_fd_sc_hd__and2_1
X_7672_ _7576_/A _7569_/C _7576_/Y _7612_/X _7644_/Y vssd1 vssd1 vccd1 vccd1 _7697_/B
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6623_ _6623_/A _6623_/B vssd1 vssd1 vccd1 vccd1 _6623_/Y sky130_fd_sc_hd__nand2_1
X_4884_ _4884_/A _4884_/B vssd1 vssd1 vccd1 vccd1 _4911_/B sky130_fd_sc_hd__xor2_4
X_6554_ _6581_/A _6554_/B vssd1 vssd1 vccd1 vccd1 _6555_/B sky130_fd_sc_hd__nand2_4
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6485_ _6492_/A _6485_/B vssd1 vssd1 vccd1 vccd1 _6485_/Y sky130_fd_sc_hd__nor2_1
X_5505_ _6842_/B _5755_/A _5303_/Y vssd1 vssd1 vccd1 vccd1 _5505_/X sky130_fd_sc_hd__o21ba_1
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5436_ _5191_/X _5338_/Y _5398_/X _5401_/B vssd1 vssd1 vccd1 vccd1 _5439_/A sky130_fd_sc_hd__o22a_4
XFILLER_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5367_ _5367_/A _5647_/B vssd1 vssd1 vccd1 vccd1 _5594_/A sky130_fd_sc_hd__or2_4
XFILLER_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4318_ _4548_/A _4319_/B vssd1 vssd1 vccd1 vccd1 _4356_/B sky130_fd_sc_hd__nor2_1
X_7106_ _7106_/A _7106_/B vssd1 vssd1 vccd1 vccd1 _7439_/A sky130_fd_sc_hd__nand2_1
X_5298_ _5298_/A _5298_/B vssd1 vssd1 vccd1 vccd1 _5314_/A sky130_fd_sc_hd__xnor2_4
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4249_ _4241_/B _4227_/X _4231_/X _4204_/Y vssd1 vssd1 vccd1 vccd1 _4249_/X sky130_fd_sc_hd__o211a_1
X_7037_ _7039_/A _7037_/B vssd1 vssd1 vccd1 vccd1 _7053_/B sky130_fd_sc_hd__nand2_1
XFILLER_47_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7939_ _7939_/A _7939_/B vssd1 vssd1 vccd1 vccd1 _7940_/B sky130_fd_sc_hd__nand2_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6270_ _6267_/B _7568_/B _7611_/D vssd1 vssd1 vccd1 vccd1 _6270_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5221_ _5239_/A _5239_/B _5218_/Y vssd1 vssd1 vccd1 vccd1 _5284_/B sky130_fd_sc_hd__a21oi_1
XFILLER_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5152_ _5183_/A _5152_/B vssd1 vssd1 vccd1 vccd1 _5154_/B sky130_fd_sc_hd__xnor2_2
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4103_ _4103_/A _4107_/A _4088_/X vssd1 vssd1 vccd1 vccd1 _4103_/X sky130_fd_sc_hd__or3b_4
XFILLER_111_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5083_ _6278_/A _5134_/A2 _4292_/X _4303_/B vssd1 vssd1 vccd1 vccd1 _5083_/X sky130_fd_sc_hd__a211o_4
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4034_ _8023_/Q _8024_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _8024_/D sky130_fd_sc_hd__mux2_1
XFILLER_92_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7724_ _7706_/X _7715_/X _7723_/X _7903_/B1 vssd1 vssd1 vccd1 vccd1 _7724_/X sky130_fd_sc_hd__a31o_2
X_5985_ _5986_/S _7213_/C _5984_/Y vssd1 vssd1 vccd1 vccd1 _5985_/X sky130_fd_sc_hd__o21a_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4936_ _4936_/A _4936_/B vssd1 vssd1 vccd1 vccd1 _4971_/B sky130_fd_sc_hd__xnor2_4
X_7655_ _7654_/A _7654_/B _7654_/Y _6774_/X vssd1 vssd1 vccd1 vccd1 _7655_/X sky130_fd_sc_hd__a211o_1
XANTENNA_10 _7085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4867_ _4867_/A _4867_/B vssd1 vssd1 vccd1 vccd1 _4884_/A sky130_fd_sc_hd__and2_2
X_6606_ _6617_/C _6606_/B vssd1 vssd1 vccd1 vccd1 _6621_/A sky130_fd_sc_hd__nor2_2
X_7586_ _7619_/A _7619_/B vssd1 vssd1 vccd1 vccd1 _7587_/B sky130_fd_sc_hd__or2_1
X_6537_ _6538_/B vssd1 vssd1 vccd1 vccd1 _6537_/Y sky130_fd_sc_hd__inv_2
X_4798_ _4798_/A _4820_/S _4923_/B vssd1 vssd1 vccd1 vccd1 _4798_/X sky130_fd_sc_hd__or3b_1
XFILLER_106_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6468_ _6468_/A _6468_/B vssd1 vssd1 vccd1 vccd1 _6472_/B sky130_fd_sc_hd__nand2_2
XFILLER_106_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6399_ _6399_/A _6399_/B vssd1 vssd1 vccd1 vccd1 _6527_/A sky130_fd_sc_hd__nand2_4
X_5419_ _5419_/A _5419_/B vssd1 vssd1 vccd1 vccd1 _5421_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8069_ _8075_/CLK _8069_/D vssd1 vssd1 vccd1 vccd1 _8069_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5770_ _5800_/A _5796_/B _5800_/D vssd1 vssd1 vccd1 vccd1 _5798_/B sky130_fd_sc_hd__or3_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _4720_/A _4720_/B _4720_/C vssd1 vssd1 vccd1 vccd1 _4721_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_21_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7440_ _7440_/A _7440_/B vssd1 vssd1 vccd1 vccd1 _7440_/X sky130_fd_sc_hd__xor2_1
X_4652_ _4652_/A _4652_/B _4652_/C vssd1 vssd1 vccd1 vccd1 _4673_/A sky130_fd_sc_hd__nand3_1
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7371_ _7371_/A _7371_/B _7371_/C vssd1 vssd1 vccd1 vccd1 _7516_/C sky130_fd_sc_hd__or3_1
X_4583_ _4583_/A _4583_/B vssd1 vssd1 vccd1 vccd1 _4614_/A sky130_fd_sc_hd__nor2_4
X_6322_ _7400_/A _6322_/B vssd1 vssd1 vccd1 vccd1 _6488_/A sky130_fd_sc_hd__xnor2_4
X_6253_ _6166_/S _6245_/C _6208_/X _6245_/B vssd1 vssd1 vccd1 vccd1 _6253_/X sky130_fd_sc_hd__a211o_1
XFILLER_88_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5204_ _7213_/A _7170_/B vssd1 vssd1 vccd1 vccd1 _5204_/X sky130_fd_sc_hd__and2_4
XFILLER_97_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6184_ _6179_/X _6183_/X _7570_/B vssd1 vssd1 vccd1 vccd1 _6184_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5135_ _4088_/A _5993_/B _4127_/X _5135_/C1 vssd1 vssd1 vccd1 vccd1 _5977_/D sky130_fd_sc_hd__a211o_4
X_5066_ _5268_/A _5066_/B vssd1 vssd1 vccd1 vccd1 _5066_/Y sky130_fd_sc_hd__nor2_2
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4017_ _8027_/Q input2/X vssd1 vssd1 vccd1 vccd1 _7879_/B sky130_fd_sc_hd__and2b_4
XFILLER_65_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5968_ _4360_/Y _5969_/B _5969_/C vssd1 vssd1 vccd1 vccd1 _6174_/A sky130_fd_sc_hd__and3b_4
X_7707_ _7707_/A _7707_/B vssd1 vssd1 vccd1 vccd1 _7744_/A sky130_fd_sc_hd__nand2_1
X_4919_ _4989_/A _5013_/C _4919_/C vssd1 vssd1 vccd1 vccd1 _4931_/A sky130_fd_sc_hd__or3_4
XFILLER_21_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5899_ _5896_/A _5896_/C _5896_/B vssd1 vssd1 vccd1 vccd1 _5912_/B sky130_fd_sc_hd__o21ai_1
X_7638_ _7928_/A _7638_/B vssd1 vssd1 vccd1 vccd1 _8030_/D sky130_fd_sc_hd__nor2_1
XFILLER_119_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7569_ _7607_/A _7576_/A _7569_/C vssd1 vssd1 vccd1 vccd1 _7577_/A sky130_fd_sc_hd__and3_1
XFILLER_79_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6940_ _6940_/A _6940_/B vssd1 vssd1 vccd1 vccd1 _6941_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6871_ _7025_/A _6871_/B _6871_/C vssd1 vssd1 vccd1 vccd1 _6872_/A sky130_fd_sc_hd__or3_2
X_5822_ _5822_/A _5822_/B vssd1 vssd1 vccd1 vccd1 _5823_/B sky130_fd_sc_hd__and2_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5753_ _7281_/C _5858_/B vssd1 vssd1 vccd1 vccd1 _5822_/A sky130_fd_sc_hd__nand2_2
X_4704_ _4611_/A _4611_/C _4611_/B vssd1 vssd1 vccd1 vccd1 _4704_/Y sky130_fd_sc_hd__a21oi_4
X_5684_ _5684_/A _5684_/B vssd1 vssd1 vccd1 vccd1 _5730_/B sky130_fd_sc_hd__xnor2_4
X_7423_ _7423_/A _7423_/B vssd1 vssd1 vccd1 vccd1 _7424_/B sky130_fd_sc_hd__xnor2_4
XFILLER_8_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4635_ _4641_/B _4634_/C _4634_/A vssd1 vssd1 vccd1 vccd1 _4636_/C sky130_fd_sc_hd__a21o_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7354_ _7354_/A _7354_/B vssd1 vssd1 vccd1 vccd1 _7365_/B sky130_fd_sc_hd__nand2_2
X_4566_ _4566_/A _4566_/B _4566_/C vssd1 vssd1 vccd1 vccd1 _4574_/A sky130_fd_sc_hd__and3_4
X_6305_ _6305_/A _6305_/B vssd1 vssd1 vccd1 vccd1 _6308_/B sky130_fd_sc_hd__xnor2_4
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7285_ _7285_/A _7285_/B _7285_/C vssd1 vssd1 vccd1 vccd1 _7286_/B sky130_fd_sc_hd__and3_4
X_4497_ _4497_/A _4497_/B _4497_/C vssd1 vssd1 vccd1 vccd1 _4498_/B sky130_fd_sc_hd__or3_4
X_6236_ _6236_/A _6236_/B vssd1 vssd1 vccd1 vccd1 _6236_/X sky130_fd_sc_hd__and2_1
X_6167_ _6081_/Y _6111_/B _6111_/C _6009_/X vssd1 vssd1 vccd1 vccd1 _6167_/X sky130_fd_sc_hd__a31o_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _4998_/A _4751_/C _5090_/X vssd1 vssd1 vccd1 vccd1 _5118_/X sky130_fd_sc_hd__a21o_1
X_6098_ _7639_/A _6092_/B _6096_/Y _6092_/A vssd1 vssd1 vccd1 vccd1 _6099_/B sky130_fd_sc_hd__a211o_4
XFILLER_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5049_ _5703_/A _5703_/B vssd1 vssd1 vccd1 vccd1 _5908_/A sky130_fd_sc_hd__or2_4
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4420_ _7165_/A _7319_/A _4268_/X _4377_/A _4436_/A vssd1 vssd1 vccd1 vccd1 _4420_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_99_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4351_ _7136_/A _4349_/Y _4494_/A vssd1 vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__o21ai_4
X_4282_ _4192_/B _4260_/C _4251_/Y _4315_/B vssd1 vssd1 vccd1 vccd1 _4282_/X sky130_fd_sc_hd__a211o_1
X_7070_ _7013_/A _7013_/B _7013_/C vssd1 vssd1 vccd1 vccd1 _7071_/B sky130_fd_sc_hd__a21oi_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6021_ _6021_/A0 _6020_/Y _6021_/S vssd1 vssd1 vccd1 vccd1 _6024_/B sky130_fd_sc_hd__mux2_1
XFILLER_86_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7972_ _8050_/Q _7970_/X _7961_/B _7961_/A vssd1 vssd1 vccd1 vccd1 _7972_/X sky130_fd_sc_hd__a211o_1
XFILLER_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6923_ _6923_/A _6923_/B vssd1 vssd1 vccd1 vccd1 _6964_/B sky130_fd_sc_hd__xnor2_2
Xfanout16 _6635_/Y vssd1 vssd1 vccd1 vccd1 _7894_/A sky130_fd_sc_hd__buf_4
Xfanout27 _7437_/Y vssd1 vssd1 vccd1 vccd1 _7624_/S sky130_fd_sc_hd__buf_6
Xfanout38 _7394_/X vssd1 vssd1 vccd1 vccd1 _7513_/S sky130_fd_sc_hd__buf_6
X_6854_ _7101_/A _7012_/A vssd1 vssd1 vccd1 vccd1 _6903_/A sky130_fd_sc_hd__or2_2
X_6785_ _5275_/A _6783_/B _6838_/A vssd1 vssd1 vccd1 vccd1 _6788_/B sky130_fd_sc_hd__o21ba_1
Xfanout49 _5647_/B vssd1 vssd1 vccd1 vccd1 _5796_/B sky130_fd_sc_hd__clkbuf_4
X_5805_ _5806_/B _5806_/A vssd1 vssd1 vccd1 vccd1 _5805_/Y sky130_fd_sc_hd__nand2b_1
X_5736_ _5736_/A _5736_/B _5736_/C vssd1 vssd1 vccd1 vccd1 _5779_/A sky130_fd_sc_hd__and3_4
XFILLER_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5667_ _5621_/Y _5716_/A _5666_/Y vssd1 vssd1 vccd1 vccd1 _5713_/B sky130_fd_sc_hd__a21o_2
XFILLER_108_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7406_ _7413_/A _7413_/B _6022_/X vssd1 vssd1 vccd1 vccd1 _7416_/B sky130_fd_sc_hd__o21bai_4
X_4618_ _7281_/A _5040_/A _7281_/B _5020_/A vssd1 vssd1 vccd1 vccd1 _4619_/C sky130_fd_sc_hd__a22o_2
X_5598_ _5650_/A _5599_/B vssd1 vssd1 vccd1 vccd1 _5598_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_104_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7337_ _7354_/A _7338_/B vssd1 vssd1 vccd1 vccd1 _7351_/A sky130_fd_sc_hd__nand2b_4
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4549_ _5090_/A _4654_/A _7001_/A _4585_/B vssd1 vssd1 vccd1 vccd1 _4552_/A sky130_fd_sc_hd__or4b_4
XFILLER_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7268_ _7268_/A _7268_/B vssd1 vssd1 vccd1 vccd1 _7274_/A sky130_fd_sc_hd__xnor2_4
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6219_ _6219_/A _6219_/B _6219_/C vssd1 vssd1 vccd1 vccd1 _6219_/X sky130_fd_sc_hd__and3_1
XFILLER_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7199_ _7199_/A _7199_/B vssd1 vssd1 vccd1 vccd1 _7474_/A sky130_fd_sc_hd__nand2_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6570_ _6570_/A _6570_/B vssd1 vssd1 vccd1 vccd1 _6570_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5521_ _5521_/A _5521_/B vssd1 vssd1 vccd1 vccd1 _5562_/A sky130_fd_sc_hd__xor2_4
XFILLER_117_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5452_ _5453_/A _5453_/B vssd1 vssd1 vccd1 vccd1 _5477_/A sky130_fd_sc_hd__nand2_1
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4403_ _7245_/A _4407_/A _4430_/C _4436_/A vssd1 vssd1 vccd1 vccd1 _4403_/X sky130_fd_sc_hd__o211a_1
X_5383_ _5542_/B _6970_/A _5375_/A _5375_/B vssd1 vssd1 vccd1 vccd1 _5391_/A sky130_fd_sc_hd__a22o_4
X_4334_ _4334_/A _4334_/B vssd1 vssd1 vccd1 vccd1 _4334_/Y sky130_fd_sc_hd__nand2_1
X_7122_ _7122_/A _7216_/A vssd1 vssd1 vccd1 vccd1 _7122_/X sky130_fd_sc_hd__or2_1
XFILLER_115_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout217 _7562_/X vssd1 vssd1 vccd1 vccd1 _7857_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_99_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout206 _7974_/X vssd1 vssd1 vccd1 vccd1 _7986_/S sky130_fd_sc_hd__buf_6
Xfanout228 _4168_/B1 vssd1 vssd1 vccd1 vccd1 _4211_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7053_ _7053_/A _7053_/B vssd1 vssd1 vccd1 vccd1 _7054_/B sky130_fd_sc_hd__nand2_1
Xfanout239 _7952_/B1 vssd1 vssd1 vccd1 vccd1 _7991_/D sky130_fd_sc_hd__buf_4
X_6004_ _7398_/A _6003_/Y _6084_/A vssd1 vssd1 vccd1 vccd1 _6078_/A sky130_fd_sc_hd__o21a_4
XFILLER_86_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4265_ _4200_/B _4260_/C _4264_/X _4548_/B vssd1 vssd1 vccd1 vccd1 _4266_/B sky130_fd_sc_hd__a211o_4
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4196_ _4211_/B _4196_/B vssd1 vssd1 vccd1 vccd1 _4204_/B sky130_fd_sc_hd__nand2_4
XFILLER_55_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7955_ _8043_/Q _8044_/Q _7955_/S vssd1 vssd1 vccd1 vccd1 _8044_/D sky130_fd_sc_hd__mux2_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7886_ _7886_/A _7908_/A _7886_/C vssd1 vssd1 vccd1 vccd1 _7910_/C sky130_fd_sc_hd__or3_1
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6906_ _7057_/A _7150_/B _6900_/X vssd1 vssd1 vccd1 vccd1 _6906_/X sky130_fd_sc_hd__o21a_1
X_6837_ _6873_/A _6878_/B _6784_/C vssd1 vssd1 vccd1 vccd1 _6838_/B sky130_fd_sc_hd__a21oi_2
XFILLER_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6768_ _7580_/C _6768_/B vssd1 vssd1 vccd1 vccd1 _7579_/B sky130_fd_sc_hd__xor2_1
XFILLER_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6699_ _6693_/X _6698_/X _6751_/S vssd1 vssd1 vccd1 vccd1 _6699_/X sky130_fd_sc_hd__mux2_1
X_5719_ _5720_/A _5720_/B vssd1 vssd1 vccd1 vccd1 _5719_/X sky130_fd_sc_hd__and2b_1
XFILLER_104_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4050_ _8059_/Q _4050_/B vssd1 vssd1 vccd1 vccd1 _4050_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_64_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7740_ _7721_/B _7720_/Y _7935_/A vssd1 vssd1 vccd1 vccd1 _7741_/B sky130_fd_sc_hd__o21a_1
X_4952_ _4923_/X _4952_/B vssd1 vssd1 vccd1 vccd1 _4960_/B sky130_fd_sc_hd__and2b_2
XFILLER_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7671_ _7671_/A _7731_/A vssd1 vssd1 vccd1 vccd1 _7760_/A sky130_fd_sc_hd__xor2_4
XFILLER_60_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4883_ _4998_/A _4947_/C _4876_/A _4877_/X vssd1 vssd1 vccd1 vccd1 _4911_/A sky130_fd_sc_hd__a31o_2
X_6622_ _6622_/A vssd1 vssd1 vccd1 vccd1 _6623_/B sky130_fd_sc_hd__inv_2
XFILLER_60_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6553_ _6581_/B vssd1 vssd1 vccd1 vccd1 _6554_/B sky130_fd_sc_hd__inv_2
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6484_ _6439_/X _6483_/Y _6484_/S vssd1 vssd1 vccd1 vccd1 _6485_/B sky130_fd_sc_hd__mux2_1
X_5504_ _5504_/A _5504_/B vssd1 vssd1 vccd1 vccd1 _5526_/A sky130_fd_sc_hd__xnor2_4
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5435_ _5407_/A _5407_/B _5408_/A _5408_/B vssd1 vssd1 vccd1 vccd1 _5440_/A sky130_fd_sc_hd__a22o_4
X_5366_ _5889_/A vssd1 vssd1 vccd1 vccd1 _5369_/B sky130_fd_sc_hd__inv_2
X_4317_ _4317_/A _4317_/B vssd1 vssd1 vccd1 vccd1 _4319_/B sky130_fd_sc_hd__and2_1
XFILLER_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7105_ _7104_/B _7105_/B vssd1 vssd1 vccd1 vccd1 _7106_/B sky130_fd_sc_hd__nand2b_1
X_5297_ _5298_/A _5298_/B vssd1 vssd1 vccd1 vccd1 _5347_/A sky130_fd_sc_hd__nand2_2
XFILLER_101_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4248_ _4212_/Y _5989_/B _4246_/X _4315_/B _4322_/A vssd1 vssd1 vccd1 vccd1 _4248_/X
+ sky130_fd_sc_hd__o2111a_2
X_7036_ _7036_/A _7036_/B _7036_/C vssd1 vssd1 vccd1 vccd1 _7037_/B sky130_fd_sc_hd__nand3_1
X_4179_ _8075_/Q _4179_/B vssd1 vssd1 vccd1 vccd1 _4228_/B sky130_fd_sc_hd__xnor2_4
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7938_ _7766_/B _7746_/Y _7913_/X _7766_/Y vssd1 vssd1 vccd1 vccd1 _7940_/A sky130_fd_sc_hd__a31o_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7869_ _7869_/A _7869_/B vssd1 vssd1 vccd1 vccd1 _7869_/X sky130_fd_sc_hd__xor2_1
XFILLER_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_3__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _8063_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5220_ _5220_/A _5220_/B vssd1 vssd1 vccd1 vccd1 _5239_/B sky130_fd_sc_hd__xor2_4
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5151_ _5264_/A _6783_/A _5151_/C vssd1 vssd1 vccd1 vccd1 _5154_/A sky130_fd_sc_hd__and3b_2
XFILLER_110_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4102_ _4102_/A _4102_/B vssd1 vssd1 vccd1 vccd1 _4107_/A sky130_fd_sc_hd__or2_1
X_5082_ _5080_/X _5081_/X _5268_/A vssd1 vssd1 vccd1 vccd1 _5082_/X sky130_fd_sc_hd__a21o_2
XFILLER_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4033_ _8022_/Q _8023_/Q _7955_/S vssd1 vssd1 vccd1 vccd1 _8023_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7723_ _7720_/Y _7721_/X _7722_/Y vssd1 vssd1 vccd1 vccd1 _7723_/X sky130_fd_sc_hd__a21o_1
X_5984_ _5986_/S _5984_/B vssd1 vssd1 vccd1 vccd1 _5984_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4935_ _5033_/B _4935_/B vssd1 vssd1 vccd1 vccd1 _4971_/A sky130_fd_sc_hd__xnor2_4
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7654_ _7654_/A _7654_/B vssd1 vssd1 vccd1 vccd1 _7654_/Y sky130_fd_sc_hd__nor2_1
X_4866_ _4866_/A _4866_/B vssd1 vssd1 vccd1 vccd1 _4867_/B sky130_fd_sc_hd__or2_1
X_6605_ _6605_/A _6605_/B _6612_/A vssd1 vssd1 vccd1 vccd1 _6606_/B sky130_fd_sc_hd__nor3_1
X_7585_ _7619_/A _7619_/B vssd1 vssd1 vccd1 vccd1 _7620_/A sky130_fd_sc_hd__nand2_2
X_4797_ _4795_/A _4795_/B _4795_/C vssd1 vssd1 vccd1 vccd1 _4923_/C sky130_fd_sc_hd__a21oi_2
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6536_ _6536_/A _6536_/B vssd1 vssd1 vccd1 vccd1 _6538_/B sky130_fd_sc_hd__xnor2_4
XFILLER_118_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6467_ _6378_/Y _6466_/Y _6373_/X vssd1 vssd1 vccd1 vccd1 _6467_/Y sky130_fd_sc_hd__o21ai_4
X_6398_ _6398_/A vssd1 vssd1 vccd1 vccd1 _6399_/B sky130_fd_sc_hd__inv_2
X_5418_ _5419_/A _5419_/B vssd1 vssd1 vccd1 vccd1 _5450_/A sky130_fd_sc_hd__nor2_4
X_5349_ _5294_/A _5294_/B _5296_/A _5296_/B vssd1 vssd1 vccd1 vccd1 _5356_/A sky130_fd_sc_hd__a2bb2oi_4
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8068_ _8075_/CLK _8068_/D vssd1 vssd1 vccd1 vccd1 _8068_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_75_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7019_ _7036_/B _7036_/C _7036_/A vssd1 vssd1 vccd1 vccd1 _7039_/A sky130_fd_sc_hd__a21o_1
XFILLER_28_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4720_/A _4720_/B _4720_/C vssd1 vssd1 vccd1 vccd1 _4720_/X sky130_fd_sc_hd__and3_1
XFILLER_42_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4651_ _4650_/B _4650_/C _4650_/A vssd1 vssd1 vccd1 vccd1 _4652_/C sky130_fd_sc_hd__a21o_1
XFILLER_30_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7370_ _7370_/A _7370_/B vssd1 vssd1 vccd1 vccd1 _7371_/C sky130_fd_sc_hd__xnor2_1
X_4582_ _4577_/A _4578_/X _4569_/X _4571_/Y vssd1 vssd1 vccd1 vccd1 _4583_/B sky130_fd_sc_hd__a211oi_4
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6321_ _6374_/A vssd1 vssd1 vccd1 vccd1 _6386_/A sky130_fd_sc_hd__inv_2
X_6252_ _6210_/X _6249_/X _6250_/Y _6251_/X vssd1 vssd1 vccd1 vccd1 _6258_/B sky130_fd_sc_hd__o31a_1
XFILLER_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6183_ _6182_/X _6012_/A _6199_/S vssd1 vssd1 vccd1 vccd1 _6183_/X sky130_fd_sc_hd__mux2_1
X_5203_ _5241_/A _5241_/B vssd1 vssd1 vccd1 vccd1 _5215_/B sky130_fd_sc_hd__nand2_4
XFILLER_111_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5134_ _4084_/B _5134_/A2 _4122_/X _4303_/B vssd1 vssd1 vccd1 vccd1 _5977_/C sky130_fd_sc_hd__a211o_4
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5065_ _4124_/X _4125_/X _5977_/B vssd1 vssd1 vccd1 vccd1 _5065_/Y sky130_fd_sc_hd__a21oi_4
X_4016_ _8018_/Q _8010_/Q _4016_/S vssd1 vssd1 vccd1 vccd1 _8010_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5967_ _7025_/A _7334_/A _7284_/A _7334_/B vssd1 vssd1 vccd1 vccd1 _5969_/C sky130_fd_sc_hd__and4_2
X_7706_ _7706_/A _7706_/B vssd1 vssd1 vccd1 vccd1 _7706_/X sky130_fd_sc_hd__or2_1
X_4918_ _4989_/A _5013_/C vssd1 vssd1 vccd1 vccd1 _4957_/A sky130_fd_sc_hd__or2_4
XFILLER_40_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7637_ _8030_/Q _7857_/B _7636_/X vssd1 vssd1 vccd1 vccd1 _7638_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5898_ _5897_/B _5912_/A _5897_/A vssd1 vssd1 vccd1 vccd1 _5933_/B sky130_fd_sc_hd__a21o_1
X_4849_ _4847_/X _4848_/Y _4773_/A vssd1 vssd1 vccd1 vccd1 _4868_/D sky130_fd_sc_hd__a21oi_4
XFILLER_32_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7568_ _7611_/D _7568_/B vssd1 vssd1 vccd1 vccd1 _7569_/C sky130_fd_sc_hd__or2_2
XFILLER_106_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6519_ _6465_/X _6507_/Y _7607_/A vssd1 vssd1 vccd1 vccd1 _6520_/B sky130_fd_sc_hd__mux2_2
X_7499_ _7456_/X _7450_/X _7624_/S vssd1 vssd1 vccd1 vccd1 _7500_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6870_ _6870_/A _6870_/B vssd1 vssd1 vccd1 vccd1 _6877_/A sky130_fd_sc_hd__nand2_1
X_5821_ _5822_/B _5821_/B vssd1 vssd1 vccd1 vccd1 _5825_/A sky130_fd_sc_hd__or2_1
XFILLER_34_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5752_ _5755_/A _5855_/A _5716_/Y vssd1 vssd1 vccd1 vccd1 _5759_/B sky130_fd_sc_hd__o21bai_4
X_4703_ _4709_/B _4703_/B vssd1 vssd1 vccd1 vccd1 _4836_/A sky130_fd_sc_hd__or2_4
X_5683_ _5683_/A _5683_/B _5684_/B vssd1 vssd1 vccd1 vccd1 _5694_/A sky130_fd_sc_hd__or3_4
XFILLER_8_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7422_ _7766_/A _7422_/B vssd1 vssd1 vccd1 vccd1 _7423_/B sky130_fd_sc_hd__or2_4
X_4634_ _4634_/A _4641_/B _4634_/C vssd1 vssd1 vccd1 vccd1 _4636_/B sky130_fd_sc_hd__nand3_4
X_4565_ _4453_/B _4453_/C _4453_/A vssd1 vssd1 vccd1 vccd1 _4566_/C sky130_fd_sc_hd__a21o_2
X_7353_ _7281_/B _7281_/D _7085_/B _7281_/A vssd1 vssd1 vccd1 vccd1 _7354_/B sky130_fd_sc_hd__a22o_1
XFILLER_116_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6304_ _6304_/A _6564_/A vssd1 vssd1 vccd1 vccd1 _6305_/B sky130_fd_sc_hd__or2_4
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7284_ _7284_/A _7358_/B vssd1 vssd1 vccd1 vccd1 _7366_/C sky130_fd_sc_hd__or2_2
X_4496_ _7247_/A _4496_/B vssd1 vssd1 vccd1 vccd1 _4497_/C sky130_fd_sc_hd__xnor2_4
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6235_ _5923_/A _7085_/B _5858_/B _5880_/Y vssd1 vssd1 vccd1 vccd1 _6238_/B sky130_fd_sc_hd__o22a_1
XFILLER_103_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6166_ _6142_/X _6165_/Y _6166_/S vssd1 vssd1 vccd1 vccd1 _6166_/X sky130_fd_sc_hd__mux2_2
XFILLER_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6097_ _6088_/Y _6092_/B _6096_/Y _7639_/A vssd1 vssd1 vccd1 vccd1 _6099_/A sky130_fd_sc_hd__o211ai_4
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _5062_/A _5062_/B _5100_/A _4787_/A vssd1 vssd1 vccd1 vccd1 _5121_/B sky130_fd_sc_hd__a211o_2
XFILLER_57_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5048_ _5029_/X _5714_/A _5299_/A vssd1 vssd1 vccd1 vccd1 _5703_/B sky130_fd_sc_hd__a21o_2
XFILLER_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6999_ _6999_/A _7269_/B vssd1 vssd1 vccd1 vccd1 _7056_/A sky130_fd_sc_hd__nand2_4
XFILLER_40_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4350_ _7136_/A _4349_/Y _4494_/A vssd1 vssd1 vccd1 vccd1 _4350_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4281_ _4178_/X _4260_/C _4235_/X _4548_/B vssd1 vssd1 vccd1 vccd1 _4281_/X sky130_fd_sc_hd__a211o_1
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6020_ _6020_/A vssd1 vssd1 vccd1 vccd1 _6020_/Y sky130_fd_sc_hd__inv_2
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7971_ _7970_/X _7971_/B _7971_/C vssd1 vssd1 vccd1 vccd1 _8049_/D sky130_fd_sc_hd__and3b_1
XFILLER_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6922_ _7030_/A _7235_/B vssd1 vssd1 vccd1 vccd1 _6964_/A sky130_fd_sc_hd__nor2_2
X_6853_ _6863_/A _6863_/B vssd1 vssd1 vccd1 vccd1 _6857_/B sky130_fd_sc_hd__nand2b_1
XFILLER_35_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout17 _6635_/Y vssd1 vssd1 vccd1 vccd1 _7718_/S sky130_fd_sc_hd__buf_2
Xfanout28 _7433_/X vssd1 vssd1 vccd1 vccd1 _7535_/A sky130_fd_sc_hd__buf_6
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5804_ _5804_/A _5804_/B vssd1 vssd1 vccd1 vccd1 _5806_/B sky130_fd_sc_hd__xnor2_4
XFILLER_35_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout39 _7394_/X vssd1 vssd1 vccd1 vccd1 _7479_/S sky130_fd_sc_hd__clkbuf_4
X_6784_ _6873_/A _6878_/B _6784_/C vssd1 vssd1 vccd1 vccd1 _6838_/A sky130_fd_sc_hd__and3_2
X_5735_ _5736_/B _5736_/C vssd1 vssd1 vccd1 vccd1 _5771_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5666_ _5666_/A _5666_/B vssd1 vssd1 vccd1 vccd1 _5666_/Y sky130_fd_sc_hd__nor2_1
X_7405_ _5997_/Y _7398_/B _6000_/B vssd1 vssd1 vccd1 vccd1 _7413_/B sky130_fd_sc_hd__a21oi_4
X_4617_ _7214_/A _5013_/A vssd1 vssd1 vccd1 vccd1 _4619_/B sky130_fd_sc_hd__nor2_2
XFILLER_116_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5597_ _5597_/A _5597_/B vssd1 vssd1 vccd1 vccd1 _5599_/B sky130_fd_sc_hd__xor2_4
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4548_ _4548_/A _4548_/B _4548_/C _4547_/D vssd1 vssd1 vccd1 vccd1 _4548_/X sky130_fd_sc_hd__or4b_4
X_7336_ _7336_/A _7336_/B vssd1 vssd1 vccd1 vccd1 _7338_/B sky130_fd_sc_hd__and2_4
X_7267_ _7275_/A _7275_/B _7265_/X vssd1 vssd1 vccd1 vccd1 _7268_/B sky130_fd_sc_hd__o21a_2
X_4479_ _4474_/X _4478_/Y _7085_/A vssd1 vssd1 vccd1 vccd1 _4570_/A sky130_fd_sc_hd__o21a_4
X_6218_ _6203_/Y _6217_/Y _6226_/S vssd1 vssd1 vccd1 vccd1 _6255_/C sky130_fd_sc_hd__mux2_2
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7198_ _7197_/B _7198_/B vssd1 vssd1 vccd1 vccd1 _7199_/B sky130_fd_sc_hd__nand2b_1
X_6149_ _5204_/X _6139_/B _6127_/A _6148_/Y _6146_/X vssd1 vssd1 vccd1 vccd1 _6149_/X
+ sky130_fd_sc_hd__o221a_2
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5520_ _5521_/A _5521_/B vssd1 vssd1 vccd1 vccd1 _5520_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5451_ _5451_/A _5451_/B vssd1 vssd1 vccd1 vccd1 _5453_/B sky130_fd_sc_hd__xor2_2
X_4402_ _7245_/A _4407_/A _4430_/C vssd1 vssd1 vccd1 vccd1 _4402_/X sky130_fd_sc_hd__o21a_1
X_5382_ _5336_/A _5334_/Y _5333_/Y vssd1 vssd1 vccd1 vccd1 _5394_/A sky130_fd_sc_hd__o21a_4
XFILLER_113_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7121_ _5087_/B _4296_/Y _7284_/A _5145_/X _5322_/A vssd1 vssd1 vccd1 vccd1 _7216_/A
+ sky130_fd_sc_hd__a2111o_4
X_4333_ _4334_/A _4334_/B vssd1 vssd1 vccd1 vccd1 _7068_/A sky130_fd_sc_hd__and2_4
Xfanout218 _7562_/X vssd1 vssd1 vccd1 vccd1 _7944_/B sky130_fd_sc_hd__clkbuf_4
Xfanout207 _7974_/X vssd1 vssd1 vccd1 vccd1 _7990_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout229 _6770_/A vssd1 vssd1 vccd1 vccd1 _4168_/B1 sky130_fd_sc_hd__clkbuf_4
X_4264_ _4241_/B _4227_/X _4231_/X _6278_/B vssd1 vssd1 vccd1 vccd1 _4264_/X sky130_fd_sc_hd__o211a_1
X_7052_ _7052_/A _7052_/B vssd1 vssd1 vccd1 vccd1 _7102_/A sky130_fd_sc_hd__xor2_4
X_6003_ _4258_/X _6009_/A _6001_/X vssd1 vssd1 vccd1 vccd1 _6003_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_67_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4195_ _4216_/B _4200_/B vssd1 vssd1 vccd1 vccd1 _4195_/X sky130_fd_sc_hd__or2_1
XFILLER_39_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7954_ _7974_/A _7954_/B _7954_/C vssd1 vssd1 vccd1 vccd1 _8043_/D sky130_fd_sc_hd__and3b_1
XFILLER_82_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6905_ _6913_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6942_/A sky130_fd_sc_hd__nand2_2
X_7885_ _7909_/B _7909_/C vssd1 vssd1 vccd1 vccd1 _7888_/A sky130_fd_sc_hd__nor2_1
X_6836_ _6836_/A _6836_/B vssd1 vssd1 vccd1 vccd1 _6849_/A sky130_fd_sc_hd__xnor2_1
XFILLER_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6767_ _6770_/A _6188_/A _6767_/S vssd1 vssd1 vccd1 vccd1 _7935_/A sky130_fd_sc_hd__mux2_8
XFILLER_50_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5718_ _5666_/A _5714_/X _5759_/A vssd1 vssd1 vccd1 vccd1 _5720_/B sky130_fd_sc_hd__a21bo_2
X_6698_ _6692_/X _6697_/X _6713_/S vssd1 vssd1 vccd1 vccd1 _6698_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5649_ _5367_/A _5853_/B _5648_/A vssd1 vssd1 vccd1 vccd1 _5650_/B sky130_fd_sc_hd__o21ai_1
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7319_ _7319_/A _7319_/B vssd1 vssd1 vccd1 vccd1 _7326_/A sky130_fd_sc_hd__nand2_2
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4951_ _4923_/B _4923_/C _4947_/C _5040_/A vssd1 vssd1 vccd1 vccd1 _4952_/B sky130_fd_sc_hd__a22o_1
X_7670_ _7702_/A _7731_/A _7757_/D vssd1 vssd1 vccd1 vccd1 _7703_/A sky130_fd_sc_hd__or3b_4
X_4882_ _4884_/A _4884_/B vssd1 vssd1 vccd1 vccd1 _4882_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6621_ _6621_/A _6621_/B vssd1 vssd1 vccd1 vccd1 _6622_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6552_ _6552_/A _6552_/B vssd1 vssd1 vccd1 vccd1 _6581_/B sky130_fd_sc_hd__nand2_2
X_6483_ _6483_/A _6483_/B vssd1 vssd1 vccd1 vccd1 _6483_/Y sky130_fd_sc_hd__nor2_1
X_5503_ _5503_/A _5503_/B vssd1 vssd1 vccd1 vccd1 _5549_/A sky130_fd_sc_hd__xnor2_4
XFILLER_106_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5434_ _5434_/A _5434_/B vssd1 vssd1 vccd1 vccd1 _5441_/A sky130_fd_sc_hd__nor2_4
XFILLER_114_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7104_ _7105_/B _7104_/B vssd1 vssd1 vccd1 vccd1 _7106_/A sky130_fd_sc_hd__nand2b_1
X_5365_ _5925_/A _5855_/B vssd1 vssd1 vccd1 vccd1 _5889_/A sky130_fd_sc_hd__or2_4
XFILLER_113_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4316_ _4216_/C _4259_/B _4261_/X _4548_/B vssd1 vssd1 vccd1 vccd1 _4317_/B sky130_fd_sc_hd__a211o_2
X_5296_ _5296_/A _5296_/B vssd1 vssd1 vccd1 vccd1 _5298_/B sky130_fd_sc_hd__xor2_4
XFILLER_113_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4247_ _4212_/Y _5989_/B _4246_/X vssd1 vssd1 vccd1 vccd1 _4547_/D sky130_fd_sc_hd__o21a_1
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7035_ _7035_/A _7035_/B vssd1 vssd1 vccd1 vccd1 _7053_/A sky130_fd_sc_hd__nand2_1
X_4178_ _8074_/Q _4178_/B vssd1 vssd1 vccd1 vccd1 _4178_/X sky130_fd_sc_hd__xor2_4
XFILLER_67_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7937_ _7773_/A _7920_/X _7935_/Y _7936_/Y _6774_/X vssd1 vssd1 vccd1 vccd1 _7937_/X
+ sky130_fd_sc_hd__a311o_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7868_ _7793_/Y _7823_/Y _7844_/A _7649_/A vssd1 vssd1 vccd1 vccd1 _7869_/B sky130_fd_sc_hd__a31o_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6819_ _6819_/A _6819_/B vssd1 vssd1 vccd1 vccd1 _6820_/B sky130_fd_sc_hd__or2_4
X_7799_ _7766_/Y _7798_/B _7798_/A vssd1 vssd1 vccd1 vccd1 _7800_/B sky130_fd_sc_hd__o21ai_1
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5150_ _5207_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _5275_/A sky130_fd_sc_hd__or2_2
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4101_ _6326_/A _6278_/A vssd1 vssd1 vccd1 vccd1 _4102_/B sky130_fd_sc_hd__xnor2_1
X_5081_ _4094_/B _5134_/A2 _4293_/X _5135_/C1 vssd1 vssd1 vccd1 vccd1 _5081_/X sky130_fd_sc_hd__a211o_2
XFILLER_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4032_ _8021_/Q _8022_/Q _7955_/S vssd1 vssd1 vccd1 vccd1 _8022_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5983_ _5268_/A _5080_/X _5081_/X _5981_/X _5982_/X vssd1 vssd1 vccd1 vccd1 _5984_/B
+ sky130_fd_sc_hd__a32oi_4
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7722_ _7720_/Y _7721_/X _7923_/A vssd1 vssd1 vccd1 vccd1 _7722_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4934_ _5033_/B _4935_/B vssd1 vssd1 vccd1 vccd1 _4934_/X sky130_fd_sc_hd__and2b_1
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7653_ _7677_/A _7677_/B vssd1 vssd1 vccd1 vccd1 _7654_/B sky130_fd_sc_hd__xnor2_2
X_4865_ _4865_/A _4865_/B vssd1 vssd1 vccd1 vccd1 _4887_/A sky130_fd_sc_hd__xnor2_4
X_7584_ _6732_/A _7583_/X _7894_/A vssd1 vssd1 vccd1 vccd1 _7619_/B sky130_fd_sc_hd__mux2_2
X_6604_ _6302_/A _6302_/B _6602_/A _6603_/Y vssd1 vssd1 vccd1 vccd1 _7773_/A sky130_fd_sc_hd__o22ai_4
X_4796_ _4795_/A _4795_/B _4795_/C vssd1 vssd1 vccd1 vccd1 _4798_/A sky130_fd_sc_hd__a21o_1
XFILLER_20_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6535_ _6460_/Y _6503_/Y _6544_/S vssd1 vssd1 vccd1 vccd1 _6536_/B sky130_fd_sc_hd__mux2_4
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6466_ _6520_/A _6465_/X _6386_/X vssd1 vssd1 vccd1 vccd1 _6466_/Y sky130_fd_sc_hd__a21oi_4
X_6397_ _6397_/A _6397_/B vssd1 vssd1 vccd1 vccd1 _6398_/A sky130_fd_sc_hd__and2_1
X_5417_ _5446_/B _6916_/C vssd1 vssd1 vccd1 vccd1 _5419_/B sky130_fd_sc_hd__xor2_4
X_5348_ _5325_/B _5353_/A _5332_/A _5332_/B vssd1 vssd1 vccd1 vccd1 _5357_/A sky130_fd_sc_hd__a2bb2o_4
X_8067_ _8075_/CLK _8067_/D vssd1 vssd1 vccd1 vccd1 _8067_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_101_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5279_ _5267_/A _5267_/B _5276_/A _5466_/A vssd1 vssd1 vccd1 vccd1 _5492_/A sky130_fd_sc_hd__a2bb2o_4
X_7018_ _7055_/A _7055_/B vssd1 vssd1 vccd1 vccd1 _7036_/C sky130_fd_sc_hd__or2_1
XFILLER_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _4650_/A _4650_/B _4650_/C vssd1 vssd1 vccd1 vccd1 _4652_/B sky130_fd_sc_hd__nand3_2
XFILLER_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6320_ _6320_/A _6320_/B vssd1 vssd1 vccd1 vccd1 _6374_/A sky130_fd_sc_hd__xnor2_4
X_4581_ _4581_/A _4581_/B _4583_/A vssd1 vssd1 vccd1 vccd1 _4735_/B sky130_fd_sc_hd__or3_1
XFILLER_116_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6251_ _6112_/C _6248_/X _6245_/C _6166_/S vssd1 vssd1 vccd1 vccd1 _6251_/X sky130_fd_sc_hd__a211o_1
XFILLER_103_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6182_ _5745_/A _6139_/B _6146_/A _6172_/X _6181_/Y vssd1 vssd1 vccd1 vccd1 _6182_/X
+ sky130_fd_sc_hd__o221a_1
X_5202_ _5202_/A _5202_/B vssd1 vssd1 vccd1 vccd1 _5241_/B sky130_fd_sc_hd__xor2_4
X_5133_ _5133_/A _5133_/B vssd1 vssd1 vccd1 vccd1 _5133_/Y sky130_fd_sc_hd__nand2_2
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5064_ _6806_/A _5582_/A vssd1 vssd1 vccd1 vccd1 _5174_/A sky130_fd_sc_hd__or2_4
X_4015_ _8017_/Q _8009_/Q _4016_/S vssd1 vssd1 vccd1 vccd1 _8009_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5966_ _5970_/A _5970_/B vssd1 vssd1 vccd1 vccd1 _6242_/S sky130_fd_sc_hd__and2_4
X_7705_ _6544_/S _7697_/Y _7760_/B _6269_/X vssd1 vssd1 vccd1 vccd1 _7706_/B sky130_fd_sc_hd__a31o_1
XFILLER_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4917_ _4988_/A _5013_/C _4947_/C _5019_/A vssd1 vssd1 vccd1 vccd1 _4921_/A sky130_fd_sc_hd__a2bb2o_2
X_5897_ _5897_/A _5897_/B _5912_/A vssd1 vssd1 vccd1 vccd1 _5897_/Y sky130_fd_sc_hd__nand3_1
X_7636_ _7614_/Y _7633_/X _7634_/X _7635_/X vssd1 vssd1 vccd1 vccd1 _7636_/X sky130_fd_sc_hd__o31a_2
X_4848_ _4848_/A _4848_/B vssd1 vssd1 vccd1 vccd1 _4848_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7567_ _7611_/D _7611_/C vssd1 vssd1 vccd1 vccd1 _7576_/A sky130_fd_sc_hd__nand2_4
X_4779_ _4779_/A _4779_/B vssd1 vssd1 vccd1 vccd1 _4790_/B sky130_fd_sc_hd__nor2_1
X_6518_ _6515_/Y _6709_/A vssd1 vssd1 vccd1 vccd1 _6525_/A sky130_fd_sc_hd__nand2b_2
XFILLER_106_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7498_ _7465_/X _7535_/B _7538_/S vssd1 vssd1 vccd1 vccd1 _7544_/C sky130_fd_sc_hd__mux2_2
X_6449_ _6483_/A _6483_/B vssd1 vssd1 vccd1 vccd1 _6449_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5820_ _5880_/A _7344_/B vssd1 vssd1 vccd1 vccd1 _5859_/A sky130_fd_sc_hd__or2_1
XFILLER_34_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5751_ _5751_/A _5751_/B vssd1 vssd1 vccd1 vccd1 _5786_/A sky130_fd_sc_hd__xnor2_4
X_4702_ _4709_/B _4703_/B vssd1 vssd1 vccd1 vccd1 _4702_/Y sky130_fd_sc_hd__nor2_1
X_7421_ _7421_/A _7421_/B _7421_/C vssd1 vssd1 vccd1 vccd1 _7422_/B sky130_fd_sc_hd__nor3_2
X_5682_ _5672_/A _5925_/A _5677_/B _5675_/X vssd1 vssd1 vccd1 vccd1 _5684_/B sky130_fd_sc_hd__o31a_4
X_4633_ _4641_/A _4632_/C _4632_/A vssd1 vssd1 vccd1 vccd1 _4634_/C sky130_fd_sc_hd__a21o_1
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7352_ _7352_/A _7352_/B vssd1 vssd1 vccd1 vccd1 _7367_/A sky130_fd_sc_hd__xnor2_2
X_4564_ _4563_/A _4563_/B _4563_/C _4555_/X vssd1 vssd1 vccd1 vccd1 _4566_/B sky130_fd_sc_hd__a31o_2
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6303_ _6308_/A _6303_/B vssd1 vssd1 vccd1 vccd1 _6601_/A sky130_fd_sc_hd__xnor2_2
X_7283_ _7283_/A _7304_/A vssd1 vssd1 vccd1 vccd1 _7286_/A sky130_fd_sc_hd__xor2_4
XFILLER_116_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4495_ _4495_/A _4495_/B vssd1 vssd1 vccd1 vccd1 _4496_/B sky130_fd_sc_hd__xor2_4
X_6234_ _5928_/A _6233_/X _5928_/X vssd1 vssd1 vccd1 vccd1 _6238_/A sky130_fd_sc_hd__o21ba_1
X_6165_ _6193_/A _6153_/Y _6164_/Y vssd1 vssd1 vccd1 vccd1 _6165_/Y sky130_fd_sc_hd__a21oi_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6096_ _6096_/A _6096_/B vssd1 vssd1 vccd1 vccd1 _6096_/Y sky130_fd_sc_hd__xnor2_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _4786_/A _5097_/Y _5098_/A vssd1 vssd1 vccd1 vccd1 _5121_/A sky130_fd_sc_hd__a21o_1
XFILLER_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5047_ _5047_/A _5047_/B _5047_/C vssd1 vssd1 vccd1 vccd1 _5714_/A sky130_fd_sc_hd__or3_4
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6998_ _6998_/A _6998_/B vssd1 vssd1 vccd1 vccd1 _7016_/A sky130_fd_sc_hd__and2_1
XFILLER_41_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5949_ _5499_/A _5496_/Y _5499_/B vssd1 vssd1 vccd1 vccd1 _5949_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7619_ _7619_/A _7619_/B _7620_/B vssd1 vssd1 vccd1 vccd1 _7677_/A sky130_fd_sc_hd__and3_4
XFILLER_119_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4280_ _6315_/A vssd1 vssd1 vccd1 vccd1 _6310_/A sky130_fd_sc_hd__clkinv_4
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7970_ _8049_/Q _8048_/Q _7970_/C vssd1 vssd1 vccd1 vccd1 _7970_/X sky130_fd_sc_hd__and3_1
XFILLER_94_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6921_ _6923_/B _6923_/A vssd1 vssd1 vccd1 vccd1 _6921_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6852_ _7123_/A _6951_/D _6947_/C vssd1 vssd1 vccd1 vccd1 _6863_/B sky130_fd_sc_hd__and3_2
Xfanout18 _7583_/S vssd1 vssd1 vccd1 vccd1 _6749_/S sky130_fd_sc_hd__clkbuf_8
Xfanout29 _7433_/X vssd1 vssd1 vccd1 vccd1 _7657_/B sky130_fd_sc_hd__buf_4
XFILLER_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5803_ _5795_/A _5826_/A _5837_/A vssd1 vssd1 vccd1 vccd1 _5806_/A sky130_fd_sc_hd__o21ai_4
X_6783_ _6783_/A _6783_/B vssd1 vssd1 vccd1 vccd1 _6784_/C sky130_fd_sc_hd__xnor2_2
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5734_ _5800_/A _5853_/B vssd1 vssd1 vccd1 vccd1 _5736_/C sky130_fd_sc_hd__nor2_1
X_5665_ _5755_/A _7344_/B vssd1 vssd1 vccd1 vccd1 _5713_/A sky130_fd_sc_hd__or2_4
X_7404_ _7421_/A vssd1 vssd1 vccd1 vccd1 _7419_/A sky130_fd_sc_hd__inv_2
X_4616_ _5014_/A _7001_/A _4616_/C vssd1 vssd1 vccd1 vccd1 _4620_/A sky130_fd_sc_hd__or3_4
X_5596_ _5596_/A _5596_/B vssd1 vssd1 vccd1 vccd1 _5597_/B sky130_fd_sc_hd__xnor2_4
X_7335_ _7311_/A _7371_/B _7311_/C vssd1 vssd1 vccd1 vccd1 _7336_/B sky130_fd_sc_hd__o21ai_1
X_4547_ _6034_/A _6017_/A _4547_/C _4547_/D vssd1 vssd1 vccd1 vccd1 _7281_/B sky130_fd_sc_hd__and4_4
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4478_ _4424_/A _4476_/X _4477_/X vssd1 vssd1 vccd1 vccd1 _4478_/Y sky130_fd_sc_hd__a21oi_1
X_7266_ _7266_/A _7266_/B vssd1 vssd1 vccd1 vccd1 _7275_/B sky130_fd_sc_hd__xnor2_2
XFILLER_104_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6217_ _6193_/A _6195_/X _6215_/X vssd1 vssd1 vccd1 vccd1 _6217_/Y sky130_fd_sc_hd__a21oi_1
X_7197_ _7198_/B _7197_/B vssd1 vssd1 vccd1 vccd1 _7199_/A sky130_fd_sc_hd__nand2b_4
XFILLER_85_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6148_ _6148_/A _6148_/B vssd1 vssd1 vccd1 vccd1 _6148_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_58_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _6078_/B _6078_/C _6078_/A vssd1 vssd1 vccd1 vccd1 _6081_/B sky130_fd_sc_hd__o21ai_4
XFILLER_73_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5450_ _5450_/A _5450_/B vssd1 vssd1 vccd1 vccd1 _5451_/B sky130_fd_sc_hd__xor2_4
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4401_ _4501_/A _4397_/Y _4399_/Y _4400_/X _4370_/Y vssd1 vssd1 vccd1 vccd1 _4401_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_99_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5381_ _5545_/A _5545_/B _5376_/Y vssd1 vssd1 vccd1 vccd1 _5395_/A sky130_fd_sc_hd__a21o_4
XFILLER_113_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4332_ _4341_/A1 _4287_/X _4288_/X _4356_/A vssd1 vssd1 vccd1 vccd1 _4334_/B sky130_fd_sc_hd__o31a_2
X_7120_ _7134_/B _7120_/B vssd1 vssd1 vccd1 vccd1 _7159_/A sky130_fd_sc_hd__and2_1
Xfanout219 _7886_/A vssd1 vssd1 vccd1 vccd1 _7929_/A sky130_fd_sc_hd__buf_4
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4263_ _4209_/X _4226_/X _4232_/Y _6278_/B vssd1 vssd1 vccd1 vccd1 _4263_/X sky130_fd_sc_hd__a211o_2
X_7051_ _7051_/A _7051_/B vssd1 vssd1 vccd1 vccd1 _7105_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout208 _5445_/A vssd1 vssd1 vccd1 vccd1 _4773_/A sky130_fd_sc_hd__buf_8
X_6002_ _4258_/X _6009_/A _6320_/A _6001_/X vssd1 vssd1 vccd1 vccd1 _6084_/A sky130_fd_sc_hd__a211o_4
X_4194_ _8071_/Q _4194_/B vssd1 vssd1 vccd1 vccd1 _4200_/B sky130_fd_sc_hd__xor2_4
XFILLER_67_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7953_ _8042_/Q _4020_/B _7563_/Y _8043_/Q vssd1 vssd1 vccd1 vccd1 _7954_/C sky130_fd_sc_hd__o22a_1
XFILLER_82_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6904_ _6903_/B _6903_/C _7067_/A _6903_/A vssd1 vssd1 vccd1 vccd1 _6905_/B sky130_fd_sc_hd__o22ai_2
X_7884_ _7883_/A _7883_/B _7883_/C vssd1 vssd1 vccd1 vccd1 _7909_/C sky130_fd_sc_hd__a21oi_1
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6835_ _6835_/A _6835_/B vssd1 vssd1 vccd1 vccd1 _6857_/A sky130_fd_sc_hd__or2_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6766_ _7949_/A _4005_/Y _6766_/S vssd1 vssd1 vccd1 vccd1 _7622_/A sky130_fd_sc_hd__mux2_2
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5717_ _5755_/A _5855_/A _5716_/Y vssd1 vssd1 vccd1 vccd1 _5759_/A sky130_fd_sc_hd__or3b_4
X_6697_ _6696_/X _6655_/Y _6697_/S vssd1 vssd1 vccd1 vccd1 _6697_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5648_ _5648_/A _5736_/A vssd1 vssd1 vccd1 vccd1 _5654_/A sky130_fd_sc_hd__or2_4
X_5579_ _5579_/A _5579_/B vssd1 vssd1 vccd1 vccd1 _5580_/B sky130_fd_sc_hd__and2_1
X_7318_ _7327_/A _7327_/B vssd1 vssd1 vccd1 vccd1 _7328_/A sky130_fd_sc_hd__nor2_4
XFILLER_116_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7249_ _7278_/A _7278_/B vssd1 vssd1 vccd1 vccd1 _7257_/B sky130_fd_sc_hd__and2_2
XFILLER_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4950_ _4986_/A _4986_/B _4947_/X vssd1 vssd1 vccd1 vccd1 _4960_/A sky130_fd_sc_hd__a21o_2
X_4881_ _4906_/A _4880_/B _4872_/Y vssd1 vssd1 vccd1 vccd1 _4884_/B sky130_fd_sc_hd__a21o_2
X_6620_ _6621_/A _6621_/B vssd1 vssd1 vccd1 vccd1 _6623_/A sky130_fd_sc_hd__nand2_1
X_6551_ _6550_/B _6550_/C _6550_/D _7929_/A vssd1 vssd1 vccd1 vccd1 _6552_/B sky130_fd_sc_hd__o22ai_2
X_5502_ _5502_/A _5502_/B vssd1 vssd1 vccd1 vccd1 _5947_/A sky130_fd_sc_hd__or2_1
XFILLER_118_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6482_ _6482_/A _6482_/B vssd1 vssd1 vccd1 vccd1 _6550_/C sky130_fd_sc_hd__and2_1
XFILLER_9_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5433_ _5432_/A _5432_/B _5432_/C vssd1 vssd1 vccd1 vccd1 _5434_/B sky130_fd_sc_hd__a21oi_2
X_5364_ _5364_/A _5364_/B vssd1 vssd1 vccd1 vccd1 _5364_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4315_ _4315_/A _4315_/B _5989_/B vssd1 vssd1 vccd1 vccd1 _4317_/A sky130_fd_sc_hd__or3_4
X_7103_ _7107_/A _7107_/B _7100_/X vssd1 vssd1 vccd1 vccd1 _7104_/B sky130_fd_sc_hd__o21ai_2
XFILLER_101_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5295_ _5715_/A _5672_/A vssd1 vssd1 vccd1 vccd1 _5296_/B sky130_fd_sc_hd__nor2_4
X_4246_ _4209_/X _4226_/X _4232_/Y _8067_/Q vssd1 vssd1 vccd1 vccd1 _4246_/X sky130_fd_sc_hd__a211o_1
X_7034_ _7034_/A _7034_/B vssd1 vssd1 vccd1 vccd1 _7035_/B sky130_fd_sc_hd__nand2_1
X_4177_ _8072_/Q _8071_/Q _8073_/Q _4175_/B _4211_/B vssd1 vssd1 vccd1 vccd1 _4178_/B
+ sky130_fd_sc_hd__o41a_4
XFILLER_55_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7936_ _7773_/A _7920_/X _7935_/Y vssd1 vssd1 vccd1 vccd1 _7936_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7867_ _7867_/A _7867_/B vssd1 vssd1 vccd1 vccd1 _7869_/A sky130_fd_sc_hd__or2_1
XFILLER_23_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6818_ _7025_/A _6805_/B _5164_/X vssd1 vssd1 vccd1 vccd1 _6819_/B sky130_fd_sc_hd__o21a_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7798_ _7798_/A _7798_/B vssd1 vssd1 vccd1 vccd1 _7817_/A sky130_fd_sc_hd__or2_2
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6749_ _6746_/X _6748_/X _6749_/S vssd1 vssd1 vccd1 vccd1 _7788_/B sky130_fd_sc_hd__mux2_1
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4100_ _8054_/Q _4100_/B vssd1 vssd1 vccd1 vccd1 _6278_/A sky130_fd_sc_hd__xor2_4
X_5080_ _4056_/S _5134_/A2 _4298_/X _4110_/Y vssd1 vssd1 vccd1 vccd1 _5080_/X sky130_fd_sc_hd__a211o_2
XFILLER_69_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4031_ _8020_/Q _8021_/Q _7955_/S vssd1 vssd1 vccd1 vccd1 _8021_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5982_ _4077_/B _4110_/Y _6030_/A vssd1 vssd1 vccd1 vccd1 _5982_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7721_ _7935_/A _7721_/B vssd1 vssd1 vccd1 vccd1 _7721_/X sky130_fd_sc_hd__and2_1
X_4933_ _4933_/A _4933_/B vssd1 vssd1 vccd1 vccd1 _4935_/B sky130_fd_sc_hd__xnor2_4
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7652_ _6732_/D _7651_/Y _7894_/A vssd1 vssd1 vccd1 vccd1 _7677_/B sky130_fd_sc_hd__mux2_4
X_4864_ _5058_/A vssd1 vssd1 vccd1 vccd1 _5189_/A sky130_fd_sc_hd__inv_2
XFILLER_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7583_ _6735_/X _7582_/Y _7583_/S vssd1 vssd1 vccd1 vccd1 _7583_/X sky130_fd_sc_hd__mux2_1
X_6603_ _6060_/Y _6302_/B _6303_/B _6308_/A vssd1 vssd1 vccd1 vccd1 _6603_/Y sky130_fd_sc_hd__o22ai_4
X_4795_ _4795_/A _4795_/B _4795_/C vssd1 vssd1 vccd1 vccd1 _4923_/B sky130_fd_sc_hd__or3_4
X_6534_ _6538_/A vssd1 vssd1 vccd1 vccd1 _6534_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6465_ _6393_/X _6397_/B _6464_/Y vssd1 vssd1 vccd1 vccd1 _6465_/X sky130_fd_sc_hd__a21bo_2
X_5416_ _5373_/B _6916_/C _5387_/Y _5389_/A vssd1 vssd1 vccd1 vccd1 _5419_/A sky130_fd_sc_hd__o2bb2a_4
X_6396_ _6397_/A _6397_/B vssd1 vssd1 vccd1 vccd1 _6399_/A sky130_fd_sc_hd__or2_2
XFILLER_114_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5347_ _5347_/A _5347_/B vssd1 vssd1 vccd1 vccd1 _5358_/A sky130_fd_sc_hd__xnor2_4
X_8066_ _8082_/CLK _8066_/D vssd1 vssd1 vccd1 vccd1 _8066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5278_ _5280_/A _5280_/B vssd1 vssd1 vccd1 vccd1 _5278_/Y sky130_fd_sc_hd__nor2_2
X_4229_ _4174_/A _4174_/B _4228_/Y _4172_/X _4167_/Y vssd1 vssd1 vccd1 vccd1 _4229_/X
+ sky130_fd_sc_hd__o32a_2
X_7017_ _7036_/B _7017_/B vssd1 vssd1 vccd1 vccd1 _7055_/B sky130_fd_sc_hd__nand2_2
XFILLER_101_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7919_ _6636_/Y _7717_/A _7773_/X vssd1 vssd1 vccd1 vccd1 _7921_/B sky130_fd_sc_hd__a21o_1
XFILLER_15_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4580_ _4581_/B _4583_/A _4581_/A vssd1 vssd1 vccd1 vccd1 _4580_/X sky130_fd_sc_hd__o21a_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6250_ _6250_/A _6250_/B vssd1 vssd1 vccd1 vccd1 _6250_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6181_ _6175_/B _6180_/X _6156_/A vssd1 vssd1 vccd1 vccd1 _6181_/Y sky130_fd_sc_hd__o21ai_1
X_5201_ _5103_/B _5245_/A _5255_/A _5255_/B vssd1 vssd1 vccd1 vccd1 _5202_/B sky130_fd_sc_hd__a22oi_4
X_5132_ _4098_/B _5134_/A2 _4123_/X _5135_/C1 vssd1 vssd1 vccd1 vccd1 _5133_/B sky130_fd_sc_hd__a211o_2
XFILLER_69_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5063_ _5063_/A _5063_/B vssd1 vssd1 vccd1 vccd1 _5243_/A sky130_fd_sc_hd__xnor2_4
XFILLER_38_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4014_ _8011_/Q _8008_/Q _4016_/S vssd1 vssd1 vccd1 vccd1 _8008_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5965_ _5961_/A _5961_/B _5964_/X vssd1 vssd1 vccd1 vccd1 _5970_/B sky130_fd_sc_hd__o21a_1
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7704_ _7607_/A _7697_/Y _7760_/B vssd1 vssd1 vccd1 vccd1 _7706_/A sky130_fd_sc_hd__a21oi_1
X_4916_ _4916_/A _4916_/B vssd1 vssd1 vccd1 vccd1 _4945_/A sky130_fd_sc_hd__xor2_4
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5896_ _5896_/A _5896_/B _5896_/C vssd1 vssd1 vccd1 vccd1 _5912_/A sky130_fd_sc_hd__or3_2
X_7635_ _8029_/Q _7879_/B _7562_/B vssd1 vssd1 vccd1 vccd1 _7635_/X sky130_fd_sc_hd__a21bo_1
X_4847_ _4732_/X _4844_/X _4873_/B _4929_/A _5041_/D1 vssd1 vssd1 vccd1 vccd1 _4847_/X
+ sky130_fd_sc_hd__a2111o_4
X_7566_ _7831_/A _6264_/X _6265_/X _6260_/Y vssd1 vssd1 vccd1 vccd1 _7611_/C sky130_fd_sc_hd__o211a_4
X_4778_ _4800_/A _4778_/B vssd1 vssd1 vccd1 vccd1 _4779_/B sky130_fd_sc_hd__and2_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6517_ _6517_/A _6517_/B vssd1 vssd1 vccd1 vccd1 _6709_/A sky130_fd_sc_hd__xnor2_4
X_7497_ _7483_/X _7496_/X _7515_/S vssd1 vssd1 vccd1 vccd1 _7535_/B sky130_fd_sc_hd__mux2_1
X_6448_ _7366_/B _7366_/A _6448_/S vssd1 vssd1 vccd1 vccd1 _6483_/B sky130_fd_sc_hd__mux2_1
X_6379_ _7195_/B _6878_/C _6445_/S vssd1 vssd1 vccd1 vccd1 _6379_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8049_ _8057_/CLK _8049_/D vssd1 vssd1 vccd1 vccd1 _8049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5750_ _5750_/A _5750_/B _5750_/C vssd1 vssd1 vccd1 vccd1 _5938_/B sky130_fd_sc_hd__or3_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5681_ _5681_/A _5681_/B vssd1 vssd1 vccd1 vccd1 _5730_/A sky130_fd_sc_hd__xor2_4
X_4701_ _4700_/A _4700_/B _4700_/C vssd1 vssd1 vccd1 vccd1 _4703_/B sky130_fd_sc_hd__a21oi_1
X_7420_ _7420_/A _7420_/B vssd1 vssd1 vccd1 vccd1 _7423_/A sky130_fd_sc_hd__xnor2_4
X_4632_ _4632_/A _4641_/A _4632_/C vssd1 vssd1 vccd1 vccd1 _4641_/B sky130_fd_sc_hd__nand3_4
X_7351_ _7351_/A _7351_/B vssd1 vssd1 vccd1 vccd1 _7370_/A sky130_fd_sc_hd__xnor2_4
X_4563_ _4563_/A _4563_/B _4563_/C vssd1 vssd1 vccd1 vccd1 _4599_/A sky130_fd_sc_hd__nand3_2
X_6302_ _6302_/A _6302_/B vssd1 vssd1 vccd1 vccd1 _6303_/B sky130_fd_sc_hd__xor2_4
X_7282_ _7283_/A _7304_/A vssd1 vssd1 vccd1 vccd1 _7282_/Y sky130_fd_sc_hd__nand2_1
X_4494_ _4494_/A _4495_/A _5013_/B vssd1 vssd1 vccd1 vccd1 _4494_/X sky130_fd_sc_hd__or3_2
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6233_ _5927_/C _5925_/Y _5927_/D _5927_/B _7085_/B vssd1 vssd1 vccd1 vccd1 _6233_/X
+ sky130_fd_sc_hd__a32o_1
X_6164_ _6219_/B _6219_/C _6193_/A vssd1 vssd1 vccd1 vccd1 _6164_/Y sky130_fd_sc_hd__a21oi_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6095_ _6096_/A _6096_/B vssd1 vssd1 vccd1 vccd1 _6095_/X sky130_fd_sc_hd__xor2_4
XFILLER_85_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5115_ _5182_/A _5182_/B _5182_/C vssd1 vssd1 vccd1 vccd1 _5183_/A sky130_fd_sc_hd__o21ai_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5046_ _5046_/A _5046_/B vssd1 vssd1 vccd1 vccd1 _5047_/C sky130_fd_sc_hd__xnor2_4
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6997_ _7057_/A _7235_/B _7072_/A vssd1 vssd1 vccd1 vccd1 _6998_/B sky130_fd_sc_hd__o21ai_1
X_5948_ _5476_/Y _6147_/A _5491_/B vssd1 vssd1 vccd1 vccd1 _5948_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5879_ _5879_/A _5879_/B vssd1 vssd1 vccd1 vccd1 _5900_/A sky130_fd_sc_hd__xor2_1
X_7618_ _6732_/B _7617_/Y _7894_/A vssd1 vssd1 vccd1 vccd1 _7620_/B sky130_fd_sc_hd__mux2_2
XFILLER_107_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7549_ _7403_/B _7502_/B _7502_/Y vssd1 vssd1 vccd1 vccd1 _7549_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6920_ _6968_/A _6968_/B _6919_/A vssd1 vssd1 vccd1 vccd1 _6923_/B sky130_fd_sc_hd__a21oi_2
X_6851_ _7101_/A _7057_/A vssd1 vssd1 vccd1 vccd1 _6947_/C sky130_fd_sc_hd__or2_4
Xfanout19 _6629_/Y vssd1 vssd1 vccd1 vccd1 _7583_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_50_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5802_ _5836_/A _5836_/B vssd1 vssd1 vccd1 vccd1 _5837_/A sky130_fd_sc_hd__nand2_2
X_6782_ _6782_/A _6782_/B vssd1 vssd1 vccd1 vccd1 _6788_/A sky130_fd_sc_hd__xor2_4
X_5733_ _5715_/A _5647_/B _5736_/A vssd1 vssd1 vccd1 vccd1 _5733_/Y sky130_fd_sc_hd__o21ai_1
X_5664_ _5714_/A _5842_/B _5714_/C vssd1 vssd1 vccd1 vccd1 _5716_/A sky130_fd_sc_hd__and3_1
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7403_ _7403_/A _7403_/B _7403_/C _7403_/D vssd1 vssd1 vccd1 vccd1 _7421_/A sky130_fd_sc_hd__or4_4
X_5595_ _5589_/A _5587_/Y _5586_/Y vssd1 vssd1 vccd1 vccd1 _5597_/A sky130_fd_sc_hd__o21ai_4
X_4615_ _5014_/A _7001_/A vssd1 vssd1 vccd1 vccd1 _4716_/A sky130_fd_sc_hd__nor2_1
X_7334_ _7334_/A _7334_/B _7344_/B _7371_/B vssd1 vssd1 vccd1 vccd1 _7354_/A sky130_fd_sc_hd__or4_4
X_4546_ _4546_/A _4546_/B vssd1 vssd1 vccd1 vccd1 _4581_/A sky130_fd_sc_hd__xnor2_2
XFILLER_116_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4477_ _4501_/A _4424_/B _4441_/Y _4378_/X _4494_/A vssd1 vssd1 vccd1 vccd1 _4477_/X
+ sky130_fd_sc_hd__a221o_1
X_7265_ _7266_/A _7266_/B vssd1 vssd1 vccd1 vccd1 _7265_/X sky130_fd_sc_hd__or2_1
X_6216_ _6193_/A _6195_/X _6215_/X vssd1 vssd1 vccd1 vccd1 _6216_/X sky130_fd_sc_hd__a21o_1
X_7196_ _7194_/A _7194_/B _7201_/A vssd1 vssd1 vccd1 vccd1 _7198_/B sky130_fd_sc_hd__o21ba_1
X_6147_ _6147_/A _6147_/B vssd1 vssd1 vccd1 vccd1 _6148_/B sky130_fd_sc_hd__nor2_1
XFILLER_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _6078_/A _6078_/B _6078_/C vssd1 vssd1 vccd1 vccd1 _6081_/A sky130_fd_sc_hd__or3_4
XFILLER_73_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5029_ _5030_/A _5030_/B vssd1 vssd1 vccd1 vccd1 _5029_/X sky130_fd_sc_hd__or2_2
XFILLER_72_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4400_ _6999_/A _4412_/B _4602_/A vssd1 vssd1 vccd1 vccd1 _4400_/X sky130_fd_sc_hd__a21o_1
X_5380_ _6800_/B _5853_/B vssd1 vssd1 vccd1 vccd1 _5545_/B sky130_fd_sc_hd__nor2_4
XFILLER_99_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4331_ _4281_/X _4282_/X _4322_/A vssd1 vssd1 vccd1 vccd1 _4334_/A sky130_fd_sc_hd__a21o_1
XFILLER_5_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4262_ _4216_/C _4259_/B _4261_/X _6017_/A vssd1 vssd1 vccd1 vccd1 _4266_/A sky130_fd_sc_hd__a211o_4
X_7050_ _4343_/Y _6951_/D _7045_/Y vssd1 vssd1 vccd1 vccd1 _7051_/B sky130_fd_sc_hd__a21o_1
Xfanout209 _4352_/Y vssd1 vssd1 vccd1 vccd1 _5445_/A sky130_fd_sc_hd__buf_12
XFILLER_113_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6001_ _6007_/A _6317_/A vssd1 vssd1 vccd1 vccd1 _6001_/X sky130_fd_sc_hd__and2_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4193_ _4193_/A _4193_/B vssd1 vssd1 vccd1 vccd1 _4193_/Y sky130_fd_sc_hd__nor2_2
XFILLER_94_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7952_ _7947_/X _7948_/Y _7951_/X _7952_/B1 vssd1 vssd1 vccd1 vccd1 _7954_/B sky130_fd_sc_hd__a31o_1
XFILLER_48_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6903_ _6903_/A _6903_/B _6903_/C _7067_/A vssd1 vssd1 vccd1 vccd1 _6913_/A sky130_fd_sc_hd__or4_4
X_7883_ _7883_/A _7883_/B _7883_/C vssd1 vssd1 vccd1 vccd1 _7909_/B sky130_fd_sc_hd__and3_1
X_6834_ _6834_/A _6834_/B _6834_/C vssd1 vssd1 vccd1 vccd1 _6835_/B sky130_fd_sc_hd__nor3_1
XFILLER_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6765_ _7580_/B _6760_/X _6768_/B vssd1 vssd1 vccd1 vccd1 _7579_/A sky130_fd_sc_hd__a21o_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5716_ _5716_/A _5754_/A vssd1 vssd1 vccd1 vccd1 _5716_/Y sky130_fd_sc_hd__xnor2_1
X_6696_ _6691_/A _6661_/A _6695_/X vssd1 vssd1 vccd1 vccd1 _6696_/X sky130_fd_sc_hd__a21o_1
X_5647_ _6842_/B _5647_/B vssd1 vssd1 vccd1 vccd1 _5692_/B sky130_fd_sc_hd__nor2_8
X_5578_ _5579_/A _5579_/B vssd1 vssd1 vccd1 vccd1 _5580_/A sky130_fd_sc_hd__nor2_2
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7317_ _7329_/A _7329_/B _7314_/Y vssd1 vssd1 vccd1 vccd1 _7327_/B sky130_fd_sc_hd__o21a_2
X_4529_ _4529_/A _4529_/B vssd1 vssd1 vccd1 vccd1 _4530_/B sky130_fd_sc_hd__xnor2_4
X_7248_ _7246_/X _7252_/A vssd1 vssd1 vccd1 vccd1 _7278_/B sky130_fd_sc_hd__and2b_2
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7179_ _7177_/A _7177_/B _7178_/Y vssd1 vssd1 vccd1 vccd1 _7181_/B sky130_fd_sc_hd__o21ai_4
XFILLER_100_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4880_ _4872_/Y _4880_/B vssd1 vssd1 vccd1 vccd1 _4906_/B sky130_fd_sc_hd__nand2b_2
XFILLER_45_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6550_ _7929_/A _6550_/B _6550_/C _6550_/D vssd1 vssd1 vccd1 vccd1 _6552_/A sky130_fd_sc_hd__or4_1
XFILLER_20_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5501_ _6144_/A _6148_/A vssd1 vssd1 vccd1 vccd1 _5502_/B sky130_fd_sc_hd__nand2b_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6481_ _6482_/A _6482_/B vssd1 vssd1 vccd1 vccd1 _6550_/B sky130_fd_sc_hd__nor2_2
X_5432_ _5432_/A _5432_/B _5432_/C vssd1 vssd1 vccd1 vccd1 _5434_/A sky130_fd_sc_hd__and3_2
X_5363_ _5054_/C _5054_/D _5054_/B vssd1 vssd1 vccd1 vccd1 _5364_/B sky130_fd_sc_hd__o21ai_1
XFILLER_113_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4314_ _6035_/A0 _4313_/X _4356_/A vssd1 vssd1 vccd1 vccd1 _4314_/Y sky130_fd_sc_hd__o21ai_2
X_7102_ _7102_/A _7102_/B vssd1 vssd1 vccd1 vccd1 _7107_/B sky130_fd_sc_hd__xnor2_2
X_8082_ _8082_/CLK _8082_/D vssd1 vssd1 vccd1 vccd1 _8082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5294_ _5294_/A _5294_/B vssd1 vssd1 vccd1 vccd1 _5296_/A sky130_fd_sc_hd__xor2_4
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4245_ _6289_/B _6017_/A _4244_/Y _6035_/A0 vssd1 vssd1 vccd1 vccd1 _4245_/X sky130_fd_sc_hd__a211o_1
X_7033_ _7034_/A _7034_/B vssd1 vssd1 vccd1 vccd1 _7035_/A sky130_fd_sc_hd__or2_1
X_4176_ _8072_/Q _8071_/Q _4175_/B _4211_/B vssd1 vssd1 vccd1 vccd1 _4185_/B sky130_fd_sc_hd__o31a_2
XFILLER_27_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7935_ _7935_/A _7935_/B vssd1 vssd1 vccd1 vccd1 _7935_/Y sky130_fd_sc_hd__nand2_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7866_ _7895_/A _7895_/B vssd1 vssd1 vccd1 vccd1 _7867_/B sky130_fd_sc_hd__nor2_1
X_6817_ _6806_/A _7025_/A _6807_/A _6810_/A vssd1 vssd1 vccd1 vccd1 _6820_/A sky130_fd_sc_hd__o31a_4
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7797_ _7889_/A _7797_/B vssd1 vssd1 vccd1 vccd1 _7798_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6748_ _6623_/A _6723_/X _6622_/A vssd1 vssd1 vccd1 vccd1 _6748_/X sky130_fd_sc_hd__a21o_1
X_6679_ _6691_/A _6679_/B vssd1 vssd1 vccd1 vccd1 _6679_/X sky130_fd_sc_hd__and2b_1
XFILLER_2_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4030_ _8019_/Q _8020_/Q _7955_/S vssd1 vssd1 vccd1 vccd1 _8020_/D sky130_fd_sc_hd__mux2_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5981_ _4062_/B _5993_/B _4297_/X _6021_/A0 vssd1 vssd1 vccd1 vccd1 _5981_/X sky130_fd_sc_hd__a211o_1
XFILLER_24_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7720_ _7720_/A _7720_/B vssd1 vssd1 vccd1 vccd1 _7720_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_92_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4932_ _4998_/A _5040_/B vssd1 vssd1 vccd1 vccd1 _4933_/B sky130_fd_sc_hd__nand2_2
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7651_ _7651_/A vssd1 vssd1 vccd1 vccd1 _7651_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6602_ _6602_/A _6602_/B vssd1 vssd1 vccd1 vccd1 _6635_/A sky130_fd_sc_hd__or2_4
X_4863_ _4860_/Y _4863_/B vssd1 vssd1 vccd1 vccd1 _5058_/A sky130_fd_sc_hd__nand2b_2
XFILLER_119_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7582_ _7582_/A vssd1 vssd1 vccd1 vccd1 _7582_/Y sky130_fd_sc_hd__inv_2
X_4794_ _4795_/A _4795_/C vssd1 vssd1 vccd1 vccd1 _4949_/A sky130_fd_sc_hd__nor2_4
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6533_ _6533_/A _6533_/B vssd1 vssd1 vccd1 vccd1 _6538_/A sky130_fd_sc_hd__xor2_4
XFILLER_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6464_ _6463_/X _6527_/A vssd1 vssd1 vccd1 vccd1 _6464_/Y sky130_fd_sc_hd__nand2b_1
X_5415_ _5357_/A _5357_/B _5355_/Y vssd1 vssd1 vccd1 vccd1 _5421_/A sky130_fd_sc_hd__a21bo_4
X_6395_ _7123_/A _5842_/B _6456_/S vssd1 vssd1 vccd1 vccd1 _6397_/B sky130_fd_sc_hd__mux2_2
XFILLER_114_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5346_ _5346_/A _5346_/B vssd1 vssd1 vccd1 vccd1 _5347_/B sky130_fd_sc_hd__xor2_4
X_8065_ _8065_/CLK _8065_/D vssd1 vssd1 vccd1 vccd1 _8065_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5277_ _5482_/A _5482_/B _5261_/X vssd1 vssd1 vccd1 vccd1 _5280_/B sky130_fd_sc_hd__a21oi_2
XFILLER_87_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4228_ _4228_/A _4228_/B vssd1 vssd1 vccd1 vccd1 _4228_/Y sky130_fd_sc_hd__xnor2_1
X_7016_ _7016_/A _7016_/B vssd1 vssd1 vccd1 vccd1 _7017_/B sky130_fd_sc_hd__or2_1
XFILLER_101_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4159_ _6326_/B _6289_/B _4242_/A vssd1 vssd1 vccd1 vccd1 _4159_/Y sky130_fd_sc_hd__nand3_4
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7918_ _7918_/A _7918_/B _7939_/B vssd1 vssd1 vccd1 vccd1 _7918_/X sky130_fd_sc_hd__or3b_1
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7849_ _7766_/A _7766_/B _7848_/A _7848_/B _7872_/A vssd1 vssd1 vccd1 vccd1 _7874_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6180_ _6180_/A _6180_/B _6180_/C vssd1 vssd1 vccd1 vccd1 _6180_/X sky130_fd_sc_hd__and3_1
X_5200_ _5200_/A _5200_/B vssd1 vssd1 vccd1 vccd1 _5255_/B sky130_fd_sc_hd__xnor2_4
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5131_ _6274_/A _5134_/A2 _4132_/X _4303_/B vssd1 vssd1 vccd1 vccd1 _5133_/A sky130_fd_sc_hd__a211o_2
X_5062_ _5062_/A _5062_/B vssd1 vssd1 vccd1 vccd1 _5063_/B sky130_fd_sc_hd__nand2_4
X_4013_ _7974_/A _4013_/B _7991_/D vssd1 vssd1 vccd1 vccd1 _4016_/S sky130_fd_sc_hd__or3b_4
XFILLER_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7703_ _7703_/A _7703_/B vssd1 vssd1 vccd1 vccd1 _7760_/B sky130_fd_sc_hd__xnor2_4
X_5964_ _5226_/Y _7558_/A _5960_/A _5956_/A vssd1 vssd1 vccd1 vccd1 _5964_/X sky130_fd_sc_hd__o211a_1
X_4915_ _4915_/A _4915_/B vssd1 vssd1 vccd1 vccd1 _5290_/A sky130_fd_sc_hd__or2_4
X_5895_ _5893_/A _5893_/B _5901_/A vssd1 vssd1 vccd1 vccd1 _5896_/C sky130_fd_sc_hd__a21oi_1
X_7634_ _7923_/A _7621_/Y _7622_/X _7903_/B1 vssd1 vssd1 vccd1 vccd1 _7634_/X sky130_fd_sc_hd__a31o_1
X_4846_ _4846_/A _4846_/B vssd1 vssd1 vccd1 vccd1 _4873_/B sky130_fd_sc_hd__xor2_4
X_7565_ _7928_/A _7565_/B vssd1 vssd1 vccd1 vccd1 _8028_/D sky130_fd_sc_hd__nor2_1
XFILLER_20_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6516_ _6467_/Y _6510_/Y _7728_/A vssd1 vssd1 vccd1 vccd1 _6517_/B sky130_fd_sc_hd__mux2_4
X_4777_ _4800_/A _4792_/A _4778_/B vssd1 vssd1 vccd1 vccd1 _4779_/A sky130_fd_sc_hd__a21oi_1
XFILLER_119_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7496_ _7475_/X _7478_/X _7527_/S vssd1 vssd1 vccd1 vccd1 _7496_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6447_ _6447_/A _6447_/B vssd1 vssd1 vccd1 vccd1 _6480_/B sky130_fd_sc_hd__nand2_1
X_6378_ _6523_/A vssd1 vssd1 vccd1 vccd1 _6378_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5329_ _5352_/A _5352_/B _7281_/C vssd1 vssd1 vccd1 vccd1 _5330_/B sky130_fd_sc_hd__and3_4
X_8048_ _8057_/CLK _8048_/D vssd1 vssd1 vccd1 vccd1 _8048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _5681_/A _5681_/B vssd1 vssd1 vccd1 vccd1 _5680_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4700_ _4700_/A _4700_/B _4700_/C vssd1 vssd1 vccd1 vccd1 _4709_/B sky130_fd_sc_hd__and3_2
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4631_ _7285_/A _5020_/A _5040_/A _4551_/A vssd1 vssd1 vccd1 vccd1 _4632_/C sky130_fd_sc_hd__a22o_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7350_ _7350_/A _7350_/B vssd1 vssd1 vccd1 vccd1 _7359_/A sky130_fd_sc_hd__xnor2_2
X_4562_ _4561_/B _4561_/C _4561_/A vssd1 vssd1 vccd1 vccd1 _4563_/C sky130_fd_sc_hd__a21o_1
X_6301_ _6047_/X _6050_/Y _6767_/S vssd1 vssd1 vccd1 vccd1 _6302_/B sky130_fd_sc_hd__mux2_8
X_7281_ _7281_/A _7281_/B _7281_/C _7281_/D vssd1 vssd1 vccd1 vccd1 _7304_/A sky130_fd_sc_hd__and4_4
X_4493_ _4494_/A _4642_/B vssd1 vssd1 vccd1 vccd1 _4495_/B sky130_fd_sc_hd__nor2_2
XFILLER_89_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6232_ _6146_/A _6240_/A _6231_/Y _6242_/S vssd1 vssd1 vccd1 vccd1 _6232_/Y sky130_fd_sc_hd__o22ai_2
X_6163_ _6259_/A _6192_/B _6192_/C _6163_/D vssd1 vssd1 vccd1 vccd1 _6219_/C sky130_fd_sc_hd__or4_1
XFILLER_69_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6094_ _6084_/A _6045_/X _6071_/A vssd1 vssd1 vccd1 vccd1 _6096_/B sky130_fd_sc_hd__a21oi_4
XFILLER_84_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5114_ _5182_/A _5182_/B _5182_/C vssd1 vssd1 vccd1 vccd1 _5114_/X sky130_fd_sc_hd__o21a_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5037_/Y _5039_/Y _5042_/Y _5044_/X vssd1 vssd1 vccd1 vccd1 _5047_/B sky130_fd_sc_hd__a31o_2
XFILLER_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6996_ _6996_/A _6996_/B vssd1 vssd1 vccd1 vccd1 _7036_/A sky130_fd_sc_hd__xnor2_1
X_5947_ _5947_/A _6135_/A _5944_/Y _5615_/Y vssd1 vssd1 vccd1 vccd1 _5951_/B sky130_fd_sc_hd__or4bb_2
XFILLER_25_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7617_ _7617_/A vssd1 vssd1 vccd1 vccd1 _7617_/Y sky130_fd_sc_hd__inv_2
X_5878_ _5869_/A _5868_/C _5868_/A vssd1 vssd1 vccd1 vccd1 _5893_/B sky130_fd_sc_hd__a21o_1
X_4829_ _4829_/A _4829_/B _4833_/A vssd1 vssd1 vccd1 vccd1 _4830_/B sky130_fd_sc_hd__or3_2
X_7548_ _7554_/B _7541_/Y _7547_/Y _7554_/A vssd1 vssd1 vccd1 vccd1 _7553_/B sky130_fd_sc_hd__a31o_1
X_7479_ _7477_/X _7439_/X _7479_/S vssd1 vssd1 vccd1 vccd1 _7479_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6850_ _6862_/A _6850_/B vssd1 vssd1 vccd1 vccd1 _6863_/A sky130_fd_sc_hd__or2_4
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6781_ _5151_/C _6783_/B _6780_/Y vssd1 vssd1 vccd1 vccd1 _6782_/B sky130_fd_sc_hd__o21ai_4
X_5801_ _5736_/C _5798_/C _5799_/Y _5800_/X vssd1 vssd1 vccd1 vccd1 _5836_/B sky130_fd_sc_hd__o211a_1
X_5732_ _5732_/A _5732_/B vssd1 vssd1 vccd1 vccd1 _5776_/A sky130_fd_sc_hd__xor2_4
X_5663_ _5663_/A _5663_/B vssd1 vssd1 vccd1 vccd1 _5670_/B sky130_fd_sc_hd__xnor2_1
X_7402_ _7402_/A _7513_/S vssd1 vssd1 vccd1 vccd1 _7403_/D sky130_fd_sc_hd__xnor2_4
X_5594_ _5594_/A _5692_/A vssd1 vssd1 vccd1 vccd1 _5650_/A sky130_fd_sc_hd__or2_4
X_4614_ _4614_/A _4614_/B vssd1 vssd1 vccd1 vccd1 _4846_/A sky130_fd_sc_hd__xnor2_4
X_7333_ _7366_/A _7371_/B vssd1 vssd1 vccd1 vccd1 _7333_/Y sky130_fd_sc_hd__nor2_1
X_4545_ _4545_/A _4545_/B vssd1 vssd1 vccd1 vccd1 _4738_/A sky130_fd_sc_hd__xnor2_4
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4476_ _4406_/A _4441_/A _7311_/A _4475_/X vssd1 vssd1 vccd1 vccd1 _4476_/X sky130_fd_sc_hd__a22o_1
X_7264_ _7276_/A _7276_/B _7259_/X vssd1 vssd1 vccd1 vccd1 _7266_/B sky130_fd_sc_hd__a21oi_2
X_6215_ _6012_/A _6113_/X _6213_/X _6254_/S vssd1 vssd1 vccd1 vccd1 _6215_/X sky130_fd_sc_hd__o211a_1
X_7195_ _7319_/A _7195_/B _7195_/C vssd1 vssd1 vccd1 vccd1 _7201_/A sky130_fd_sc_hd__and3_2
XFILLER_112_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6146_ _6146_/A _6146_/B vssd1 vssd1 vccd1 vccd1 _6146_/X sky130_fd_sc_hd__or2_1
XFILLER_38_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _6077_/A _6077_/B vssd1 vssd1 vccd1 vccd1 _7639_/A sky130_fd_sc_hd__nand2_8
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5028_ _5046_/A _5046_/B _5026_/X vssd1 vssd1 vccd1 vccd1 _5030_/B sky130_fd_sc_hd__a21oi_4
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6979_ _6983_/B _6979_/B vssd1 vssd1 vccd1 vccd1 _6994_/B sky130_fd_sc_hd__and2_1
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4330_ _4266_/X _4328_/Y _4327_/X _6034_/A vssd1 vssd1 vccd1 vccd1 _4330_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4261_ _4241_/B _4227_/X _4231_/X _4221_/B vssd1 vssd1 vccd1 vccd1 _4261_/X sky130_fd_sc_hd__o211a_1
X_6000_ _6000_/A _6000_/B vssd1 vssd1 vccd1 vccd1 _7398_/A sky130_fd_sc_hd__or2_4
X_4192_ _4216_/B _4192_/B vssd1 vssd1 vccd1 vccd1 _4192_/X sky130_fd_sc_hd__xor2_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7951_ _6188_/A _6805_/B _6354_/A _7939_/A _7950_/Y vssd1 vssd1 vccd1 vccd1 _7951_/X
+ sky130_fd_sc_hd__a221o_1
X_7882_ _7831_/A _7667_/Y _7908_/A vssd1 vssd1 vccd1 vccd1 _7883_/C sky130_fd_sc_hd__a21oi_4
XFILLER_70_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6902_ _6902_/A _7235_/B vssd1 vssd1 vccd1 vccd1 _7067_/A sky130_fd_sc_hd__or2_4
X_6833_ _6833_/A _6833_/B vssd1 vssd1 vccd1 vccd1 _6861_/A sky130_fd_sc_hd__and2_2
XFILLER_62_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6764_ _6744_/Y _6763_/X _7718_/S vssd1 vssd1 vccd1 vccd1 _6768_/B sky130_fd_sc_hd__mux2_2
XFILLER_50_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6695_ _6694_/X _6683_/X _6695_/S vssd1 vssd1 vccd1 vccd1 _6695_/X sky130_fd_sc_hd__mux2_1
X_5715_ _5715_/A _5880_/A vssd1 vssd1 vccd1 vccd1 _5754_/A sky130_fd_sc_hd__or2_2
X_5646_ _6842_/B _5853_/B vssd1 vssd1 vccd1 vccd1 _5736_/A sky130_fd_sc_hd__or2_2
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5577_ _5635_/A _5635_/B _5570_/A vssd1 vssd1 vccd1 vccd1 _5579_/B sky130_fd_sc_hd__a21oi_2
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7316_ _7316_/A _7316_/B vssd1 vssd1 vccd1 vccd1 _7329_/B sky130_fd_sc_hd__xnor2_2
X_4528_ _4528_/A _4528_/B vssd1 vssd1 vccd1 vccd1 _4529_/B sky130_fd_sc_hd__nand2_2
X_7247_ _7247_/A _7334_/B _7247_/C _7247_/D vssd1 vssd1 vccd1 vccd1 _7252_/A sky130_fd_sc_hd__or4_4
X_4459_ _4457_/A _4503_/A _4458_/X vssd1 vssd1 vccd1 vccd1 _4460_/B sky130_fd_sc_hd__o21ai_4
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7178_ _7204_/A _7204_/B vssd1 vssd1 vccd1 vccd1 _7178_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_85_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6129_ _6081_/Y _6111_/B _6111_/C _6192_/D vssd1 vssd1 vccd1 vccd1 _6129_/X sky130_fd_sc_hd__a31o_1
XFILLER_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5500_ _6155_/A _6159_/A vssd1 vssd1 vccd1 vccd1 _5502_/A sky130_fd_sc_hd__or2_1
XFILLER_9_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6480_ _6446_/Y _6480_/B vssd1 vssd1 vccd1 vccd1 _6545_/A sky130_fd_sc_hd__and2b_4
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5431_ _5431_/A _5431_/B vssd1 vssd1 vccd1 vccd1 _5432_/C sky130_fd_sc_hd__xnor2_2
XFILLER_114_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5362_ _5986_/S _5362_/B vssd1 vssd1 vccd1 vccd1 _5362_/Y sky130_fd_sc_hd__nand2_2
XFILLER_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8081_ _8082_/CLK _8081_/D vssd1 vssd1 vccd1 vccd1 _8081_/Q sky130_fd_sc_hd__dfxtp_4
X_4313_ _4272_/Y _4276_/X _6017_/A vssd1 vssd1 vccd1 vccd1 _4313_/X sky130_fd_sc_hd__mux2_1
X_7101_ _7101_/A _7371_/A vssd1 vssd1 vccd1 vccd1 _7107_/A sky130_fd_sc_hd__or2_2
XFILLER_113_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5293_ _6878_/B _5338_/B vssd1 vssd1 vccd1 vccd1 _5294_/B sky130_fd_sc_hd__nand2_8
X_7032_ _7079_/A _7079_/B _7029_/X vssd1 vssd1 vccd1 vccd1 _7034_/B sky130_fd_sc_hd__a21oi_1
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4244_ _4244_/A _4244_/B vssd1 vssd1 vccd1 vccd1 _4244_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4175_ _4211_/B _4175_/B vssd1 vssd1 vccd1 vccd1 _4194_/B sky130_fd_sc_hd__nand2_2
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7934_ _7934_/A _7934_/B vssd1 vssd1 vccd1 vccd1 _7934_/X sky130_fd_sc_hd__or2_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7865_ _7895_/A _7895_/B vssd1 vssd1 vccd1 vccd1 _7867_/A sky130_fd_sc_hd__and2_1
XFILLER_82_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7796_ _7837_/A _7874_/A vssd1 vssd1 vccd1 vccd1 _7801_/A sky130_fd_sc_hd__nand2_2
X_6816_ _6835_/A _6832_/B vssd1 vssd1 vccd1 vccd1 _6833_/A sky130_fd_sc_hd__nand2_2
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6747_ _6745_/X _6746_/X _6749_/S vssd1 vssd1 vccd1 vccd1 _6757_/C sky130_fd_sc_hd__mux2_1
X_6678_ _6677_/Y _6666_/A _6695_/S vssd1 vssd1 vccd1 vccd1 _6679_/B sky130_fd_sc_hd__mux2_1
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5629_ _5722_/A _5722_/B _5919_/A vssd1 vssd1 vccd1 vccd1 _5632_/B sky130_fd_sc_hd__and3_2
XFILLER_117_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5980_ _6349_/B _6010_/B _5972_/Y vssd1 vssd1 vccd1 vccd1 _5987_/B sky130_fd_sc_hd__a21oi_4
XFILLER_37_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4931_ _4931_/A _4931_/B vssd1 vssd1 vccd1 vccd1 _4933_/A sky130_fd_sc_hd__nand2_4
X_7650_ _7616_/S _6762_/X _6631_/X vssd1 vssd1 vccd1 vccd1 _7651_/A sky130_fd_sc_hd__a21o_1
X_4862_ _4863_/B vssd1 vssd1 vccd1 vccd1 _4862_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6601_ _6601_/A _6601_/B _6627_/A vssd1 vssd1 vccd1 vccd1 _6602_/B sky130_fd_sc_hd__and3_1
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7581_ _6761_/Y _7773_/A _7581_/S vssd1 vssd1 vccd1 vccd1 _7582_/A sky130_fd_sc_hd__mux2_1
X_4793_ _4795_/B _4795_/C _4820_/S _4772_/Y vssd1 vssd1 vccd1 vccd1 _4793_/X sky130_fd_sc_hd__o211a_1
XFILLER_119_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6532_ _6544_/S _6504_/Y _6531_/Y vssd1 vssd1 vccd1 vccd1 _6533_/B sky130_fd_sc_hd__a21oi_4
X_6463_ _6406_/X _6462_/Y _6474_/B vssd1 vssd1 vccd1 vccd1 _6463_/X sky130_fd_sc_hd__o21a_1
X_5414_ _5414_/A _5414_/B vssd1 vssd1 vccd1 vccd1 _5423_/A sky130_fd_sc_hd__xor2_4
X_6394_ _6443_/A _6394_/B vssd1 vssd1 vccd1 vccd1 _6397_/A sky130_fd_sc_hd__nand2_1
XFILLER_114_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5345_ _5346_/A _5346_/B vssd1 vssd1 vccd1 vccd1 _5403_/A sky130_fd_sc_hd__nand2_2
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8064_ _8065_/CLK _8064_/D vssd1 vssd1 vccd1 vccd1 _8064_/Q sky130_fd_sc_hd__dfxtp_4
X_5276_ _5276_/A _5466_/A vssd1 vssd1 vccd1 vccd1 _5482_/B sky130_fd_sc_hd__xor2_4
XFILLER_101_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4227_ _4223_/Y _4224_/Y _4227_/S vssd1 vssd1 vccd1 vccd1 _4227_/X sky130_fd_sc_hd__mux2_4
X_7015_ _7015_/A _7015_/B vssd1 vssd1 vccd1 vccd1 _7055_/A sky130_fd_sc_hd__xnor2_4
XFILLER_101_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4158_ _4228_/A _6289_/B _4242_/A vssd1 vssd1 vccd1 vccd1 _4158_/X sky130_fd_sc_hd__or3_4
X_4089_ _8056_/Q _8055_/Q _4096_/B _4096_/A vssd1 vssd1 vccd1 vccd1 _4090_/B sky130_fd_sc_hd__o31a_2
X_7917_ _7917_/A _7917_/B vssd1 vssd1 vccd1 vccd1 _7918_/A sky130_fd_sc_hd__nor2_1
XFILLER_102_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7848_ _7848_/A _7848_/B vssd1 vssd1 vccd1 vccd1 _7872_/A sky130_fd_sc_hd__nand2_2
XFILLER_51_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7779_ _7935_/A _7743_/A _7777_/Y _7778_/Y _6774_/X vssd1 vssd1 vccd1 vccd1 _7779_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_11_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5130_ _5367_/A _5386_/A vssd1 vssd1 vccd1 vccd1 _5369_/A sky130_fd_sc_hd__nor2_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5061_ _4814_/B _5074_/B _4831_/X _5071_/B _4812_/Y vssd1 vssd1 vccd1 vccd1 _5062_/B
+ sky130_fd_sc_hd__o221a_2
X_4012_ _4008_/X _4009_/X _7961_/A vssd1 vssd1 vccd1 vccd1 _4013_/B sky130_fd_sc_hd__o21ai_1
XFILLER_97_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5963_ _6180_/A _6180_/B _6180_/C vssd1 vssd1 vccd1 vccd1 _5970_/A sky130_fd_sc_hd__a21o_1
XFILLER_65_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7702_ _7702_/A _7702_/B _7757_/D vssd1 vssd1 vccd1 vccd1 _7702_/X sky130_fd_sc_hd__or3b_1
X_4914_ _4914_/A _4914_/B _4914_/C vssd1 vssd1 vccd1 vccd1 _4915_/B sky130_fd_sc_hd__and3_1
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5894_ _7281_/C _5927_/B vssd1 vssd1 vccd1 vccd1 _5896_/B sky130_fd_sc_hd__nand2_1
X_7633_ _7929_/A _7656_/A _7656_/B _7632_/Y vssd1 vssd1 vccd1 vccd1 _7633_/X sky130_fd_sc_hd__o31a_1
X_4845_ _4732_/X _4844_/X _5041_/D1 _4929_/A vssd1 vssd1 vccd1 vccd1 _4897_/A sky130_fd_sc_hd__a211o_4
XFILLER_20_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7564_ _8028_/Q _7857_/B _7561_/X _7562_/B vssd1 vssd1 vccd1 vccd1 _7565_/B sky130_fd_sc_hd__o2bb2a_1
X_4776_ _4447_/Y _4751_/C _4775_/A _4775_/B vssd1 vssd1 vccd1 vccd1 _4778_/B sky130_fd_sc_hd__a22oi_2
XFILLER_119_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6515_ _6739_/S _6515_/B vssd1 vssd1 vccd1 vccd1 _6515_/Y sky130_fd_sc_hd__nand2b_2
X_7495_ _7542_/A vssd1 vssd1 vccd1 vccd1 _7495_/Y sky130_fd_sc_hd__inv_2
X_6446_ _6447_/A _6447_/B vssd1 vssd1 vccd1 vccd1 _6446_/Y sky130_fd_sc_hd__nor2_1
X_6377_ _6377_/A _6377_/B vssd1 vssd1 vccd1 vccd1 _6523_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5328_ _5582_/A _5800_/A vssd1 vssd1 vccd1 vccd1 _5353_/A sky130_fd_sc_hd__or2_4
X_8047_ _8057_/CLK _8047_/D vssd1 vssd1 vccd1 vccd1 _8047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5259_ _5259_/A _5259_/B vssd1 vssd1 vccd1 vccd1 _5459_/B sky130_fd_sc_hd__xnor2_4
XFILLER_113_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout190 _4244_/A vssd1 vssd1 vccd1 vccd1 _6017_/A sky130_fd_sc_hd__buf_6
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4630_ _4654_/A _4630_/B _4630_/C vssd1 vssd1 vccd1 vccd1 _4641_/A sky130_fd_sc_hd__or3_4
X_6300_ _6299_/A _6564_/A _6305_/A _6304_/A vssd1 vssd1 vccd1 vccd1 _6302_/A sky130_fd_sc_hd__a31o_4
X_4561_ _4561_/A _4561_/B _4561_/C vssd1 vssd1 vccd1 vccd1 _4563_/B sky130_fd_sc_hd__nand3_2
X_7280_ _7311_/A _7294_/B _7311_/C _7279_/X vssd1 vssd1 vccd1 vccd1 _7283_/A sky130_fd_sc_hd__o31a_4
X_4492_ _4360_/A _4487_/X _4490_/X _4570_/A vssd1 vssd1 vccd1 vccd1 _5034_/A sky130_fd_sc_hd__a31o_4
X_6231_ _6231_/A vssd1 vssd1 vccd1 vccd1 _6231_/Y sky130_fd_sc_hd__inv_2
X_6162_ _6081_/Y _6111_/B _6111_/C _6161_/Y vssd1 vssd1 vccd1 vccd1 _6219_/B sky130_fd_sc_hd__a31o_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5113_/A _5113_/B vssd1 vssd1 vccd1 vccd1 _5182_/C sky130_fd_sc_hd__xor2_4
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6093_ _6110_/A _6093_/B _6132_/B vssd1 vssd1 vccd1 vccd1 _6093_/X sky130_fd_sc_hd__or3_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5037_/Y _5042_/Y _5043_/Y vssd1 vssd1 vccd1 vccd1 _5044_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6995_ _6995_/A _6995_/B vssd1 vssd1 vccd1 vccd1 _7041_/A sky130_fd_sc_hd__nand2_4
X_5946_ _5947_/A _5946_/B vssd1 vssd1 vccd1 vccd1 _5951_/A sky130_fd_sc_hd__nand2b_1
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5877_ _5877_/A _5877_/B vssd1 vssd1 vccd1 vccd1 _5897_/A sky130_fd_sc_hd__xor2_1
X_7616_ _6632_/X _6725_/Y _7616_/S vssd1 vssd1 vccd1 vccd1 _7617_/A sky130_fd_sc_hd__mux2_2
X_4828_ _4829_/B _4833_/A _4829_/A vssd1 vssd1 vccd1 vccd1 _5074_/B sky130_fd_sc_hd__o21ai_4
XFILLER_21_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7547_ _7536_/X _7537_/X _7546_/X vssd1 vssd1 vccd1 vccd1 _7547_/Y sky130_fd_sc_hd__a21oi_1
X_4759_ _5090_/B _4759_/B vssd1 vssd1 vccd1 vccd1 _4761_/B sky130_fd_sc_hd__nand2_1
X_7478_ _7474_/X _7477_/X _7513_/S vssd1 vssd1 vccd1 vccd1 _7478_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6429_ _6475_/A _6429_/B vssd1 vssd1 vccd1 vccd1 _6476_/B sky130_fd_sc_hd__or2_2
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6780_ _6780_/A _6791_/B vssd1 vssd1 vccd1 vccd1 _6780_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5800_ _5800_/A _5919_/A _5855_/B _5800_/D vssd1 vssd1 vccd1 vccd1 _5800_/X sky130_fd_sc_hd__or4_1
XFILLER_35_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5731_ _5732_/A _5732_/B vssd1 vssd1 vccd1 vccd1 _5731_/Y sky130_fd_sc_hd__nor2_1
X_5662_ _5662_/A _5662_/B vssd1 vssd1 vccd1 vccd1 _5706_/A sky130_fd_sc_hd__xor2_4
X_7401_ _7401_/A _7401_/B vssd1 vssd1 vccd1 vccd1 _7403_/C sky130_fd_sc_hd__xor2_2
X_5593_ _5621_/A _5647_/B vssd1 vssd1 vccd1 vccd1 _5648_/A sky130_fd_sc_hd__or2_1
X_4613_ _4614_/B _4614_/A vssd1 vssd1 vccd1 vccd1 _4613_/X sky130_fd_sc_hd__and2b_2
X_7332_ _7332_/A _7332_/B vssd1 vssd1 vccd1 vccd1 _7352_/A sky130_fd_sc_hd__nor2_2
X_4544_ _4544_/A _4544_/B vssd1 vssd1 vccd1 vccd1 _4545_/B sky130_fd_sc_hd__xnor2_4
X_7263_ _7263_/A _7263_/B vssd1 vssd1 vccd1 vccd1 _7276_/B sky130_fd_sc_hd__xnor2_4
XFILLER_89_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6214_ _6012_/A _6262_/S _6213_/X vssd1 vssd1 vccd1 vccd1 _6214_/X sky130_fd_sc_hd__o21a_1
X_4475_ _4268_/X _7319_/A _4441_/A vssd1 vssd1 vccd1 vccd1 _4475_/X sky130_fd_sc_hd__a21o_1
X_7194_ _7194_/A _7194_/B vssd1 vssd1 vccd1 vccd1 _7195_/C sky130_fd_sc_hd__xor2_2
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6145_ _6147_/B _6145_/B vssd1 vssd1 vccd1 vccd1 _6146_/B sky130_fd_sc_hd__nor2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6078_/B _6078_/C vssd1 vssd1 vccd1 vccd1 _7755_/A sky130_fd_sc_hd__nor2_4
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5027_ _5027_/A _5027_/B vssd1 vssd1 vccd1 vccd1 _5046_/B sky130_fd_sc_hd__xnor2_4
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6978_ _6978_/A _6978_/B _6978_/C vssd1 vssd1 vccd1 vccd1 _6979_/B sky130_fd_sc_hd__nand3_1
XFILLER_41_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5929_ _5924_/A _5924_/B _5928_/X vssd1 vssd1 vccd1 vccd1 _5929_/X sky130_fd_sc_hd__o21ba_1
XFILLER_70_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4260_ _8067_/Q _4315_/B _4260_/C vssd1 vssd1 vccd1 vccd1 _4260_/X sky130_fd_sc_hd__and3_1
XFILLER_69_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4191_ _4216_/B _4192_/B vssd1 vssd1 vccd1 vccd1 _4193_/B sky130_fd_sc_hd__xnor2_2
XFILLER_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7950_ _8009_/Q _6770_/Y _7949_/Y _8010_/Q vssd1 vssd1 vccd1 vccd1 _7950_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_67_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7881_ _7857_/Y _7880_/X _7928_/A vssd1 vssd1 vccd1 vccd1 _8039_/D sky130_fd_sc_hd__a21oi_1
XFILLER_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6901_ _7012_/A _7124_/A2 _7046_/B _6902_/A vssd1 vssd1 vccd1 vccd1 _6903_/C sky130_fd_sc_hd__o22a_1
X_6832_ _6835_/A _6832_/B vssd1 vssd1 vccd1 vccd1 _6833_/B sky130_fd_sc_hd__or2_1
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6763_ _6730_/Y _6762_/X _7583_/S vssd1 vssd1 vccd1 vccd1 _6763_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6694_ _6524_/B _6524_/A _6737_/B vssd1 vssd1 vccd1 vccd1 _6694_/X sky130_fd_sc_hd__mux2_1
X_5714_ _5714_/A _7269_/B _5714_/C vssd1 vssd1 vccd1 vccd1 _5714_/X sky130_fd_sc_hd__and3_1
X_5645_ _5645_/A _5645_/B vssd1 vssd1 vccd1 vccd1 _5697_/A sky130_fd_sc_hd__xnor2_4
XFILLER_40_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5576_ _5576_/A _5576_/B vssd1 vssd1 vccd1 vccd1 _5635_/B sky130_fd_sc_hd__xnor2_4
XFILLER_117_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7315_ _7312_/A _7336_/A _7309_/Y vssd1 vssd1 vccd1 vccd1 _7329_/A sky130_fd_sc_hd__o21a_2
XFILLER_2_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4527_ _4642_/A _7116_/A _5090_/A _4920_/A vssd1 vssd1 vccd1 vccd1 _4528_/B sky130_fd_sc_hd__or4b_1
XFILLER_116_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7246_ _7334_/B _7247_/C _7247_/D _7247_/A vssd1 vssd1 vccd1 vccd1 _7246_/X sky130_fd_sc_hd__o22a_1
X_4458_ _4551_/A _4456_/B _4585_/B _7319_/A vssd1 vssd1 vccd1 vccd1 _4458_/X sky130_fd_sc_hd__a22o_2
X_7177_ _7177_/A _7177_/B vssd1 vssd1 vccd1 vccd1 _7204_/B sky130_fd_sc_hd__xor2_4
XFILLER_49_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6128_ _5797_/A _6174_/A _6125_/X vssd1 vssd1 vccd1 vccd1 _6192_/D sky130_fd_sc_hd__a21oi_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4389_ _4551_/A _4585_/B vssd1 vssd1 vccd1 vccd1 _4457_/A sky130_fd_sc_hd__nand2_2
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6059_/A _6059_/B vssd1 vssd1 vccd1 vccd1 _6096_/A sky130_fd_sc_hd__or2_4
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5430_ _5346_/A _5346_/B _5403_/B _5412_/A _5412_/B vssd1 vssd1 vccd1 vccd1 _5443_/A
+ sky130_fd_sc_hd__a32oi_4
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5361_ _5986_/S _5362_/B vssd1 vssd1 vccd1 vccd1 _7085_/B sky130_fd_sc_hd__and2_4
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8080_ _8080_/CLK _8080_/D vssd1 vssd1 vccd1 vccd1 _8080_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4312_ _4548_/A _4312_/B _4312_/C vssd1 vssd1 vccd1 vccd1 _4312_/X sky130_fd_sc_hd__and3_2
X_5292_ _6842_/B _5516_/A vssd1 vssd1 vccd1 vccd1 _5294_/A sky130_fd_sc_hd__or2_4
X_7100_ _7102_/A _7102_/B vssd1 vssd1 vccd1 vccd1 _7100_/X sky130_fd_sc_hd__or2_1
X_4243_ _4172_/B _4259_/B _4242_/X vssd1 vssd1 vccd1 vccd1 _4244_/B sky130_fd_sc_hd__o21ai_1
X_7031_ _7031_/A _7031_/B vssd1 vssd1 vccd1 vccd1 _7079_/B sky130_fd_sc_hd__xnor2_4
XFILLER_113_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4174_ _4174_/A _4174_/B vssd1 vssd1 vccd1 vccd1 _4210_/B sky130_fd_sc_hd__nor2_4
XFILLER_67_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7933_ _7911_/B _7929_/X _7931_/X _6269_/X vssd1 vssd1 vccd1 vccd1 _7934_/B sky130_fd_sc_hd__a31o_1
XFILLER_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7864_ _6636_/Y _7651_/A _7773_/X vssd1 vssd1 vccd1 vccd1 _7895_/B sky130_fd_sc_hd__a21oi_1
X_7795_ _7795_/A _7795_/B vssd1 vssd1 vccd1 vccd1 _7874_/A sky130_fd_sc_hd__nand2_2
X_6815_ _6815_/A _6815_/B vssd1 vssd1 vccd1 vccd1 _6832_/B sky130_fd_sc_hd__xnor2_1
X_6746_ _6714_/X _6722_/X _6753_/S vssd1 vssd1 vccd1 vccd1 _6746_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6677_ _6677_/A vssd1 vssd1 vccd1 vccd1 _6677_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5628_ _5672_/A _5855_/A vssd1 vssd1 vccd1 vccd1 _5633_/A sky130_fd_sc_hd__or2_4
X_5559_ _5614_/A _5559_/B vssd1 vssd1 vccd1 vccd1 _5611_/A sky130_fd_sc_hd__and2_2
XFILLER_104_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7229_ _7229_/A _7229_/B vssd1 vssd1 vccd1 vccd1 _7241_/B sky130_fd_sc_hd__xnor2_4
XFILLER_100_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4930_ _4930_/A _4930_/B vssd1 vssd1 vccd1 vccd1 _5033_/B sky130_fd_sc_hd__or2_4
X_4861_ _4860_/B _4860_/C _4860_/A vssd1 vssd1 vccd1 vccd1 _4863_/B sky130_fd_sc_hd__o21ai_2
XFILLER_33_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6600_ _6601_/B _6627_/A _6601_/A vssd1 vssd1 vccd1 vccd1 _6602_/A sky130_fd_sc_hd__a21oi_4
X_7580_ _6768_/B _7580_/B _7580_/C vssd1 vssd1 vccd1 vccd1 _7619_/A sky130_fd_sc_hd__and3b_2
X_4792_ _4792_/A _4792_/B vssd1 vssd1 vccd1 vccd1 _4806_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6531_ _6544_/S _6531_/B vssd1 vssd1 vccd1 vccd1 _6531_/Y sky130_fd_sc_hd__nor2_1
X_6462_ _6533_/A _6531_/B _6415_/X vssd1 vssd1 vccd1 vccd1 _6462_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6393_ _6443_/A _6394_/B vssd1 vssd1 vccd1 vccd1 _6393_/X sky130_fd_sc_hd__and2_1
X_5413_ _5414_/A _5414_/B vssd1 vssd1 vccd1 vccd1 _5413_/Y sky130_fd_sc_hd__nor2_1
X_5344_ _5541_/A _5344_/B vssd1 vssd1 vccd1 vccd1 _5346_/B sky130_fd_sc_hd__nor2_8
XFILLER_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8063_ _8063_/CLK _8063_/D vssd1 vssd1 vccd1 vccd1 _8063_/Q sky130_fd_sc_hd__dfxtp_4
X_5275_ _5275_/A _5464_/B _5275_/C vssd1 vssd1 vccd1 vccd1 _5466_/A sky130_fd_sc_hd__and3_4
XFILLER_101_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4226_ _4222_/X _4225_/X _4227_/S vssd1 vssd1 vccd1 vccd1 _4226_/X sky130_fd_sc_hd__mux2_8
X_7014_ _7013_/B _7013_/C _7013_/A vssd1 vssd1 vccd1 vccd1 _7015_/B sky130_fd_sc_hd__a21bo_4
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4157_ _6326_/B _6289_/B vssd1 vssd1 vccd1 vccd1 _4230_/B sky130_fd_sc_hd__and2_1
XFILLER_110_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4088_ _4088_/A _8053_/Q _8052_/Q _6060_/A vssd1 vssd1 vccd1 vccd1 _4088_/X sky130_fd_sc_hd__or4_1
XFILLER_71_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7916_ _7917_/A _7917_/B vssd1 vssd1 vccd1 vccd1 _7939_/B sky130_fd_sc_hd__nand2_1
XFILLER_70_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7847_ _7847_/A _7847_/B vssd1 vssd1 vccd1 vccd1 _7848_/B sky130_fd_sc_hd__or2_1
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7778_ _7935_/A _7743_/A _7777_/Y vssd1 vssd1 vccd1 vccd1 _7778_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6729_ _6699_/X _6728_/X _6753_/S vssd1 vssd1 vccd1 vccd1 _6730_/A sky130_fd_sc_hd__mux2_2
XFILLER_109_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5060_ _4862_/Y _5189_/B _4860_/Y vssd1 vssd1 vccd1 vccd1 _5071_/B sky130_fd_sc_hd__o21bai_4
X_4011_ _8050_/Q _8045_/Q _7956_/C _8049_/Q vssd1 vssd1 vccd1 vccd1 _7961_/A sky130_fd_sc_hd__nor4b_4
XFILLER_96_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5962_ _6180_/A _6180_/B _6180_/C vssd1 vssd1 vccd1 vccd1 _6175_/B sky130_fd_sc_hd__a21oi_1
X_7701_ _7731_/A _7703_/B vssd1 vssd1 vccd1 vccd1 _7702_/B sky130_fd_sc_hd__nand2b_1
X_4913_ _4915_/A vssd1 vssd1 vccd1 vccd1 _4913_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5893_ _5893_/A _5893_/B _5901_/A vssd1 vssd1 vccd1 vccd1 _5897_/B sky130_fd_sc_hd__nand3_1
X_7632_ _7918_/B _7632_/B vssd1 vssd1 vccd1 vccd1 _7632_/Y sky130_fd_sc_hd__nor2_1
X_4844_ _4702_/Y _4836_/B _4707_/Y _4709_/B vssd1 vssd1 vccd1 vccd1 _4844_/X sky130_fd_sc_hd__a211o_2
XFILLER_20_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7563_ _7944_/B vssd1 vssd1 vccd1 vccd1 _7563_/Y sky130_fd_sc_hd__inv_2
X_4775_ _4775_/A _4775_/B _4800_/A _4775_/D vssd1 vssd1 vccd1 vccd1 _4792_/A sky130_fd_sc_hd__nand4_2
XFILLER_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6514_ _6514_/A _6514_/B vssd1 vssd1 vccd1 vccd1 _6515_/B sky130_fd_sc_hd__xor2_2
XFILLER_20_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7494_ _7531_/B _7493_/X _7535_/A vssd1 vssd1 vccd1 vccd1 _7542_/A sky130_fd_sc_hd__mux2_1
X_6445_ _7284_/A _7210_/B _6445_/S vssd1 vssd1 vccd1 vccd1 _6447_/B sky130_fd_sc_hd__mux2_4
X_6376_ _6376_/A vssd1 vssd1 vccd1 vccd1 _6377_/B sky130_fd_sc_hd__inv_2
XFILLER_114_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5327_ _5294_/A _5518_/A _5311_/B _5307_/X vssd1 vssd1 vccd1 vccd1 _5335_/A sky130_fd_sc_hd__o22ai_4
X_8046_ _8057_/CLK _8046_/D vssd1 vssd1 vccd1 vccd1 _8046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5258_ _5258_/A _5258_/B vssd1 vssd1 vccd1 vccd1 _5459_/A sky130_fd_sc_hd__xor2_4
X_4209_ _4210_/A _4210_/B _4210_/C vssd1 vssd1 vccd1 vccd1 _4209_/X sky130_fd_sc_hd__and3_4
X_5189_ _5189_/A _5189_/B _5248_/A vssd1 vssd1 vccd1 vccd1 _5722_/B sky130_fd_sc_hd__or3_4
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout180 _7558_/X vssd1 vssd1 vccd1 vccd1 _7918_/B sky130_fd_sc_hd__buf_4
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout191 _4219_/Y vssd1 vssd1 vccd1 vccd1 _4548_/B sky130_fd_sc_hd__buf_6
XFILLER_14_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4560_ _7116_/A _4630_/B _4630_/C vssd1 vssd1 vccd1 vccd1 _4561_/C sky130_fd_sc_hd__o21ai_4
XFILLER_116_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4491_ _4360_/A _4487_/X _4490_/X _4570_/A vssd1 vssd1 vccd1 vccd1 _4642_/B sky130_fd_sc_hd__a31oi_4
X_6230_ _5847_/Y _6228_/X _6229_/Y vssd1 vssd1 vccd1 vccd1 _6231_/A sky130_fd_sc_hd__o21a_2
XFILLER_97_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6161_ _6778_/B _6174_/A _6156_/A _6177_/B _6160_/X vssd1 vssd1 vccd1 vccd1 _6161_/Y
+ sky130_fd_sc_hd__a221oi_4
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5112_ _5113_/A _5113_/B vssd1 vssd1 vccd1 vccd1 _5155_/B sky130_fd_sc_hd__or2_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6092_ _6092_/A _6092_/B vssd1 vssd1 vccd1 vccd1 _6132_/B sky130_fd_sc_hd__xnor2_4
XFILLER_69_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5043_/A _5043_/B vssd1 vssd1 vccd1 vccd1 _5043_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_65_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6994_ _6994_/A _6994_/B vssd1 vssd1 vccd1 vccd1 _6995_/B sky130_fd_sc_hd__or2_2
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5945_ _5615_/Y _5940_/X _5944_/Y _5946_/B vssd1 vssd1 vccd1 vccd1 _6144_/B sky130_fd_sc_hd__a31oi_4
XFILLER_25_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5876_ _5874_/Y _5876_/B vssd1 vssd1 vccd1 vccd1 _6241_/A sky130_fd_sc_hd__nand2b_2
X_7615_ _7648_/A _7648_/B vssd1 vssd1 vccd1 vccd1 _7622_/B sky130_fd_sc_hd__and2_1
X_4827_ _4832_/A _4832_/B vssd1 vssd1 vccd1 vccd1 _4833_/A sky130_fd_sc_hd__nor2_2
XFILLER_21_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7546_ _7889_/A _7537_/D _7545_/X _7544_/X vssd1 vssd1 vccd1 vccd1 _7546_/X sky130_fd_sc_hd__o31a_1
X_4758_ _4746_/A _4757_/B _4757_/Y vssd1 vssd1 vccd1 vccd1 _4759_/B sky130_fd_sc_hd__o21ai_1
XFILLER_107_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7477_ _7477_/A _7477_/B vssd1 vssd1 vccd1 vccd1 _7477_/X sky130_fd_sc_hd__xor2_2
X_4689_ _4689_/A _4689_/B _4689_/C vssd1 vssd1 vccd1 vccd1 _4712_/A sky130_fd_sc_hd__and3_2
X_6428_ _6475_/A _6429_/B vssd1 vssd1 vccd1 vccd1 _6476_/A sky130_fd_sc_hd__nand2_2
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6359_ _6359_/A _6492_/B vssd1 vssd1 vccd1 vccd1 _6451_/A sky130_fd_sc_hd__nand2_4
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8029_ _8065_/CLK _8029_/D vssd1 vssd1 vccd1 vccd1 _8029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5730_ _5730_/A _5730_/B vssd1 vssd1 vccd1 vccd1 _5732_/B sky130_fd_sc_hd__xnor2_4
XFILLER_22_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7400_ _7400_/A _7400_/B vssd1 vssd1 vccd1 vccd1 _7403_/B sky130_fd_sc_hd__xnor2_2
X_5661_ _5708_/B _5708_/A vssd1 vssd1 vccd1 vccd1 _5943_/B sky130_fd_sc_hd__and2b_4
X_5592_ _5621_/A _5853_/B vssd1 vssd1 vccd1 vccd1 _5692_/A sky130_fd_sc_hd__or2_4
X_4612_ _4611_/B _4611_/C _4611_/A vssd1 vssd1 vccd1 vccd1 _4614_/B sky130_fd_sc_hd__a21boi_4
X_4543_ _4543_/A _4543_/B vssd1 vssd1 vccd1 vccd1 _4544_/B sky130_fd_sc_hd__xnor2_4
X_7331_ _7366_/A _7247_/D _7358_/B _7334_/A vssd1 vssd1 vccd1 vccd1 _7332_/B sky130_fd_sc_hd__o22a_1
XFILLER_7_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7262_ _7262_/A _7262_/B vssd1 vssd1 vccd1 vccd1 _7276_/A sky130_fd_sc_hd__xnor2_4
X_6213_ _6081_/Y _6111_/B _6111_/C _6012_/B vssd1 vssd1 vccd1 vccd1 _6213_/X sky130_fd_sc_hd__a31o_1
X_4474_ _4377_/A _4551_/A _4472_/Y _4473_/X _4411_/A vssd1 vssd1 vccd1 vccd1 _4474_/X
+ sky130_fd_sc_hd__o221a_1
X_7193_ _7190_/A _7190_/B _7192_/Y vssd1 vssd1 vccd1 vccd1 _7194_/B sky130_fd_sc_hd__a21oi_4
X_6144_ _6144_/A _6144_/B vssd1 vssd1 vccd1 vccd1 _6145_/B sky130_fd_sc_hd__and2_1
XFILLER_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6075_ _6084_/A _6045_/X _6069_/Y _6073_/X vssd1 vssd1 vccd1 vccd1 _6077_/B sky130_fd_sc_hd__a31o_4
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5026_ _5027_/B _5027_/A vssd1 vssd1 vccd1 vccd1 _5026_/X sky130_fd_sc_hd__and2b_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6977_ _6977_/A _6977_/B vssd1 vssd1 vccd1 vccd1 _6994_/A sky130_fd_sc_hd__xor2_4
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5928_ _5928_/A _5928_/B vssd1 vssd1 vccd1 vccd1 _5928_/X sky130_fd_sc_hd__and2_1
XFILLER_41_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5859_ _5859_/A _5881_/D vssd1 vssd1 vccd1 vccd1 _5925_/B sky130_fd_sc_hd__nor2_1
XFILLER_107_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7529_ _7535_/A _7529_/B vssd1 vssd1 vccd1 vccd1 _7529_/X sky130_fd_sc_hd__or2_1
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4190_ _4192_/B vssd1 vssd1 vccd1 vccd1 _4190_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7880_ _7863_/X _7878_/X _7879_/Y _7991_/D vssd1 vssd1 vccd1 vccd1 _7880_/X sky130_fd_sc_hd__a2bb2o_1
X_6900_ _6943_/A _6943_/B vssd1 vssd1 vccd1 vccd1 _6900_/X sky130_fd_sc_hd__or2_1
XFILLER_90_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6831_ _6831_/A _6831_/B vssd1 vssd1 vccd1 vccd1 _7454_/A sky130_fd_sc_hd__xor2_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6762_ _6734_/Y _6761_/Y _7581_/S vssd1 vssd1 vccd1 vccd1 _6762_/X sky130_fd_sc_hd__mux2_1
X_6693_ _6685_/Y _6692_/X _6713_/S vssd1 vssd1 vccd1 vccd1 _6693_/X sky130_fd_sc_hd__mux2_1
X_5713_ _5713_/A _5713_/B vssd1 vssd1 vccd1 vccd1 _5720_/A sky130_fd_sc_hd__xnor2_4
X_5644_ _5645_/B _5645_/A vssd1 vssd1 vccd1 vccd1 _5644_/X sky130_fd_sc_hd__and2b_1
XFILLER_31_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7314_ _7316_/A _7316_/B vssd1 vssd1 vccd1 vccd1 _7314_/Y sky130_fd_sc_hd__nand2_1
X_5575_ _5575_/A _5631_/C vssd1 vssd1 vccd1 vccd1 _5576_/B sky130_fd_sc_hd__xnor2_4
XFILLER_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4526_ _7165_/A _4456_/B _4920_/A _4430_/B vssd1 vssd1 vccd1 vccd1 _4528_/A sky130_fd_sc_hd__a22o_1
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7245_ _7245_/A _7371_/B vssd1 vssd1 vccd1 vccd1 _7278_/A sky130_fd_sc_hd__nor2_4
X_4457_ _4457_/A _4503_/A vssd1 vssd1 vccd1 vccd1 _4457_/Y sky130_fd_sc_hd__nor2_1
X_7176_ _7176_/A _7176_/B vssd1 vssd1 vccd1 vccd1 _7204_/A sky130_fd_sc_hd__xor2_4
XFILLER_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6127_ _6127_/A vssd1 vssd1 vccd1 vccd1 _6156_/A sky130_fd_sc_hd__clkinv_4
XFILLER_58_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4388_ _7165_/A _5019_/A vssd1 vssd1 vccd1 vccd1 _4393_/A sky130_fd_sc_hd__nand2_4
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6058_ _6058_/A _6058_/B vssd1 vssd1 vccd1 vccd1 _6059_/B sky130_fd_sc_hd__and2_1
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5009_ _5009_/A _5009_/B vssd1 vssd1 vccd1 vccd1 _5299_/A sky130_fd_sc_hd__xnor2_1
XFILLER_39_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5360_ _5360_/A _5360_/B vssd1 vssd1 vccd1 vccd1 _5551_/A sky130_fd_sc_hd__xor2_4
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4311_ _4200_/B _5989_/B _4263_/X _4548_/B vssd1 vssd1 vccd1 vccd1 _4312_/C sky130_fd_sc_hd__o211ai_4
X_5291_ _5367_/A _5344_/B vssd1 vssd1 vccd1 vccd1 _5298_/A sky130_fd_sc_hd__nor2_8
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4242_ _4242_/A _5989_/B vssd1 vssd1 vccd1 vccd1 _4242_/X sky130_fd_sc_hd__or2_1
XFILLER_4_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7030_ _7030_/A _7294_/B vssd1 vssd1 vccd1 vccd1 _7079_/A sky130_fd_sc_hd__nor2_2
X_4173_ _4228_/A _4172_/B _4170_/X vssd1 vssd1 vccd1 vccd1 _4174_/B sky130_fd_sc_hd__a21oi_4
XFILLER_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7932_ _7911_/B _7929_/X _7931_/X vssd1 vssd1 vccd1 vccd1 _7934_/A sky130_fd_sc_hd__a21oi_1
XFILLER_95_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7863_ _7887_/A _7860_/Y _7887_/B _7862_/Y _6268_/X vssd1 vssd1 vccd1 vccd1 _7863_/X
+ sky130_fd_sc_hd__o311a_2
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7794_ _7793_/A _7793_/B _6774_/X vssd1 vssd1 vccd1 vccd1 _7794_/X sky130_fd_sc_hd__a21o_1
X_6814_ _6804_/A _6804_/B _6815_/B vssd1 vssd1 vccd1 vccd1 _6824_/A sky130_fd_sc_hd__a21o_1
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6745_ _6707_/B _6708_/X _7581_/S vssd1 vssd1 vccd1 vccd1 _6745_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6676_ _6539_/B _6538_/A _6737_/B vssd1 vssd1 vccd1 vccd1 _6677_/A sky130_fd_sc_hd__mux2_1
X_5627_ _5627_/A _5627_/B vssd1 vssd1 vccd1 vccd1 _5679_/A sky130_fd_sc_hd__xnor2_4
X_5558_ _5558_/A _5608_/A _5558_/C vssd1 vssd1 vccd1 vccd1 _5559_/B sky130_fd_sc_hd__nand3_1
XFILLER_105_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4509_ _4509_/A _4509_/B vssd1 vssd1 vccd1 vccd1 _4511_/B sky130_fd_sc_hd__xnor2_4
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5489_ _5490_/A _5490_/B vssd1 vssd1 vccd1 vccd1 _5497_/A sky130_fd_sc_hd__nor2_2
X_7228_ _7228_/A _7228_/B vssd1 vssd1 vccd1 vccd1 _7241_/A sky130_fd_sc_hd__xnor2_4
XFILLER_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7159_ _7159_/A _7159_/B vssd1 vssd1 vccd1 vccd1 _7160_/B sky130_fd_sc_hd__or2_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _4860_/A _4860_/B _4860_/C vssd1 vssd1 vccd1 vccd1 _4860_/Y sky130_fd_sc_hd__nor3_1
XFILLER_17_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6530_ _6539_/A _6539_/B vssd1 vssd1 vccd1 vccd1 _6530_/Y sky130_fd_sc_hd__nor2_1
X_4791_ _4775_/A _4775_/B _4800_/A _4775_/D vssd1 vssd1 vccd1 vccd1 _4792_/B sky130_fd_sc_hd__a22o_1
X_6461_ _6476_/A _6460_/A _6476_/B vssd1 vssd1 vccd1 vccd1 _6531_/B sky130_fd_sc_hd__a21boi_2
X_6392_ _6354_/X _6391_/Y _6441_/S vssd1 vssd1 vccd1 vccd1 _6394_/B sky130_fd_sc_hd__mux2_4
X_5412_ _5412_/A _5412_/B vssd1 vssd1 vccd1 vccd1 _5414_/B sky130_fd_sc_hd__xnor2_4
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5343_ _5343_/A _5343_/B vssd1 vssd1 vccd1 vccd1 _5346_/A sky130_fd_sc_hd__xor2_4
XFILLER_114_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8062_ _8063_/CLK _8062_/D vssd1 vssd1 vccd1 vccd1 _8062_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5274_ _5445_/A _6871_/C vssd1 vssd1 vccd1 vccd1 _5275_/C sky130_fd_sc_hd__nor2_4
XFILLER_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4225_ _4192_/X _4195_/X _4200_/Y _4193_/A vssd1 vssd1 vccd1 vccd1 _4225_/X sky130_fd_sc_hd__a31o_1
X_7013_ _7013_/A _7013_/B _7013_/C vssd1 vssd1 vccd1 vccd1 _7071_/A sky130_fd_sc_hd__and3_1
X_4156_ _8078_/Q _4156_/B vssd1 vssd1 vccd1 vccd1 _4242_/A sky130_fd_sc_hd__xnor2_4
XFILLER_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4087_ _4087_/A _4087_/B vssd1 vssd1 vccd1 vccd1 _4087_/X sky130_fd_sc_hd__xor2_1
XFILLER_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7915_ _7877_/B _7891_/Y _7939_/A vssd1 vssd1 vccd1 vccd1 _7917_/B sky130_fd_sc_hd__o21ai_1
XFILLER_70_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7846_ _7874_/A _7874_/B _7874_/C _7837_/A vssd1 vssd1 vccd1 vccd1 _7846_/X sky130_fd_sc_hd__o31a_1
XFILLER_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7777_ _7777_/A _7777_/B vssd1 vssd1 vccd1 vccd1 _7777_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4989_ _4989_/A _5033_/B vssd1 vssd1 vccd1 vccd1 _5022_/A sky130_fd_sc_hd__or2_4
X_6728_ _6713_/X _6721_/X _6733_/S vssd1 vssd1 vccd1 vccd1 _6728_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6659_ _6689_/S _6659_/B vssd1 vssd1 vccd1 vccd1 _6659_/X sky130_fd_sc_hd__and2b_1
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4010_ _8048_/Q _8047_/Q _8046_/Q vssd1 vssd1 vccd1 vccd1 _7956_/C sky130_fd_sc_hd__or3_2
XFILLER_96_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5961_ _5961_/A _5961_/B vssd1 vssd1 vccd1 vccd1 _6180_/C sky130_fd_sc_hd__xnor2_2
XFILLER_18_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7700_ _7784_/A _6255_/C _7699_/Y vssd1 vssd1 vccd1 vccd1 _7703_/B sky130_fd_sc_hd__o21ai_4
XFILLER_52_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4912_ _4914_/A _4914_/B _4914_/C vssd1 vssd1 vccd1 vccd1 _4915_/A sky130_fd_sc_hd__a21oi_2
X_7631_ _7929_/A _7656_/A _7656_/B vssd1 vssd1 vccd1 vccd1 _7632_/B sky130_fd_sc_hd__o21a_1
X_5892_ _5893_/A _5893_/B _5901_/A vssd1 vssd1 vccd1 vccd1 _5896_/A sky130_fd_sc_hd__and3_1
X_4843_ _4929_/A _5020_/B vssd1 vssd1 vccd1 vccd1 _4930_/A sky130_fd_sc_hd__nor2_1
X_7562_ _7964_/C _7562_/B vssd1 vssd1 vccd1 vccd1 _7562_/X sky130_fd_sc_hd__and2b_1
X_4774_ _4947_/A _4795_/C _4820_/S vssd1 vssd1 vccd1 vccd1 _4775_/D sky130_fd_sc_hd__a21bo_2
X_6513_ _7728_/A _6469_/Y _6512_/X vssd1 vssd1 vccd1 vccd1 _6514_/B sky130_fd_sc_hd__o21bai_2
X_7493_ _7444_/X _7480_/X _7515_/S vssd1 vssd1 vccd1 vccd1 _7493_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6444_ _6444_/A _6444_/B vssd1 vssd1 vccd1 vccd1 _6447_/A sky130_fd_sc_hd__nand2_1
X_6375_ _6374_/A _6374_/B _6374_/C vssd1 vssd1 vccd1 vccd1 _6376_/A sky130_fd_sc_hd__o21a_1
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5326_ _5530_/A _7358_/B _5534_/B _5321_/X vssd1 vssd1 vccd1 vccd1 _5336_/A sky130_fd_sc_hd__o31a_4
XFILLER_114_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8045_ _8057_/CLK _8045_/D vssd1 vssd1 vccd1 vccd1 _8045_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5257_ _5257_/A _5257_/B vssd1 vssd1 vccd1 vccd1 _5258_/B sky130_fd_sc_hd__xor2_4
X_4208_ _4184_/Y _4206_/X _4210_/A vssd1 vssd1 vccd1 vccd1 _4208_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_96_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5188_ _5189_/B _5248_/A _5189_/A vssd1 vssd1 vccd1 vccd1 _5722_/A sky130_fd_sc_hd__o21ai_4
XFILLER_29_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4139_ _7170_/B _4138_/X _5986_/S vssd1 vssd1 vccd1 vccd1 _6007_/A sky130_fd_sc_hd__mux2_8
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7829_ _7562_/B _7827_/Y _7828_/X vssd1 vssd1 vccd1 vccd1 _7830_/B sky130_fd_sc_hd__o21ba_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout181 _7558_/X vssd1 vssd1 vccd1 vccd1 _7802_/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout192 _4208_/Y vssd1 vssd1 vccd1 vccd1 _4341_/A1 sky130_fd_sc_hd__buf_8
Xfanout170 _4080_/X vssd1 vssd1 vccd1 vccd1 _5322_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_19_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_4__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _8080_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4490_ _4377_/A _4489_/X _4488_/X _4411_/A vssd1 vssd1 vccd1 vccd1 _4490_/X sky130_fd_sc_hd__a211o_2
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6160_ _6177_/A _6160_/B vssd1 vssd1 vccd1 vccd1 _6160_/X sky130_fd_sc_hd__and2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5111_ _5174_/A _5111_/B vssd1 vssd1 vccd1 vccd1 _5113_/B sky130_fd_sc_hd__xnor2_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6091_ _6091_/A _6091_/B vssd1 vssd1 vccd1 vccd1 _6092_/B sky130_fd_sc_hd__xnor2_4
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5039_/A _5039_/B _5041_/X vssd1 vssd1 vccd1 vccd1 _5042_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6993_ _6993_/A _6993_/B vssd1 vssd1 vccd1 vccd1 _7045_/A sky130_fd_sc_hd__xnor2_2
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5944_ _6135_/B _6115_/A vssd1 vssd1 vccd1 vccd1 _5944_/Y sky130_fd_sc_hd__nor2_2
X_5875_ _5875_/A _5875_/B vssd1 vssd1 vccd1 vccd1 _5876_/B sky130_fd_sc_hd__nand2_1
X_7614_ _7607_/X _7612_/X _7613_/Y vssd1 vssd1 vccd1 vccd1 _7614_/Y sky130_fd_sc_hd__a21oi_2
X_4826_ _4826_/A _4826_/B vssd1 vssd1 vccd1 vccd1 _4832_/B sky130_fd_sc_hd__xnor2_1
X_7545_ _7527_/S _7523_/X _7525_/Y _7515_/X _7535_/A vssd1 vssd1 vccd1 vccd1 _7545_/X
+ sky130_fd_sc_hd__a32o_1
X_4757_ _5090_/A _4757_/B vssd1 vssd1 vccd1 vccd1 _4757_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7476_ _7473_/X _7475_/X _7527_/S vssd1 vssd1 vccd1 vccd1 _7476_/X sky130_fd_sc_hd__mux2_1
X_4688_ _4687_/A _4727_/A _4687_/B vssd1 vssd1 vccd1 vccd1 _4689_/C sky130_fd_sc_hd__o21a_1
X_6427_ _6475_/B vssd1 vssd1 vccd1 vccd1 _6429_/B sky130_fd_sc_hd__inv_2
XFILLER_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6358_ _6359_/A _6492_/B vssd1 vssd1 vccd1 vccd1 _6484_/S sky130_fd_sc_hd__and2_4
XFILLER_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5309_ _5294_/A _5518_/A _5307_/X vssd1 vssd1 vccd1 vccd1 _5311_/A sky130_fd_sc_hd__o21ba_2
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6289_ _6289_/A _6289_/B vssd1 vssd1 vccd1 vccd1 _6289_/X sky130_fd_sc_hd__or2_1
XFILLER_102_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8028_ _8065_/CLK _8028_/D vssd1 vssd1 vccd1 vccd1 _8028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5660_ _5660_/A _5660_/B vssd1 vssd1 vccd1 vccd1 _5708_/B sky130_fd_sc_hd__xor2_2
XFILLER_30_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4611_ _4611_/A _4611_/B _4611_/C vssd1 vssd1 vccd1 vccd1 _4611_/X sky130_fd_sc_hd__and3_2
X_5591_ _5600_/A _5600_/B vssd1 vssd1 vccd1 vccd1 _5591_/Y sky130_fd_sc_hd__nand2b_1
X_7330_ _7330_/A _7330_/B vssd1 vssd1 vccd1 vccd1 _7340_/A sky130_fd_sc_hd__xnor2_4
X_4542_ _4519_/A _4519_/B _4512_/Y vssd1 vssd1 vccd1 vccd1 _4543_/B sky130_fd_sc_hd__o21a_2
XFILLER_116_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4473_ _4472_/A _4419_/X _6878_/C vssd1 vssd1 vccd1 vccd1 _4473_/X sky130_fd_sc_hd__a21o_1
X_7261_ _7261_/A _7371_/B _7262_/B vssd1 vssd1 vccd1 vccd1 _7275_/A sky130_fd_sc_hd__or3_4
XFILLER_89_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6212_ _6254_/S _6199_/X _6209_/X _6166_/S vssd1 vssd1 vccd1 vccd1 _6212_/X sky130_fd_sc_hd__a211o_1
X_7192_ _7202_/A _7202_/B vssd1 vssd1 vccd1 vccd1 _7192_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6143_ _6144_/A _6144_/B vssd1 vssd1 vccd1 vccd1 _6147_/B sky130_fd_sc_hd__nor2_2
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6074_ _6084_/A _6045_/X _6069_/Y _6073_/X vssd1 vssd1 vccd1 vccd1 _6078_/C sky130_fd_sc_hd__a31oi_4
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _5043_/A _5024_/B _5018_/X vssd1 vssd1 vccd1 vccd1 _5027_/B sky130_fd_sc_hd__a21oi_4
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6976_ _7030_/A _7247_/C _7021_/B _6973_/Y vssd1 vssd1 vccd1 vccd1 _6977_/B sky130_fd_sc_hd__o31ai_4
XFILLER_80_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5927_ _7085_/B _5927_/B _5927_/C _5927_/D vssd1 vssd1 vccd1 vccd1 _5928_/B sky130_fd_sc_hd__and4_1
X_5858_ _7285_/B _5858_/B vssd1 vssd1 vccd1 vccd1 _5881_/D sky130_fd_sc_hd__nand2_1
X_4809_ _4809_/A _4809_/B vssd1 vssd1 vccd1 vccd1 _4815_/B sky130_fd_sc_hd__xor2_2
X_5789_ _5762_/A _5761_/C _5761_/A vssd1 vssd1 vccd1 vccd1 _5794_/B sky130_fd_sc_hd__a21o_1
X_7528_ _7527_/S _7513_/X _7523_/X vssd1 vssd1 vccd1 vccd1 _7529_/B sky130_fd_sc_hd__a21o_1
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7459_ _7459_/A vssd1 vssd1 vccd1 vccd1 _7459_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6830_ _7392_/C _6830_/B vssd1 vssd1 vccd1 vccd1 _6831_/B sky130_fd_sc_hd__nor2_1
XFILLER_63_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6761_ _6608_/X _6616_/B _6610_/A vssd1 vssd1 vccd1 vccd1 _6761_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5712_ _5615_/Y _5710_/X _5711_/Y vssd1 vssd1 vccd1 vccd1 _5946_/B sky130_fd_sc_hd__a21o_2
X_6692_ _6697_/S _6691_/Y _6690_/X vssd1 vssd1 vccd1 vccd1 _6692_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5643_ _5643_/A _5643_/B vssd1 vssd1 vccd1 vccd1 _5645_/B sky130_fd_sc_hd__xnor2_4
XFILLER_117_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5574_ _5574_/A _5632_/A vssd1 vssd1 vccd1 vccd1 _5574_/Y sky130_fd_sc_hd__nor2_1
X_7313_ _7330_/A _7330_/B vssd1 vssd1 vccd1 vccd1 _7316_/B sky130_fd_sc_hd__and2b_2
X_4525_ _7085_/A _4551_/B vssd1 vssd1 vccd1 vccd1 _4529_/A sky130_fd_sc_hd__nand2_2
X_7244_ _7244_/A _7244_/B vssd1 vssd1 vccd1 vccd1 _7257_/A sky130_fd_sc_hd__xnor2_4
X_4456_ _7319_/A _4456_/B vssd1 vssd1 vccd1 vccd1 _4503_/A sky130_fd_sc_hd__nand2_8
X_4387_ _4387_/A _4555_/A vssd1 vssd1 vccd1 vccd1 _4395_/A sky130_fd_sc_hd__nand2_4
X_7175_ _7176_/A _7176_/B vssd1 vssd1 vccd1 vccd1 _7184_/B sky130_fd_sc_hd__nand2b_1
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6126_ _6242_/S _6174_/A vssd1 vssd1 vccd1 vccd1 _6127_/A sky130_fd_sc_hd__or2_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _6058_/A _6058_/B vssd1 vssd1 vccd1 vccd1 _6059_/A sky130_fd_sc_hd__nor2_1
XFILLER_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5008_ _5008_/A _5008_/B vssd1 vssd1 vccd1 vccd1 _5703_/A sky130_fd_sc_hd__xnor2_4
XFILLER_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6959_ _5745_/A _6999_/A _7114_/C _6943_/X vssd1 vssd1 vccd1 vccd1 _6960_/B sky130_fd_sc_hd__a31o_1
XFILLER_41_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4310_ _4187_/B _4259_/B _4270_/X _4548_/B vssd1 vssd1 vccd1 vccd1 _4312_/B sky130_fd_sc_hd__a211o_2
X_5290_ _5290_/A _5290_/B vssd1 vssd1 vccd1 vccd1 _5344_/B sky130_fd_sc_hd__xnor2_4
XFILLER_114_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4241_ _4241_/A _4241_/B vssd1 vssd1 vccd1 vccd1 _4241_/X sky130_fd_sc_hd__or2_1
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4172_ _4228_/A _4172_/B vssd1 vssd1 vccd1 vccd1 _4172_/X sky130_fd_sc_hd__and2_1
XFILLER_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7931_ _7729_/X _7930_/Y _7908_/A vssd1 vssd1 vccd1 vccd1 _7931_/X sky130_fd_sc_hd__a21o_1
XFILLER_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7862_ _7887_/A _7887_/B _7860_/Y vssd1 vssd1 vccd1 vccd1 _7862_/Y sky130_fd_sc_hd__o21ai_1
X_7793_ _7793_/A _7793_/B vssd1 vssd1 vccd1 vccd1 _7793_/Y sky130_fd_sc_hd__nor2_4
X_6813_ _6827_/B _6813_/B vssd1 vssd1 vccd1 vccd1 _6815_/B sky130_fd_sc_hd__nand2_1
X_6744_ _6757_/B vssd1 vssd1 vccd1 vccd1 _6744_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6675_ _6753_/S _6675_/B vssd1 vssd1 vccd1 vccd1 _6675_/X sky130_fd_sc_hd__and2_1
XFILLER_50_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5626_ _5627_/A _5627_/B vssd1 vssd1 vccd1 vccd1 _5626_/X sky130_fd_sc_hd__and2b_1
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5557_ _5558_/A _5608_/A _5558_/C vssd1 vssd1 vccd1 vccd1 _5614_/A sky130_fd_sc_hd__a21o_2
XFILLER_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5488_ _5474_/A _5474_/B _5472_/X vssd1 vssd1 vccd1 vccd1 _5490_/B sky130_fd_sc_hd__a21oi_4
X_4508_ _4508_/A _4508_/B vssd1 vssd1 vccd1 vccd1 _4509_/B sky130_fd_sc_hd__xnor2_4
XFILLER_105_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7227_ _7227_/A _7228_/A _7227_/C vssd1 vssd1 vccd1 vccd1 _7240_/A sky130_fd_sc_hd__and3_4
X_4439_ _4602_/A _4359_/Y _4405_/Y _4379_/Y vssd1 vssd1 vccd1 vccd1 _4439_/X sky130_fd_sc_hd__a31o_1
XFILLER_59_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7158_ _7158_/A _7158_/B vssd1 vssd1 vccd1 vccd1 _7190_/A sky130_fd_sc_hd__xnor2_4
XFILLER_86_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6109_ _6111_/B _6111_/C vssd1 vssd1 vccd1 vccd1 _6134_/A sky130_fd_sc_hd__nand2_4
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7089_ _4329_/X _7247_/D _7141_/A _7087_/B _7087_/A vssd1 vssd1 vccd1 vccd1 _7090_/B
+ sky130_fd_sc_hd__o32a_4
XFILLER_100_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4790_ _4854_/A _4790_/B vssd1 vssd1 vccd1 vccd1 _4809_/A sky130_fd_sc_hd__xnor2_2
XFILLER_60_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6460_ _6460_/A vssd1 vssd1 vccd1 vccd1 _6460_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6391_ _6451_/A _6369_/Y _6390_/Y vssd1 vssd1 vccd1 vccd1 _6391_/Y sky130_fd_sc_hd__a21oi_2
X_5411_ _5411_/A _5411_/B vssd1 vssd1 vccd1 vccd1 _5412_/B sky130_fd_sc_hd__xor2_4
XFILLER_114_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5342_ _6842_/B _5342_/B vssd1 vssd1 vccd1 vccd1 _5343_/B sky130_fd_sc_hd__nor2_4
X_8061_ _8063_/CLK _8061_/D vssd1 vssd1 vccd1 vccd1 _8061_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_114_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7012_ _7012_/A _7294_/B vssd1 vssd1 vccd1 vccd1 _7013_/C sky130_fd_sc_hd__nor2_1
X_5273_ _5273_/A _7247_/D vssd1 vssd1 vccd1 vccd1 _5446_/B sky130_fd_sc_hd__or2_4
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4224_ _4192_/X _4195_/X _4200_/Y _4193_/A vssd1 vssd1 vccd1 vccd1 _4224_/Y sky130_fd_sc_hd__a31oi_1
X_4155_ _4175_/B _4147_/B _4144_/X _4211_/B vssd1 vssd1 vccd1 vccd1 _4156_/B sky130_fd_sc_hd__o31a_2
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4086_ _8052_/Q _4086_/B vssd1 vssd1 vccd1 vccd1 _4087_/B sky130_fd_sc_hd__xnor2_4
X_7914_ _7914_/A _7914_/B vssd1 vssd1 vccd1 vccd1 _7917_/A sky130_fd_sc_hd__xor2_2
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7845_ _7844_/A _7844_/B _7923_/A vssd1 vssd1 vccd1 vccd1 _7845_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7776_ _7789_/A _7789_/B vssd1 vssd1 vccd1 vccd1 _7777_/B sky130_fd_sc_hd__nor2_1
X_4988_ _4988_/A _5033_/B vssd1 vssd1 vccd1 vccd1 _4990_/B sky130_fd_sc_hd__nor2_2
X_6727_ _6675_/B _6687_/X _6753_/S vssd1 vssd1 vccd1 vccd1 _6727_/X sky130_fd_sc_hd__mux2_1
X_6658_ _6534_/Y _6537_/Y _6688_/S vssd1 vssd1 vccd1 vccd1 _6659_/B sky130_fd_sc_hd__mux2_1
X_5609_ _5616_/A _5616_/B _5616_/C vssd1 vssd1 vccd1 vccd1 _5617_/A sky130_fd_sc_hd__a21oi_4
X_6589_ _6590_/A _6590_/B vssd1 vssd1 vccd1 vccd1 _6592_/B sky130_fd_sc_hd__and2b_2
XFILLER_105_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5960_ _5960_/A _5960_/B vssd1 vssd1 vccd1 vccd1 _5961_/B sky130_fd_sc_hd__nand2_2
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4911_ _4911_/A _4911_/B vssd1 vssd1 vccd1 vccd1 _4914_/C sky130_fd_sc_hd__xnor2_1
XFILLER_33_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5891_ _5900_/A _5900_/B vssd1 vssd1 vccd1 vccd1 _5901_/A sky130_fd_sc_hd__nor2_1
X_7630_ _7687_/A _7630_/B vssd1 vssd1 vccd1 vccd1 _7656_/B sky130_fd_sc_hd__or2_1
X_4842_ _4730_/Y _4841_/X _4840_/X vssd1 vssd1 vccd1 vccd1 _4842_/X sky130_fd_sc_hd__a21bo_1
XFILLER_20_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7561_ _7557_/Y _7918_/B _7559_/X _7560_/X vssd1 vssd1 vccd1 vccd1 _7561_/X sky130_fd_sc_hd__o31a_1
X_4773_ _4773_/A _5013_/A _5014_/A _4795_/C vssd1 vssd1 vccd1 vccd1 _4800_/A sky130_fd_sc_hd__or4_4
X_6512_ _6517_/A _6510_/Y _6511_/X _7728_/A vssd1 vssd1 vccd1 vccd1 _6512_/X sky130_fd_sc_hd__o211a_1
X_7492_ _7476_/X _7491_/X _7515_/S vssd1 vssd1 vccd1 vccd1 _7531_/B sky130_fd_sc_hd__mux2_1
XFILLER_107_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6443_ _6443_/A _6443_/B vssd1 vssd1 vccd1 vccd1 _6444_/B sky130_fd_sc_hd__or2_1
X_6374_ _6374_/A _6374_/B _6374_/C vssd1 vssd1 vccd1 vccd1 _6377_/A sky130_fd_sc_hd__or3_2
X_5325_ _5325_/A _5325_/B vssd1 vssd1 vccd1 vccd1 _5534_/B sky130_fd_sc_hd__xnor2_4
XFILLER_114_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8044_ _8082_/CLK _8044_/D vssd1 vssd1 vccd1 vccd1 _8044_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_88_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5256_ _5257_/A _5257_/B vssd1 vssd1 vccd1 vccd1 _5256_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4207_ _4184_/Y _4206_/X _4210_/A vssd1 vssd1 vccd1 vccd1 _4207_/X sky130_fd_sc_hd__o21a_1
X_5187_ _5187_/A _5187_/B vssd1 vssd1 vccd1 vccd1 _5196_/A sky130_fd_sc_hd__xnor2_4
X_4138_ _5066_/B _4137_/X _5087_/B vssd1 vssd1 vccd1 vccd1 _4138_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4069_ _4071_/B vssd1 vssd1 vccd1 vccd1 _6273_/A sky130_fd_sc_hd__inv_2
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7828_ _8036_/Q _4018_/X _7944_/B _8037_/Q vssd1 vssd1 vccd1 vccd1 _7828_/X sky130_fd_sc_hd__a22o_1
X_7759_ _7833_/A _7759_/B vssd1 vssd1 vccd1 vccd1 _7759_/Y sky130_fd_sc_hd__nor2_2
XFILLER_12_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout171 _4080_/X vssd1 vssd1 vccd1 vccd1 _5977_/A sky130_fd_sc_hd__buf_4
Xfanout182 _4547_/C vssd1 vssd1 vccd1 vccd1 _4356_/A sky130_fd_sc_hd__buf_6
Xfanout160 _4329_/X vssd1 vssd1 vccd1 vccd1 _7030_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_47_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout193 _4208_/Y vssd1 vssd1 vccd1 vccd1 _6034_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6090_ _6084_/A _6088_/B _6026_/X vssd1 vssd1 vccd1 vccd1 _6091_/B sky130_fd_sc_hd__a21boi_4
X_5110_ _5110_/A _5156_/C vssd1 vssd1 vccd1 vccd1 _5155_/A sky130_fd_sc_hd__or2_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _4984_/B _5040_/Y _5034_/C _5034_/A _5041_/D1 vssd1 vssd1 vccd1 vccd1 _5041_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_111_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6992_ _6992_/A _6992_/B vssd1 vssd1 vccd1 vccd1 _7048_/A sky130_fd_sc_hd__nand2_1
XFILLER_80_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5943_ _5943_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _6115_/A sky130_fd_sc_hd__xnor2_4
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5874_ _5875_/A _5875_/B vssd1 vssd1 vccd1 vccd1 _5874_/Y sky130_fd_sc_hd__nor2_1
X_7613_ _7607_/X _7612_/X _6268_/X vssd1 vssd1 vccd1 vccd1 _7613_/Y sky130_fd_sc_hd__o21ai_1
X_4825_ _4826_/A _4826_/B vssd1 vssd1 vccd1 vccd1 _4829_/B sky130_fd_sc_hd__and2_2
X_7544_ _7544_/A _7544_/B _7544_/C _7544_/D vssd1 vssd1 vccd1 vccd1 _7544_/X sky130_fd_sc_hd__or4_1
XFILLER_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4756_ _5020_/A _4751_/C _5090_/B _4991_/A vssd1 vssd1 vccd1 vccd1 _4761_/A sky130_fd_sc_hd__a22o_1
XFILLER_107_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7475_ _7472_/X _7474_/X _7513_/S vssd1 vssd1 vccd1 vccd1 _7475_/X sky130_fd_sc_hd__mux2_1
X_4687_ _4687_/A _4687_/B vssd1 vssd1 vccd1 vccd1 _4720_/A sky130_fd_sc_hd__nand2_1
X_6426_ _6902_/A _7247_/D _6445_/S vssd1 vssd1 vccd1 vccd1 _6475_/B sky130_fd_sc_hd__mux2_4
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6357_ _6386_/A _6359_/A vssd1 vssd1 vccd1 vccd1 _6488_/B sky130_fd_sc_hd__nand2_2
X_5308_ _6873_/B _5723_/A vssd1 vssd1 vccd1 vccd1 _5518_/A sky130_fd_sc_hd__nand2_8
X_6288_ _4077_/B _4242_/A _4172_/B _4059_/B vssd1 vssd1 vccd1 vccd1 _6288_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8027_ _8057_/CLK _8027_/D vssd1 vssd1 vccd1 vccd1 _8027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5239_ _5239_/A _5239_/B vssd1 vssd1 vccd1 vccd1 _5498_/A sky130_fd_sc_hd__xnor2_4
XFILLER_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4610_ _4574_/X _4607_/Y _4606_/Y _4606_/A vssd1 vssd1 vccd1 vccd1 _4611_/C sky130_fd_sc_hd__a211o_4
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5590_ _5643_/A _5643_/B _5580_/A vssd1 vssd1 vccd1 vccd1 _5600_/B sky130_fd_sc_hd__a21o_2
X_4541_ _7311_/A _4518_/B _4517_/A vssd1 vssd1 vccd1 vccd1 _4543_/A sky130_fd_sc_hd__o21ai_4
XFILLER_116_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4472_ _4472_/A _4472_/B vssd1 vssd1 vccd1 vccd1 _4472_/Y sky130_fd_sc_hd__nor2_1
X_7260_ _7252_/A _7252_/B _7255_/X vssd1 vssd1 vccd1 vccd1 _7262_/B sky130_fd_sc_hd__o21a_2
X_6211_ _7570_/B _6190_/X _6193_/X _6225_/S vssd1 vssd1 vccd1 vccd1 _6211_/X sky130_fd_sc_hd__a211o_1
X_7191_ _7188_/A _7227_/A _7185_/A vssd1 vssd1 vccd1 vccd1 _7202_/B sky130_fd_sc_hd__o21ba_4
X_6142_ _6131_/X _6245_/B _6193_/A vssd1 vssd1 vccd1 vccd1 _6142_/X sky130_fd_sc_hd__mux2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6073_ _6059_/A _6072_/Y _6068_/B vssd1 vssd1 vccd1 vccd1 _6073_/X sky130_fd_sc_hd__o21a_2
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5018_/X _5024_/B vssd1 vssd1 vccd1 vccd1 _5043_/B sky130_fd_sc_hd__and2b_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6975_ _6975_/A _6975_/B vssd1 vssd1 vccd1 vccd1 _7021_/B sky130_fd_sc_hd__xor2_4
XFILLER_53_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5926_ _5881_/A _7210_/B _5821_/B vssd1 vssd1 vccd1 vccd1 _5927_/D sky130_fd_sc_hd__o21ai_1
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5857_ _5857_/A _5857_/B vssd1 vssd1 vccd1 vccd1 _5879_/A sky130_fd_sc_hd__nand2_1
X_4808_ _4809_/B _4809_/A vssd1 vssd1 vccd1 vccd1 _4813_/B sky130_fd_sc_hd__and2b_1
X_5788_ _5788_/A _5788_/B vssd1 vssd1 vccd1 vccd1 _5795_/A sky130_fd_sc_hd__xor2_4
XFILLER_119_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7527_ _7523_/X _7513_/X _7527_/S vssd1 vssd1 vccd1 vccd1 _7527_/X sky130_fd_sc_hd__mux2_1
X_4739_ _5445_/A _4751_/C vssd1 vssd1 vccd1 vccd1 _5090_/B sky130_fd_sc_hd__nor2_8
X_7458_ _7403_/D _7502_/B _7457_/Y vssd1 vssd1 vccd1 vccd1 _7459_/A sky130_fd_sc_hd__o21ai_2
X_6409_ _6400_/X _6408_/X _6431_/S vssd1 vssd1 vccd1 vccd1 _6410_/B sky130_fd_sc_hd__mux2_1
XFILLER_89_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7389_ _6833_/A _6860_/Y _6823_/B vssd1 vssd1 vccd1 vccd1 _7389_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6760_ _6760_/A _6760_/B _7580_/C _6756_/X vssd1 vssd1 vccd1 vccd1 _6760_/X sky130_fd_sc_hd__or4b_1
XFILLER_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5711_ _5614_/A _5610_/Y _5614_/B vssd1 vssd1 vccd1 vccd1 _5711_/Y sky130_fd_sc_hd__a21oi_1
X_6691_ _6691_/A _6691_/B vssd1 vssd1 vccd1 vccd1 _6691_/Y sky130_fd_sc_hd__nor2_2
XFILLER_31_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5642_ _5686_/A _5686_/B _5636_/Y vssd1 vssd1 vccd1 vccd1 _5645_/A sky130_fd_sc_hd__a21bo_4
X_5573_ _5723_/A _7306_/B vssd1 vssd1 vccd1 vccd1 _5632_/A sky130_fd_sc_hd__nand2_4
XFILLER_116_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7312_ _7312_/A _7336_/A vssd1 vssd1 vccd1 vccd1 _7330_/B sky130_fd_sc_hd__xor2_4
X_4524_ _4503_/A _4503_/B _4504_/Y vssd1 vssd1 vccd1 vccd1 _4530_/A sky130_fd_sc_hd__o21a_2
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4455_ _4455_/A _5019_/A vssd1 vssd1 vccd1 vccd1 _4460_/A sky130_fd_sc_hd__nand2_2
X_7243_ _7243_/A _7243_/B vssd1 vssd1 vccd1 vccd1 _7263_/A sky130_fd_sc_hd__or2_4
X_7174_ _7123_/A _7285_/B _7211_/B _7171_/X vssd1 vssd1 vccd1 vccd1 _7176_/B sky130_fd_sc_hd__a31o_4
X_4386_ _7319_/A _4387_/A _4551_/B _4386_/D vssd1 vssd1 vccd1 vccd1 _4555_/A sky130_fd_sc_hd__nand4_4
XFILLER_98_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6125_ _6150_/B _6120_/B _6242_/S vssd1 vssd1 vccd1 vccd1 _6125_/X sky130_fd_sc_hd__mux2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _6058_/B vssd1 vssd1 vccd1 vccd1 _7420_/A sky130_fd_sc_hd__clkinv_4
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5007_ _5008_/A _5008_/B vssd1 vssd1 vccd1 vccd1 _5378_/A sky130_fd_sc_hd__or2_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6958_ _6966_/A _6958_/B vssd1 vssd1 vccd1 vccd1 _6996_/A sky130_fd_sc_hd__and2_1
X_6889_ _6894_/A _6894_/B vssd1 vssd1 vccd1 vccd1 _6895_/A sky130_fd_sc_hd__or2_2
X_5909_ _5909_/A _5918_/A vssd1 vssd1 vccd1 vccd1 _5915_/B sky130_fd_sc_hd__xnor2_1
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4240_ _4241_/A _4241_/B vssd1 vssd1 vccd1 vccd1 _4240_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4171_ _4228_/A _4172_/B _4170_/X vssd1 vssd1 vccd1 vccd1 _4174_/A sky130_fd_sc_hd__o21a_1
X_7930_ _7930_/A _7930_/B vssd1 vssd1 vccd1 vccd1 _7930_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7861_ _7837_/B _7839_/B _7728_/A vssd1 vssd1 vccd1 vccd1 _7887_/B sky130_fd_sc_hd__o21a_1
X_6812_ _6812_/A _6812_/B _6812_/C vssd1 vssd1 vccd1 vccd1 _6813_/B sky130_fd_sc_hd__or3_1
X_7792_ _7741_/A _7741_/B _7777_/Y _7935_/A vssd1 vssd1 vccd1 vccd1 _7793_/B sky130_fd_sc_hd__o31a_2
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6743_ _6727_/X _6742_/X _7616_/S vssd1 vssd1 vccd1 vccd1 _6757_/B sky130_fd_sc_hd__mux2_1
XFILLER_23_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6674_ _6674_/A vssd1 vssd1 vccd1 vccd1 _6675_/B sky130_fd_sc_hd__inv_2
X_5625_ _5566_/B _5666_/B _5663_/A _5663_/B vssd1 vssd1 vccd1 vccd1 _5627_/B sky130_fd_sc_hd__a22o_4
XFILLER_117_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5556_ _5556_/A _5556_/B vssd1 vssd1 vccd1 vccd1 _5558_/C sky130_fd_sc_hd__xnor2_1
X_5487_ _5487_/A _5487_/B vssd1 vssd1 vccd1 vccd1 _5490_/A sky130_fd_sc_hd__xnor2_4
X_4507_ _7136_/A _4630_/B vssd1 vssd1 vccd1 vccd1 _4508_/B sky130_fd_sc_hd__nor2_4
XFILLER_105_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7226_ _7227_/A _7227_/C vssd1 vssd1 vccd1 vccd1 _7228_/B sky130_fd_sc_hd__nand2_2
X_4438_ _4377_/A _5969_/B _4432_/Y _4437_/X _7085_/A vssd1 vssd1 vccd1 vccd1 _4438_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_116_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7157_ _7157_/A _7157_/B vssd1 vssd1 vccd1 vccd1 _7194_/A sky130_fd_sc_hd__xnor2_4
X_4369_ _4441_/A _7214_/A vssd1 vssd1 vccd1 vccd1 _4369_/Y sky130_fd_sc_hd__nand2_1
XFILLER_112_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6108_ _7784_/A vssd1 vssd1 vccd1 vccd1 _7831_/A sky130_fd_sc_hd__clkinv_8
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _7261_/A _7247_/D vssd1 vssd1 vccd1 vccd1 _7141_/B sky130_fd_sc_hd__nor2_2
X_6039_ _6039_/A _6039_/B vssd1 vssd1 vccd1 vccd1 _6343_/A sky130_fd_sc_hd__nor2_4
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6390_ _6451_/A _6390_/B vssd1 vssd1 vccd1 vccd1 _6390_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5410_ _5410_/A _5410_/B vssd1 vssd1 vccd1 vccd1 _5411_/B sky130_fd_sc_hd__xnor2_4
X_5341_ _5294_/B _5399_/B _5339_/Y vssd1 vssd1 vccd1 vccd1 _5343_/A sky130_fd_sc_hd__o21a_4
XFILLER_99_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8060_ _8077_/CLK _8060_/D vssd1 vssd1 vccd1 vccd1 _8060_/Q sky130_fd_sc_hd__dfxtp_4
X_5272_ _7213_/A _7213_/C vssd1 vssd1 vccd1 vccd1 _6871_/C sky130_fd_sc_hd__nand2_8
X_7011_ _7101_/A _7284_/A _7122_/A vssd1 vssd1 vccd1 vccd1 _7013_/B sky130_fd_sc_hd__o21ai_2
X_4223_ _4205_/Y _4221_/B _4215_/B _4221_/Y vssd1 vssd1 vccd1 vccd1 _4223_/Y sky130_fd_sc_hd__o22ai_1
X_4154_ _4175_/B _4147_/B _4211_/B vssd1 vssd1 vccd1 vccd1 _4179_/B sky130_fd_sc_hd__o21a_2
X_4085_ _8051_/Q _4096_/A vssd1 vssd1 vccd1 vccd1 _4086_/B sky130_fd_sc_hd__nand2_2
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7913_ _7913_/A _7913_/B _7914_/B vssd1 vssd1 vccd1 vccd1 _7913_/X sky130_fd_sc_hd__or3_1
XFILLER_83_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7844_ _7844_/A _7844_/B vssd1 vssd1 vccd1 vccd1 _7844_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7775_ _7789_/A _7789_/B vssd1 vssd1 vccd1 vccd1 _7777_/A sky130_fd_sc_hd__and2_1
XFILLER_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6726_ _6716_/B _6725_/A _6749_/S vssd1 vssd1 vccd1 vccd1 _6732_/C sky130_fd_sc_hd__mux2_1
XFILLER_11_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4987_ _4993_/B _4993_/A vssd1 vssd1 vccd1 vccd1 _4987_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6657_ _6656_/X _6653_/X _6733_/S vssd1 vssd1 vccd1 vccd1 _6657_/X sky130_fd_sc_hd__mux2_1
X_6588_ _6582_/X _6587_/Y _6588_/S vssd1 vssd1 vccd1 vccd1 _6590_/B sky130_fd_sc_hd__mux2_8
X_5608_ _5608_/A _5608_/B vssd1 vssd1 vccd1 vccd1 _5616_/C sky130_fd_sc_hd__nand2_2
XFILLER_117_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5539_ _5561_/A _5561_/B _5525_/Y vssd1 vssd1 vccd1 vccd1 _5549_/B sky130_fd_sc_hd__a21oi_4
XFILLER_3_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7209_ _7245_/A _7210_/B vssd1 vssd1 vccd1 vccd1 _7244_/B sky130_fd_sc_hd__nor2_2
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4910_ _4916_/B _4916_/A vssd1 vssd1 vccd1 vccd1 _4914_/B sky130_fd_sc_hd__nand2b_1
X_5890_ _5902_/A _5902_/B _5887_/Y vssd1 vssd1 vccd1 vccd1 _5900_/B sky130_fd_sc_hd__a21oi_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4841_ _4691_/A _4690_/Y _4730_/A _4730_/B vssd1 vssd1 vccd1 vccd1 _4841_/X sky130_fd_sc_hd__a211o_1
XFILLER_33_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7560_ _6267_/X _6269_/X _6270_/Y _6776_/Y vssd1 vssd1 vccd1 vccd1 _7560_/X sky130_fd_sc_hd__o31a_1
X_4772_ _5034_/A _4795_/C vssd1 vssd1 vccd1 vccd1 _4772_/Y sky130_fd_sc_hd__nand2_1
X_6511_ _6364_/A _6443_/B _6468_/B vssd1 vssd1 vccd1 vccd1 _6511_/X sky130_fd_sc_hd__a21o_1
X_7491_ _7489_/X _7490_/X _7527_/S vssd1 vssd1 vccd1 vccd1 _7491_/X sky130_fd_sc_hd__mux2_1
X_6442_ _6488_/B _6442_/B vssd1 vssd1 vccd1 vccd1 _6444_/A sky130_fd_sc_hd__or2_1
XFILLER_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6373_ _6374_/A _6374_/B _6374_/C vssd1 vssd1 vccd1 vccd1 _6373_/X sky130_fd_sc_hd__or3b_2
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5324_ _5530_/A _7358_/B vssd1 vssd1 vccd1 vccd1 _5534_/A sky130_fd_sc_hd__nor2_2
X_8043_ _8082_/CLK _8043_/D vssd1 vssd1 vccd1 vccd1 _8043_/Q sky130_fd_sc_hd__dfxtp_1
X_5255_ _5255_/A _5255_/B vssd1 vssd1 vccd1 vccd1 _5257_/B sky130_fd_sc_hd__xor2_4
X_4206_ _4196_/B _4205_/Y _4227_/S vssd1 vssd1 vccd1 vccd1 _4206_/X sky130_fd_sc_hd__o21ba_2
X_5186_ _7046_/B _5342_/B vssd1 vssd1 vccd1 vccd1 _5241_/A sky130_fd_sc_hd__nor2_4
X_4137_ _6289_/A _4136_/X _4303_/B vssd1 vssd1 vccd1 vccd1 _4137_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4068_ _8064_/Q _4068_/B vssd1 vssd1 vccd1 vccd1 _4071_/B sky130_fd_sc_hd__xnor2_4
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7827_ _7824_/Y _7825_/X _7826_/X vssd1 vssd1 vccd1 vccd1 _7827_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_24_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7758_ _7758_/A _7758_/B vssd1 vssd1 vccd1 vccd1 _7759_/B sky130_fd_sc_hd__nor2_1
X_6709_ _6709_/A _6737_/B vssd1 vssd1 vccd1 vccd1 _6709_/Y sky130_fd_sc_hd__nor2_1
X_7689_ _7748_/A _7689_/B vssd1 vssd1 vccd1 vccd1 _7707_/B sky130_fd_sc_hd__nand2_1
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout183 _4241_/X vssd1 vssd1 vccd1 vccd1 _4547_/C sky130_fd_sc_hd__buf_4
XFILLER_59_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout161 _4326_/X vssd1 vssd1 vccd1 vccd1 _7085_/A sky130_fd_sc_hd__clkbuf_16
Xfanout150 _4472_/A vssd1 vssd1 vccd1 vccd1 _4455_/A sky130_fd_sc_hd__buf_6
Xfanout172 _7366_/A vssd1 vssd1 vccd1 vccd1 _7001_/A sky130_fd_sc_hd__buf_12
XFILLER_47_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout194 _6035_/A0 vssd1 vssd1 vccd1 vccd1 _4548_/A sky130_fd_sc_hd__buf_4
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5040_/A _5040_/B vssd1 vssd1 vccd1 vccd1 _5040_/Y sky130_fd_sc_hd__nor2_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6991_ _6991_/A _6991_/B _6991_/C vssd1 vssd1 vccd1 vccd1 _6992_/B sky130_fd_sc_hd__or3_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5942_ _5942_/A _5942_/B vssd1 vssd1 vccd1 vccd1 _6135_/B sky130_fd_sc_hd__or2_4
XFILLER_21_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5873_ _5871_/A _5871_/B _5872_/Y vssd1 vssd1 vccd1 vccd1 _5875_/B sky130_fd_sc_hd__o21a_1
X_7612_ _7643_/A _7643_/B vssd1 vssd1 vccd1 vccd1 _7612_/X sky130_fd_sc_hd__xor2_4
XFILLER_61_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4824_ _4854_/A _4818_/Y _4822_/X _4805_/C vssd1 vssd1 vccd1 vccd1 _4826_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7543_ _7766_/B _7543_/B _7543_/C _7543_/D vssd1 vssd1 vccd1 vccd1 _7544_/D sky130_fd_sc_hd__or4_1
X_4755_ _4854_/A _4768_/B vssd1 vssd1 vccd1 vccd1 _4763_/A sky130_fd_sc_hd__or2_1
XFILLER_119_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4686_ _4685_/A _4685_/C _4727_/A vssd1 vssd1 vccd1 vccd1 _4686_/Y sky130_fd_sc_hd__a21oi_1
X_7474_ _7474_/A _7474_/B vssd1 vssd1 vccd1 vccd1 _7474_/X sky130_fd_sc_hd__xor2_2
X_6425_ _6488_/B _6425_/B vssd1 vssd1 vccd1 vccd1 _6475_/A sky130_fd_sc_hd__nor2_2
XFILLER_103_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6356_ _6386_/A _6359_/A vssd1 vssd1 vccd1 vccd1 _6364_/A sky130_fd_sc_hd__and2_2
XFILLER_115_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5307_ _5842_/B _5723_/A _5516_/A _5715_/A vssd1 vssd1 vccd1 vccd1 _5307_/X sky130_fd_sc_hd__o2bb2a_2
X_8026_ _8082_/CLK _8026_/D vssd1 vssd1 vccd1 vccd1 _8026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6287_ _6284_/X _6285_/X _6286_/Y vssd1 vssd1 vccd1 vccd1 _6287_/Y sky130_fd_sc_hd__a21oi_1
X_5238_ _5285_/A _5238_/B vssd1 vssd1 vccd1 vccd1 _6172_/A sky130_fd_sc_hd__xor2_4
XFILLER_96_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5169_ _5169_/A _5169_/B vssd1 vssd1 vccd1 vccd1 _5170_/B sky130_fd_sc_hd__and2_1
XFILLER_29_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4540_ _4540_/A _4540_/B vssd1 vssd1 vccd1 vccd1 _4544_/A sky130_fd_sc_hd__xnor2_4
X_4471_ _4451_/A _4451_/C _4451_/B vssd1 vssd1 vccd1 vccd1 _4495_/A sky130_fd_sc_hd__a21boi_4
X_6210_ _6254_/S _6199_/X _6209_/X vssd1 vssd1 vccd1 vccd1 _6210_/X sky130_fd_sc_hd__a21o_1
X_7190_ _7190_/A _7190_/B vssd1 vssd1 vccd1 vccd1 _7202_/A sky130_fd_sc_hd__xnor2_4
X_6141_ _6138_/Y _6140_/Y _6262_/S vssd1 vssd1 vccd1 vccd1 _6245_/B sky130_fd_sc_hd__mux2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6072_ _6059_/B _6071_/Y _6068_/A vssd1 vssd1 vccd1 vccd1 _6072_/Y sky130_fd_sc_hd__o21ai_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5023_ _5018_/A _5018_/B _5018_/C vssd1 vssd1 vccd1 vccd1 _5024_/B sky130_fd_sc_hd__a21o_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6974_ _7030_/A _7247_/C vssd1 vssd1 vccd1 vccd1 _7021_/A sky130_fd_sc_hd__nor2_1
X_5925_ _5925_/A _5925_/B vssd1 vssd1 vccd1 vccd1 _5925_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5856_ _5855_/A _5855_/B _5921_/A _5855_/C vssd1 vssd1 vccd1 vccd1 _5857_/B sky130_fd_sc_hd__o31ai_1
X_4807_ _4854_/A _4805_/X _4804_/Y vssd1 vssd1 vccd1 vccd1 _4809_/B sky130_fd_sc_hd__o21a_1
XFILLER_21_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5787_ _5787_/A _5787_/B vssd1 vssd1 vccd1 vccd1 _6205_/A sky130_fd_sc_hd__nor2_8
XFILLER_119_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7526_ _7510_/X _7514_/X _7515_/S vssd1 vssd1 vccd1 vccd1 _7526_/X sky130_fd_sc_hd__o21ba_1
X_4738_ _4738_/A _4738_/B vssd1 vssd1 vccd1 vccd1 _4738_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_119_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7457_ _7403_/C _7502_/B vssd1 vssd1 vccd1 vccd1 _7457_/Y sky130_fd_sc_hd__nand2b_1
X_4669_ _4668_/A _4668_/C _4668_/B vssd1 vssd1 vccd1 vccd1 _4670_/C sky130_fd_sc_hd__a21o_1
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6408_ _5204_/X _4343_/Y _6456_/S vssd1 vssd1 vccd1 vccd1 _6408_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7388_ _6892_/A _6892_/B _7448_/A vssd1 vssd1 vccd1 vccd1 _7452_/A sky130_fd_sc_hd__o21bai_2
XFILLER_1_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6339_ _6338_/A _6338_/B _6338_/C vssd1 vssd1 vccd1 vccd1 _6339_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_88_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8009_ _8057_/CLK _8009_/D vssd1 vssd1 vccd1 vccd1 _8009_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_95_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5710_ _5943_/B _5942_/A _5943_/A vssd1 vssd1 vccd1 vccd1 _5710_/X sky130_fd_sc_hd__o21a_1
X_6690_ _6689_/X _6667_/X _6691_/A vssd1 vssd1 vccd1 vccd1 _6690_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5641_ _5641_/A _5641_/B vssd1 vssd1 vccd1 vccd1 _5686_/B sky130_fd_sc_hd__xor2_4
X_5572_ _5722_/A _5722_/B _7306_/B vssd1 vssd1 vccd1 vccd1 _5631_/C sky130_fd_sc_hd__and3_2
XFILLER_116_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7311_ _7311_/A _7371_/B _7311_/C vssd1 vssd1 vccd1 vccd1 _7336_/A sky130_fd_sc_hd__or3_4
X_4523_ _4521_/A _4521_/B _4522_/Y vssd1 vssd1 vccd1 vccd1 _4545_/A sky130_fd_sc_hd__o21a_2
X_7242_ _7242_/A _7242_/B vssd1 vssd1 vccd1 vccd1 _7243_/B sky130_fd_sc_hd__and2_1
X_4454_ _4393_/A _4393_/B _4392_/A vssd1 vssd1 vccd1 vccd1 _4461_/A sky130_fd_sc_hd__o21ai_4
X_7173_ _7173_/A _7173_/B vssd1 vssd1 vccd1 vccd1 _7211_/B sky130_fd_sc_hd__xor2_4
X_4385_ _4998_/A _7285_/A _4585_/B _7281_/A vssd1 vssd1 vccd1 vccd1 _4386_/D sky130_fd_sc_hd__a22o_2
XFILLER_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6124_ _6123_/A _6123_/B _6123_/Y _6139_/B vssd1 vssd1 vccd1 vccd1 _6150_/B sky130_fd_sc_hd__o211a_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6055_ _6055_/A _6055_/B vssd1 vssd1 vccd1 vccd1 _6058_/B sky130_fd_sc_hd__or2_4
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _5009_/A _5009_/B _5004_/Y vssd1 vssd1 vccd1 vccd1 _5008_/B sky130_fd_sc_hd__a21oi_4
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ _6957_/A _6957_/B _6957_/C vssd1 vssd1 vccd1 vccd1 _6958_/B sky130_fd_sc_hd__or3_1
XFILLER_53_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6888_ _6888_/A _6888_/B vssd1 vssd1 vccd1 vccd1 _6894_/B sky130_fd_sc_hd__xnor2_1
XFILLER_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5908_ _5908_/A _7319_/B _5908_/C vssd1 vssd1 vccd1 vccd1 _5915_/A sky130_fd_sc_hd__and3_1
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5839_ _5837_/A _5838_/A _5837_/B _5851_/B _5829_/Y vssd1 vssd1 vccd1 vccd1 _5843_/A
+ sky130_fd_sc_hd__a32o_2
X_7509_ _7508_/X _7487_/Y _7513_/S vssd1 vssd1 vccd1 vccd1 _7509_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4170_ _8076_/Q _4170_/B vssd1 vssd1 vccd1 vccd1 _4170_/X sky130_fd_sc_hd__xor2_4
XFILLER_95_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7860_ _7908_/A _7886_/C vssd1 vssd1 vccd1 vccd1 _7860_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6811_ _6812_/A _6812_/B _6812_/C vssd1 vssd1 vccd1 vccd1 _6827_/B sky130_fd_sc_hd__o21ai_4
XFILLER_63_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7791_ _7822_/A _7791_/B vssd1 vssd1 vccd1 vccd1 _7793_/A sky130_fd_sc_hd__nor2_2
XFILLER_90_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6742_ _6741_/X _6657_/X _6753_/S vssd1 vssd1 vccd1 vccd1 _6742_/X sky130_fd_sc_hd__mux2_1
X_6673_ _6672_/Y _6670_/X _6751_/S vssd1 vssd1 vccd1 vccd1 _6674_/A sky130_fd_sc_hd__mux2_1
X_5624_ _5566_/B _5666_/B _5623_/Y vssd1 vssd1 vccd1 vccd1 _5663_/B sky130_fd_sc_hd__a21oi_2
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5555_ _5607_/A _5607_/B vssd1 vssd1 vccd1 vccd1 _5608_/A sky130_fd_sc_hd__nand2_2
XFILLER_117_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5486_ _5484_/Y _5486_/B vssd1 vssd1 vccd1 vccd1 _5487_/B sky130_fd_sc_hd__and2b_2
X_4506_ _4506_/A _4506_/B vssd1 vssd1 vccd1 vccd1 _4511_/A sky130_fd_sc_hd__xnor2_4
X_7225_ _7030_/A _7210_/B _7086_/B vssd1 vssd1 vccd1 vccd1 _7227_/C sky130_fd_sc_hd__o21ai_2
X_4437_ _4455_/A _4430_/C _4407_/B _4430_/A vssd1 vssd1 vccd1 vccd1 _4437_/X sky130_fd_sc_hd__a211o_1
XFILLER_104_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7156_ _7156_/A _7156_/B vssd1 vssd1 vccd1 vccd1 _7197_/B sky130_fd_sc_hd__xnor2_2
XFILLER_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6107_ _6259_/C _6192_/B _6093_/X vssd1 vssd1 vccd1 vccd1 _6107_/X sky130_fd_sc_hd__or3b_1
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ _5090_/A _7247_/A _4654_/A _4585_/B vssd1 vssd1 vccd1 vccd1 _4387_/A sky130_fd_sc_hd__or4b_4
XFILLER_86_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4299_ _4056_/S _5993_/B _4298_/X _5135_/C1 vssd1 vssd1 vccd1 vccd1 _4301_/A sky130_fd_sc_hd__a211o_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7087_ _7087_/A _7087_/B vssd1 vssd1 vccd1 vccd1 _7141_/A sky130_fd_sc_hd__xnor2_4
XFILLER_100_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6038_ _6037_/B _6038_/B vssd1 vssd1 vccd1 vccd1 _6058_/A sky130_fd_sc_hd__and2b_1
XFILLER_58_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7989_ _8025_/Q _8065_/Q _7990_/S vssd1 vssd1 vccd1 vccd1 _8065_/D sky130_fd_sc_hd__mux2_1
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5340_ _5367_/A _5516_/A vssd1 vssd1 vccd1 vccd1 _5399_/B sky130_fd_sc_hd__or2_4
XFILLER_114_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5271_ _5977_/A _5271_/B vssd1 vssd1 vccd1 vccd1 _5271_/Y sky130_fd_sc_hd__nor2_1
X_4222_ _4205_/Y _4221_/B _4215_/B _4221_/Y vssd1 vssd1 vccd1 vccd1 _4222_/X sky130_fd_sc_hd__o22a_1
X_7010_ _7101_/A _7284_/A _7122_/A vssd1 vssd1 vccd1 vccd1 _7013_/A sky130_fd_sc_hd__or3_1
X_4153_ _4216_/B _6289_/B vssd1 vssd1 vccd1 vccd1 _4230_/A sky130_fd_sc_hd__nor2_1
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4084_ _6326_/A _4084_/B vssd1 vssd1 vccd1 vccd1 _4084_/X sky130_fd_sc_hd__xor2_2
XFILLER_68_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7912_ _7766_/B _7709_/Y _7766_/Y vssd1 vssd1 vccd1 vccd1 _7914_/B sky130_fd_sc_hd__a21o_1
XFILLER_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7843_ _7793_/Y _7823_/Y _7649_/A vssd1 vssd1 vccd1 vccd1 _7844_/B sky130_fd_sc_hd__a21o_1
XFILLER_23_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7774_ _6636_/Y _6763_/X _7773_/X vssd1 vssd1 vccd1 vccd1 _7789_/B sky130_fd_sc_hd__a21oi_1
X_4986_ _4986_/A _4986_/B vssd1 vssd1 vccd1 vccd1 _4993_/B sky130_fd_sc_hd__xnor2_4
XFILLER_23_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6725_ _6725_/A vssd1 vssd1 vccd1 vccd1 _6725_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6656_ _6713_/S _6651_/Y _6652_/Y _6655_/Y vssd1 vssd1 vccd1 vccd1 _6656_/X sky130_fd_sc_hd__a22o_1
X_6587_ _6562_/A _6539_/A _6586_/Y _6585_/X _6515_/Y vssd1 vssd1 vccd1 vccd1 _6587_/Y
+ sky130_fd_sc_hd__o32ai_4
X_5607_ _5607_/A _5607_/B vssd1 vssd1 vccd1 vccd1 _5608_/B sky130_fd_sc_hd__or2_1
X_5538_ _5538_/A _5538_/B vssd1 vssd1 vccd1 vccd1 _5561_/B sky130_fd_sc_hd__xnor2_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5469_ _5470_/A _5470_/B vssd1 vssd1 vccd1 vccd1 _5469_/X sky130_fd_sc_hd__and2b_1
X_7208_ _7113_/X _7206_/Y _7212_/A vssd1 vssd1 vccd1 vccd1 _7244_/A sky130_fd_sc_hd__a21o_4
XFILLER_99_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7139_ _7182_/A _7182_/B vssd1 vssd1 vccd1 vccd1 _7143_/A sky130_fd_sc_hd__and2_2
XFILLER_86_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4840_ _5013_/A _7001_/A _4728_/X _4838_/X _4839_/X vssd1 vssd1 vccd1 vccd1 _4840_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6510_ _6377_/A _6509_/X _6376_/A vssd1 vssd1 vccd1 vccd1 _6510_/Y sky130_fd_sc_hd__a21oi_1
X_4771_ _4773_/A _5014_/A _4795_/C vssd1 vssd1 vccd1 vccd1 _4820_/S sky130_fd_sc_hd__or3_4
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7490_ _7488_/X _7471_/X _7513_/S vssd1 vssd1 vccd1 vccd1 _7490_/X sky130_fd_sc_hd__mux2_1
X_6441_ _6402_/X _6440_/X _6441_/S vssd1 vssd1 vccd1 vccd1 _6442_/B sky130_fd_sc_hd__mux2_1
X_6372_ _7085_/A _7114_/B _6456_/S vssd1 vssd1 vccd1 vccd1 _6374_/C sky130_fd_sc_hd__mux2_1
X_5323_ _5145_/B _5145_/C _5322_/A _5268_/A vssd1 vssd1 vccd1 vccd1 _5323_/X sky130_fd_sc_hd__a211o_2
XFILLER_114_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8042_ _8082_/CLK _8042_/D vssd1 vssd1 vccd1 vccd1 _8042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5254_ _5782_/A _5185_/Y _5431_/B _5250_/Y vssd1 vssd1 vccd1 vccd1 _5257_/A sky130_fd_sc_hd__a31o_4
XFILLER_87_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4205_ _4228_/A _4216_/C vssd1 vssd1 vccd1 vccd1 _4205_/Y sky130_fd_sc_hd__nand2_1
X_5185_ _5672_/A vssd1 vssd1 vccd1 vccd1 _5185_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4136_ _4059_/B _4303_/C _4135_/X vssd1 vssd1 vccd1 vccd1 _4136_/X sky130_fd_sc_hd__o21a_1
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4067_ _8063_/Q _5107_/B _4066_/A vssd1 vssd1 vccd1 vccd1 _4068_/B sky130_fd_sc_hd__o21a_2
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7826_ _6268_/X _7812_/Y _7813_/X _7819_/Y vssd1 vssd1 vccd1 vccd1 _7826_/X sky130_fd_sc_hd__a31o_2
XFILLER_24_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7757_ _7702_/A _7757_/B _7758_/B _7757_/D vssd1 vssd1 vccd1 vccd1 _7833_/A sky130_fd_sc_hd__and4b_4
XFILLER_11_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4969_ _5020_/B _4969_/B vssd1 vssd1 vccd1 vccd1 _5003_/B sky130_fd_sc_hd__xor2_4
X_6708_ _6686_/X _6693_/X _6751_/S vssd1 vssd1 vccd1 vccd1 _6708_/X sky130_fd_sc_hd__mux2_1
X_7688_ _7687_/A _7687_/B _7687_/C vssd1 vssd1 vccd1 vccd1 _7689_/B sky130_fd_sc_hd__a21o_1
X_6639_ _6751_/S _6749_/S _7718_/S _6638_/A vssd1 vssd1 vccd1 vccd1 _6640_/A sky130_fd_sc_hd__o211a_1
XFILLER_118_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout140 _7116_/A vssd1 vssd1 vccd1 vccd1 _4441_/A sky130_fd_sc_hd__buf_4
XFILLER_59_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout162 _4326_/X vssd1 vssd1 vccd1 vccd1 _6873_/A sky130_fd_sc_hd__buf_4
Xfanout173 _7366_/A vssd1 vssd1 vccd1 vccd1 _7334_/B sky130_fd_sc_hd__buf_4
Xfanout151 _4472_/A vssd1 vssd1 vccd1 vccd1 _4430_/B sky130_fd_sc_hd__buf_4
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout195 _4322_/A vssd1 vssd1 vccd1 vccd1 _6035_/A0 sky130_fd_sc_hd__buf_4
Xfanout184 _4548_/C vssd1 vssd1 vccd1 vccd1 _4354_/A sky130_fd_sc_hd__buf_12
XFILLER_74_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6990_ _6992_/A _6990_/B vssd1 vssd1 vccd1 vccd1 _7442_/A sky130_fd_sc_hd__xor2_2
XFILLER_93_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5941_ _5709_/B _5941_/B vssd1 vssd1 vccd1 vccd1 _5942_/B sky130_fd_sc_hd__and2b_1
XFILLER_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5872_ _5877_/A _5877_/B vssd1 vssd1 vccd1 vccd1 _5872_/Y sky130_fd_sc_hd__nand2b_1
X_7611_ _7643_/B _7611_/B _7611_/C _7611_/D vssd1 vssd1 vccd1 vccd1 _7757_/D sky130_fd_sc_hd__and4b_4
X_4823_ _4805_/C _4822_/X _4818_/Y vssd1 vssd1 vccd1 vccd1 _4854_/B sky130_fd_sc_hd__a21o_1
X_7542_ _7542_/A _7542_/B _7542_/C _7542_/D vssd1 vssd1 vccd1 vccd1 _7543_/D sky130_fd_sc_hd__or4_1
X_4754_ _4757_/B _4754_/B vssd1 vssd1 vccd1 vccd1 _4768_/B sky130_fd_sc_hd__nand2_2
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7473_ _7471_/X _7472_/X _7513_/S vssd1 vssd1 vccd1 vccd1 _7473_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4685_ _4685_/A _4727_/A _4685_/C vssd1 vssd1 vccd1 vccd1 _4685_/X sky130_fd_sc_hd__and3_1
X_6424_ _6383_/B _6423_/Y _6441_/S vssd1 vssd1 vccd1 vccd1 _6425_/B sky130_fd_sc_hd__mux2_1
XFILLER_108_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6355_ _6374_/A _6492_/A _6354_/X vssd1 vssd1 vccd1 vccd1 _6355_/X sky130_fd_sc_hd__or3b_4
XFILLER_115_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6286_ _4059_/B _4172_/B _4169_/Y _4062_/B vssd1 vssd1 vccd1 vccd1 _6286_/Y sky130_fd_sc_hd__o22ai_1
X_5306_ _5621_/A _5305_/Y _5306_/S vssd1 vssd1 vccd1 vccd1 _5504_/A sky130_fd_sc_hd__mux2_4
X_8025_ _8080_/CLK _8025_/D vssd1 vssd1 vccd1 vccd1 _8025_/Q sky130_fd_sc_hd__dfxtp_1
X_5237_ _5961_/A _5237_/B vssd1 vssd1 vccd1 vccd1 _5238_/B sky130_fd_sc_hd__and2_2
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5168_ _5169_/A _5169_/B vssd1 vssd1 vccd1 vccd1 _5232_/A sky130_fd_sc_hd__nor2_2
XFILLER_56_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4119_ _4063_/A _4116_/Y _4117_/Y _4078_/B vssd1 vssd1 vccd1 vccd1 _4119_/Y sky130_fd_sc_hd__o31ai_4
XFILLER_84_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5099_ _5063_/A _5063_/B _4786_/A vssd1 vssd1 vccd1 vccd1 _5100_/B sky130_fd_sc_hd__a21bo_2
XFILLER_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7809_ _7908_/A _7833_/C vssd1 vssd1 vccd1 vccd1 _7809_/X sky130_fd_sc_hd__and2b_1
XFILLER_24_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4470_ _4467_/X _4468_/Y _4394_/Y _4566_/A vssd1 vssd1 vccd1 vccd1 _4497_/B sky130_fd_sc_hd__o211a_2
XFILLER_109_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6140_ _6115_/X _6156_/A _6135_/Y _6177_/A _6139_/Y vssd1 vssd1 vccd1 vccd1 _6140_/Y
+ sky130_fd_sc_hd__a221oi_4
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6071_/A vssd1 vssd1 vccd1 vccd1 _6071_/Y sky130_fd_sc_hd__inv_2
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5022_/A _5022_/B vssd1 vssd1 vccd1 vccd1 _5043_/A sky130_fd_sc_hd__xor2_4
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6973_ _6975_/A _6975_/B vssd1 vssd1 vccd1 vccd1 _6973_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5924_ _5924_/A _5924_/B vssd1 vssd1 vccd1 vccd1 _5928_/A sky130_fd_sc_hd__xor2_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5855_ _5855_/A _5855_/B _5855_/C _5921_/A vssd1 vssd1 vccd1 vccd1 _5857_/A sky130_fd_sc_hd__or4_1
X_4806_ _4806_/A _4806_/B vssd1 vssd1 vccd1 vccd1 _4817_/B sky130_fd_sc_hd__xnor2_1
X_5786_ _5786_/A _5786_/B vssd1 vssd1 vccd1 vccd1 _5787_/B sky130_fd_sc_hd__and2_2
X_7525_ _7525_/A vssd1 vssd1 vccd1 vccd1 _7525_/Y sky130_fd_sc_hd__inv_2
X_4737_ _4846_/A _4846_/B _4848_/B _4736_/X vssd1 vssd1 vccd1 vccd1 _4738_/B sky130_fd_sc_hd__a31o_2
XFILLER_119_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7456_ _7453_/X _7455_/X _7502_/B vssd1 vssd1 vccd1 vccd1 _7456_/X sky130_fd_sc_hd__mux2_1
X_4668_ _4668_/A _4668_/B _4668_/C vssd1 vssd1 vccd1 vccd1 _4670_/B sky130_fd_sc_hd__nand3_2
X_6407_ _6407_/A _6407_/B vssd1 vssd1 vccd1 vccd1 _6474_/B sky130_fd_sc_hd__or2_2
XFILLER_115_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7387_ _7447_/B _7387_/B vssd1 vssd1 vccd1 vccd1 _7448_/A sky130_fd_sc_hd__and2b_1
X_4599_ _4599_/A _4599_/B _4599_/C vssd1 vssd1 vccd1 vccd1 _4606_/A sky130_fd_sc_hd__and3_4
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6338_ _6338_/A _6338_/B _6338_/C vssd1 vssd1 vccd1 vccd1 _6338_/X sky130_fd_sc_hd__or3_1
XFILLER_88_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6269_ _8009_/Q _7558_/A _8010_/Q vssd1 vssd1 vccd1 vccd1 _6269_/X sky130_fd_sc_hd__or3b_4
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8008_ _8057_/CLK _8008_/D vssd1 vssd1 vccd1 vccd1 _8008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5640_ _5641_/A _5641_/B vssd1 vssd1 vccd1 vccd1 _5652_/A sky130_fd_sc_hd__or2_4
XFILLER_31_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5571_ _5672_/A _5797_/A vssd1 vssd1 vccd1 vccd1 _5576_/A sky130_fd_sc_hd__or2_4
X_7310_ _7332_/A _7310_/B vssd1 vssd1 vccd1 vccd1 _7312_/A sky130_fd_sc_hd__xnor2_4
X_4522_ _4546_/B _4546_/A vssd1 vssd1 vccd1 vccd1 _4522_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4453_ _4453_/A _4453_/B _4453_/C vssd1 vssd1 vccd1 vccd1 _4566_/A sky130_fd_sc_hd__nand3_4
X_7241_ _7241_/A _7241_/B vssd1 vssd1 vccd1 vccd1 _7266_/A sky130_fd_sc_hd__xnor2_4
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7172_ _7215_/A _7210_/B vssd1 vssd1 vccd1 vccd1 _7211_/A sky130_fd_sc_hd__or2_4
X_4384_ _5019_/A vssd1 vssd1 vccd1 vccd1 _4989_/A sky130_fd_sc_hd__clkinv_4
XFILLER_112_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6123_ _6123_/A _6123_/B vssd1 vssd1 vccd1 vccd1 _6123_/Y sky130_fd_sc_hd__nand2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6054_ _6054_/A _6054_/B vssd1 vssd1 vccd1 vccd1 _6055_/B sky130_fd_sc_hd__and2_1
XFILLER_98_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5005_ _5005_/A _5005_/B vssd1 vssd1 vccd1 vccd1 _5009_/B sky130_fd_sc_hd__xor2_4
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6956_ _6957_/B _6957_/C _6957_/A vssd1 vssd1 vccd1 vccd1 _6966_/A sky130_fd_sc_hd__o21ai_2
X_5907_ _5917_/A _5922_/A vssd1 vssd1 vccd1 vccd1 _5907_/Y sky130_fd_sc_hd__nand2_1
X_6887_ _6887_/A _6887_/B vssd1 vssd1 vccd1 vccd1 _6894_/A sky130_fd_sc_hd__and2_1
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5838_ _5838_/A _5838_/B vssd1 vssd1 vccd1 vccd1 _5851_/B sky130_fd_sc_hd__xnor2_4
XFILLER_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5769_ _6971_/B _5853_/B vssd1 vssd1 vccd1 vccd1 _5800_/D sky130_fd_sc_hd__or2_1
XFILLER_108_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7508_ _7508_/A _7508_/B vssd1 vssd1 vccd1 vccd1 _7508_/X sky130_fd_sc_hd__xor2_1
XFILLER_108_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7439_ _7439_/A _7439_/B vssd1 vssd1 vccd1 vccd1 _7439_/X sky130_fd_sc_hd__xor2_1
XFILLER_103_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6810_ _6810_/A _6810_/B vssd1 vssd1 vccd1 vccd1 _6812_/C sky130_fd_sc_hd__and2_1
XFILLER_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7790_ _7777_/A _7789_/C _7773_/X vssd1 vssd1 vccd1 vccd1 _7791_/B sky130_fd_sc_hd__o21bai_1
XFILLER_90_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6741_ _6739_/X _6740_/X _6751_/S vssd1 vssd1 vccd1 vccd1 _6741_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6672_ _6672_/A vssd1 vssd1 vccd1 vccd1 _6672_/Y sky130_fd_sc_hd__inv_2
X_5623_ _7114_/B _5858_/B _5621_/Y vssd1 vssd1 vccd1 vccd1 _5623_/Y sky130_fd_sc_hd__a21oi_1
X_5554_ _5554_/A _5554_/B vssd1 vssd1 vccd1 vccd1 _5607_/B sky130_fd_sc_hd__xnor2_1
XFILLER_117_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5485_ _5485_/A _5485_/B vssd1 vssd1 vccd1 vccd1 _5486_/B sky130_fd_sc_hd__nand2_2
X_4505_ _4505_/A _4505_/B vssd1 vssd1 vccd1 vccd1 _4506_/B sky130_fd_sc_hd__xnor2_4
X_4436_ _4436_/A _4558_/B vssd1 vssd1 vccd1 vccd1 _4508_/A sky130_fd_sc_hd__nor2_8
X_7224_ _7212_/A _7212_/B _7218_/X vssd1 vssd1 vccd1 vccd1 _7228_/A sky130_fd_sc_hd__a21o_2
X_7155_ _7155_/A _7155_/B vssd1 vssd1 vccd1 vccd1 _7477_/A sky130_fd_sc_hd__nor2_2
X_4367_ _4494_/A _4363_/X _4366_/X _4362_/X vssd1 vssd1 vccd1 vccd1 _4367_/X sky130_fd_sc_hd__a31o_1
XFILLER_113_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6106_ _6099_/A _6099_/B _6110_/A _6093_/B _6132_/B vssd1 vssd1 vccd1 vccd1 _6111_/C
+ sky130_fd_sc_hd__a2111o_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4298_ _4074_/Y _4118_/X _4050_/Y _4071_/Y vssd1 vssd1 vccd1 vccd1 _4298_/X sky130_fd_sc_hd__o211a_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7086_ _7086_/A _7086_/B vssd1 vssd1 vccd1 vccd1 _7087_/B sky130_fd_sc_hd__or2_4
X_6037_ _6038_/B _6037_/B vssd1 vssd1 vccd1 vccd1 _6039_/B sky130_fd_sc_hd__and2_1
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7988_ _8024_/Q _8064_/Q _7990_/S vssd1 vssd1 vccd1 vccd1 _8064_/D sky130_fd_sc_hd__mux2_1
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6939_ _6939_/A _6939_/B vssd1 vssd1 vccd1 vccd1 _6991_/A sky130_fd_sc_hd__xnor2_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5270_ _5977_/B _5083_/X _5084_/X _5268_/X vssd1 vssd1 vccd1 vccd1 _7213_/C sky130_fd_sc_hd__a31o_4
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4221_ _8067_/Q _4221_/B vssd1 vssd1 vccd1 vccd1 _4221_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4152_ _8079_/Q _4152_/B vssd1 vssd1 vccd1 vccd1 _6289_/B sky130_fd_sc_hd__xnor2_4
X_4083_ _8053_/Q _4083_/B vssd1 vssd1 vccd1 vccd1 _4084_/B sky130_fd_sc_hd__xnor2_4
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7911_ _7929_/B _7911_/B vssd1 vssd1 vccd1 vccd1 _7911_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_48_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7842_ _7895_/A _7842_/B vssd1 vssd1 vccd1 vccd1 _7844_/A sky130_fd_sc_hd__or2_2
XFILLER_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7773_ _7773_/A _7894_/A vssd1 vssd1 vccd1 vccd1 _7773_/X sky130_fd_sc_hd__and2_2
X_4985_ _4984_/B _4984_/C _4984_/A vssd1 vssd1 vccd1 vccd1 _4993_/A sky130_fd_sc_hd__a21bo_4
X_6724_ _6722_/X _6723_/X _7581_/S vssd1 vssd1 vccd1 vccd1 _6725_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6655_ _6691_/A _6655_/B vssd1 vssd1 vccd1 vccd1 _6655_/Y sky130_fd_sc_hd__nor2_2
X_6586_ _6534_/Y _6538_/B _6539_/B vssd1 vssd1 vccd1 vccd1 _6586_/Y sky130_fd_sc_hd__a21oi_2
X_5606_ _5660_/B _5660_/A vssd1 vssd1 vccd1 vccd1 _5616_/B sky130_fd_sc_hd__nand2b_2
X_5537_ _5537_/A _5537_/B vssd1 vssd1 vccd1 vccd1 _5538_/B sky130_fd_sc_hd__xor2_4
XFILLER_117_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5468_ _5468_/A _5468_/B vssd1 vssd1 vccd1 vccd1 _5470_/B sky130_fd_sc_hd__xnor2_4
X_7207_ _7334_/A _7334_/B _7235_/B _7294_/B vssd1 vssd1 vccd1 vccd1 _7212_/A sky130_fd_sc_hd__nor4_4
XFILLER_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4419_ _4441_/A _4662_/A _4483_/A vssd1 vssd1 vccd1 vccd1 _4419_/X sky130_fd_sc_hd__a21o_1
X_5399_ _5399_/A _5399_/B vssd1 vssd1 vccd1 vccd1 _5401_/A sky130_fd_sc_hd__xor2_4
X_7138_ _7261_/A _7344_/B vssd1 vssd1 vccd1 vccd1 _7182_/B sky130_fd_sc_hd__nor2_2
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7069_ _7123_/A _7306_/B _7127_/A _7066_/Y vssd1 vssd1 vccd1 vccd1 _7076_/A sky130_fd_sc_hd__a31o_4
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4770_ _4775_/A _4775_/B vssd1 vssd1 vccd1 vccd1 _4851_/A sky130_fd_sc_hd__and2_4
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6440_ _6422_/B _6439_/X _6484_/S vssd1 vssd1 vccd1 vccd1 _6440_/X sky130_fd_sc_hd__mux2_1
X_6371_ _6492_/A _6371_/B vssd1 vssd1 vccd1 vccd1 _6374_/B sky130_fd_sc_hd__or2_4
X_5322_ _5322_/A _5322_/B vssd1 vssd1 vccd1 vccd1 _5923_/A sky130_fd_sc_hd__nor2_8
XFILLER_114_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8041_ _8082_/CLK _8041_/D vssd1 vssd1 vccd1 vccd1 _8041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5253_ _5259_/A _5399_/A _5252_/X vssd1 vssd1 vccd1 vccd1 _5431_/B sky130_fd_sc_hd__o21a_2
X_4204_ _8069_/Q _4204_/B vssd1 vssd1 vccd1 vccd1 _4204_/Y sky130_fd_sc_hd__xnor2_2
X_5184_ _5184_/A _5184_/B vssd1 vssd1 vccd1 vccd1 _5342_/B sky130_fd_sc_hd__xor2_4
X_4135_ _4078_/A _4119_/Y _4077_/B _4111_/A vssd1 vssd1 vccd1 vccd1 _4135_/X sky130_fd_sc_hd__a211o_1
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4066_ _4066_/A _5107_/B vssd1 vssd1 vccd1 vccd1 _4072_/B sky130_fd_sc_hd__nand2_2
XFILLER_83_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7825_ _7649_/A _7793_/Y _7823_/Y _7923_/A vssd1 vssd1 vccd1 vccd1 _7825_/X sky130_fd_sc_hd__o31a_2
X_7756_ _7784_/A _6264_/X _7908_/A vssd1 vssd1 vccd1 vccd1 _7758_/B sky130_fd_sc_hd__o21ba_1
XFILLER_51_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4968_ _4968_/A _4968_/B vssd1 vssd1 vccd1 vccd1 _4969_/B sky130_fd_sc_hd__xor2_4
X_6707_ _6753_/S _6707_/B vssd1 vssd1 vccd1 vccd1 _6707_/X sky130_fd_sc_hd__and2_1
X_7687_ _7687_/A _7687_/B _7687_/C vssd1 vssd1 vccd1 vccd1 _7748_/A sky130_fd_sc_hd__nand3_2
X_4899_ _5090_/A _5013_/C vssd1 vssd1 vccd1 vccd1 _4900_/B sky130_fd_sc_hd__nor2_2
X_6638_ _6638_/A vssd1 vssd1 vccd1 vccd1 _6638_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6569_ _6584_/A _6583_/B _6572_/A _7886_/A vssd1 vssd1 vccd1 vccd1 _6570_/B sky130_fd_sc_hd__a31o_2
XFILLER_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout130 _6021_/A0 vssd1 vssd1 vccd1 vccd1 _5135_/C1 sky130_fd_sc_hd__buf_6
XFILLER_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout152 _7123_/A vssd1 vssd1 vccd1 vccd1 _4472_/A sky130_fd_sc_hd__buf_4
Xfanout141 _7116_/A vssd1 vssd1 vccd1 vccd1 _7245_/A sky130_fd_sc_hd__buf_4
Xfanout174 _4548_/X vssd1 vssd1 vccd1 vccd1 _7366_/A sky130_fd_sc_hd__buf_8
Xfanout163 _7027_/A vssd1 vssd1 vccd1 vccd1 _7136_/A sky130_fd_sc_hd__buf_6
Xfanout185 _4240_/Y vssd1 vssd1 vccd1 vccd1 _4548_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_59_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout196 _4207_/X vssd1 vssd1 vccd1 vccd1 _4322_/A sky130_fd_sc_hd__buf_2
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5940_ _6205_/A _6205_/B _6137_/A _5785_/X vssd1 vssd1 vccd1 vccd1 _5940_/X sky130_fd_sc_hd__a31o_2
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7610_ _6225_/X _7831_/B _7784_/A vssd1 vssd1 vccd1 vccd1 _7643_/B sky130_fd_sc_hd__mux2_4
X_5871_ _5871_/A _5871_/B vssd1 vssd1 vccd1 vccd1 _5877_/B sky130_fd_sc_hd__xor2_2
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4822_ _4851_/A _4927_/A _4926_/A vssd1 vssd1 vccd1 vccd1 _4822_/X sky130_fd_sc_hd__a21o_1
X_7541_ _7526_/X _7529_/B _7535_/A vssd1 vssd1 vccd1 vccd1 _7541_/Y sky130_fd_sc_hd__o21ai_1
X_4753_ _4991_/A _5090_/B _4750_/X vssd1 vssd1 vccd1 vccd1 _4754_/B sky130_fd_sc_hd__a21o_1
X_7472_ _7472_/A _7472_/B vssd1 vssd1 vccd1 vccd1 _7472_/X sky130_fd_sc_hd__xor2_2
X_6423_ _6484_/S _6401_/X _6422_/X vssd1 vssd1 vccd1 vccd1 _6423_/Y sky130_fd_sc_hd__o21ai_1
X_4684_ _4685_/A _4685_/C vssd1 vssd1 vccd1 vccd1 _4687_/B sky130_fd_sc_hd__and2_1
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6354_ _6354_/A _6492_/B _6431_/S vssd1 vssd1 vccd1 vccd1 _6354_/X sky130_fd_sc_hd__and3_1
XFILLER_103_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6285_ _4062_/B _4169_/Y _4180_/Y _4055_/B vssd1 vssd1 vccd1 vccd1 _6285_/X sky130_fd_sc_hd__o2bb2a_1
X_5305_ _5621_/A _5344_/B vssd1 vssd1 vccd1 vccd1 _5305_/Y sky130_fd_sc_hd__nor2_1
X_8024_ _8065_/CLK _8024_/D vssd1 vssd1 vccd1 vccd1 _8024_/Q sky130_fd_sc_hd__dfxtp_1
X_5236_ _5236_/A _5236_/B vssd1 vssd1 vccd1 vccd1 _5237_/B sky130_fd_sc_hd__nand2_1
XFILLER_75_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5167_ _6807_/A _5956_/A _5165_/X _5166_/X vssd1 vssd1 vccd1 vccd1 _5169_/B sky130_fd_sc_hd__a211o_1
X_4118_ _4063_/A _4116_/Y _4117_/Y _4078_/B vssd1 vssd1 vccd1 vccd1 _4118_/X sky130_fd_sc_hd__o31a_4
XFILLER_83_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5098_ _5098_/A _5098_/B vssd1 vssd1 vccd1 vccd1 _5100_/A sky130_fd_sc_hd__or2_4
X_4049_ _8059_/Q _4050_/B vssd1 vssd1 vccd1 vccd1 _4055_/B sky130_fd_sc_hd__xor2_4
XFILLER_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7808_ _6225_/S _6216_/X _7572_/X _7930_/A vssd1 vssd1 vccd1 vccd1 _7833_/C sky130_fd_sc_hd__a211o_4
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7739_ _7789_/A _7739_/B vssd1 vssd1 vccd1 vccd1 _7741_/A sky130_fd_sc_hd__nor2_1
XFILLER_12_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6026_/X _6042_/A _6044_/B vssd1 vssd1 vccd1 vccd1 _6071_/A sky130_fd_sc_hd__a21oi_4
XFILLER_85_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5021_ _5022_/A _5022_/B vssd1 vssd1 vccd1 vccd1 _5046_/A sky130_fd_sc_hd__nor2_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6972_ _6970_/A _6970_/B _7024_/A vssd1 vssd1 vccd1 vccd1 _6975_/B sky130_fd_sc_hd__a21bo_2
X_5923_ _5923_/A _5927_/B vssd1 vssd1 vccd1 vccd1 _5924_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5854_ _5797_/A _5855_/B _5369_/B _5889_/B vssd1 vssd1 vccd1 vccd1 _5868_/A sky130_fd_sc_hd__o211a_1
X_4805_ _4806_/A _4805_/B _4805_/C vssd1 vssd1 vccd1 vccd1 _4805_/X sky130_fd_sc_hd__and3_1
XFILLER_21_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7524_ _7538_/S _7524_/B vssd1 vssd1 vccd1 vccd1 _7525_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5785_ _5749_/X _5787_/A _5938_/B vssd1 vssd1 vccd1 vccd1 _5785_/X sky130_fd_sc_hd__o21a_2
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4736_ _4580_/X _4613_/X _4735_/B vssd1 vssd1 vccd1 vccd1 _4736_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7455_ _7452_/X _7454_/X _7455_/S vssd1 vssd1 vccd1 vccd1 _7455_/X sky130_fd_sc_hd__mux2_1
X_4667_ _4639_/A _4639_/B _4639_/C vssd1 vssd1 vccd1 vccd1 _4668_/C sky130_fd_sc_hd__a21o_1
X_6406_ _6407_/A _6407_/B vssd1 vssd1 vccd1 vccd1 _6406_/X sky130_fd_sc_hd__and2_1
X_7386_ _6938_/Y _7445_/B _6937_/A vssd1 vssd1 vccd1 vccd1 _7447_/B sky130_fd_sc_hd__a21oi_1
X_6337_ _6050_/Y _6047_/X _6767_/S vssd1 vssd1 vccd1 vccd1 _6338_/C sky130_fd_sc_hd__mux2_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4598_ _4563_/B _4563_/C _4563_/A vssd1 vssd1 vccd1 vccd1 _4599_/C sky130_fd_sc_hd__a21o_2
XFILLER_103_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6268_ _8009_/Q _6354_/A _8010_/Q vssd1 vssd1 vccd1 vccd1 _6268_/X sky130_fd_sc_hd__and3b_4
X_8007_ _6770_/A _8026_/Q _8007_/S vssd1 vssd1 vccd1 vccd1 _8082_/D sky130_fd_sc_hd__mux2_1
X_6199_ _6140_/Y _6121_/Y _6199_/S vssd1 vssd1 vccd1 vccd1 _6199_/X sky130_fd_sc_hd__mux2_2
X_5219_ _5212_/A _5212_/B _5213_/X vssd1 vssd1 vccd1 vccd1 _5239_/A sky130_fd_sc_hd__a21o_2
XFILLER_28_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5570_ _5570_/A _5570_/B vssd1 vssd1 vccd1 vccd1 _5635_/A sky130_fd_sc_hd__nor2_4
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4521_ _4521_/A _4521_/B vssd1 vssd1 vccd1 vccd1 _4546_/B sky130_fd_sc_hd__xnor2_2
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4452_ _4451_/B _4451_/C _4451_/A vssd1 vssd1 vccd1 vccd1 _4453_/C sky130_fd_sc_hd__a21o_1
X_7240_ _7240_/A _7240_/B vssd1 vssd1 vccd1 vccd1 _7268_/A sky130_fd_sc_hd__xnor2_4
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7171_ _7173_/A _7173_/B vssd1 vssd1 vccd1 vccd1 _7171_/X sky130_fd_sc_hd__and2_1
X_4383_ _6916_/A _4374_/X _4380_/X _4382_/X vssd1 vssd1 vccd1 vccd1 _4383_/X sky130_fd_sc_hd__a22o_2
XFILLER_112_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _6118_/A _6118_/B _5610_/Y vssd1 vssd1 vccd1 vccd1 _6123_/B sky130_fd_sc_hd__o21ai_1
XFILLER_112_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6053_ _6054_/A _6054_/B vssd1 vssd1 vccd1 vccd1 _6055_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5004_ _5005_/A _5005_/B vssd1 vssd1 vccd1 vccd1 _5004_/Y sky130_fd_sc_hd__nor2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6955_ _7068_/A _7269_/B _7006_/B vssd1 vssd1 vccd1 vccd1 _6957_/C sky130_fd_sc_hd__and3_1
X_5906_ _5917_/A _5922_/A vssd1 vssd1 vccd1 vccd1 _5918_/A sky130_fd_sc_hd__and2_1
X_6886_ _6896_/B _6896_/A vssd1 vssd1 vccd1 vccd1 _6888_/B sky130_fd_sc_hd__nand2b_2
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5837_ _5837_/A _5837_/B vssd1 vssd1 vccd1 vccd1 _5838_/B sky130_fd_sc_hd__nand2_2
X_5768_ _5800_/A _5796_/B vssd1 vssd1 vccd1 vccd1 _5768_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7507_ _7496_/X _7506_/X _7515_/S vssd1 vssd1 vccd1 vccd1 _7531_/C sky130_fd_sc_hd__mux2_1
X_4719_ _4726_/A _4726_/B vssd1 vssd1 vccd1 vccd1 _4720_/C sky130_fd_sc_hd__and2_1
X_7438_ _7438_/A _7438_/B vssd1 vssd1 vccd1 vccd1 _7483_/S sky130_fd_sc_hd__or2_4
X_5699_ _5692_/B _5691_/B _5695_/B _5693_/X vssd1 vssd1 vccd1 vccd1 _5743_/A sky130_fd_sc_hd__a31o_4
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7369_ _7369_/A _7369_/B vssd1 vssd1 vccd1 vccd1 _7370_/B sky130_fd_sc_hd__or2_1
XFILLER_103_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6740_ _6713_/S _6655_/Y _6691_/Y _6652_/Y vssd1 vssd1 vccd1 vccd1 _6740_/X sky130_fd_sc_hd__a22o_1
XFILLER_63_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6671_ _6645_/Y _6669_/A _6713_/S vssd1 vssd1 vccd1 vccd1 _6672_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5622_ _6971_/B _5755_/A vssd1 vssd1 vccd1 vccd1 _5663_/A sky130_fd_sc_hd__nor2_1
X_5553_ _5548_/A _5548_/B _5546_/Y vssd1 vssd1 vccd1 vccd1 _5607_/A sky130_fd_sc_hd__o21ai_2
XFILLER_117_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4504_ _4505_/A _4505_/B vssd1 vssd1 vccd1 vccd1 _4504_/Y sky130_fd_sc_hd__nand2b_1
X_5484_ _5485_/A _5485_/B vssd1 vssd1 vccd1 vccd1 _5484_/Y sky130_fd_sc_hd__nor2_2
XFILLER_117_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4435_ _4988_/A vssd1 vssd1 vccd1 vccd1 _5020_/A sky130_fd_sc_hd__inv_6
X_7223_ _7229_/B _7229_/A vssd1 vssd1 vccd1 vccd1 _7223_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_116_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4366_ _4412_/A _4407_/B _7085_/A _4602_/A vssd1 vssd1 vccd1 vccd1 _4366_/X sky130_fd_sc_hd__a211o_1
X_7154_ _7154_/A _7154_/B vssd1 vssd1 vccd1 vccd1 _7155_/B sky130_fd_sc_hd__and2_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6105_ _6099_/A _6099_/B _6110_/A _6093_/B _6132_/B vssd1 vssd1 vccd1 vccd1 _6192_/C
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4297_ _4074_/Y _4118_/X _4059_/B _4071_/Y vssd1 vssd1 vccd1 vccd1 _4297_/X sky130_fd_sc_hd__o211a_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7085_ _7085_/A _7085_/B vssd1 vssd1 vccd1 vccd1 _7086_/B sky130_fd_sc_hd__nand2_1
X_6036_ _6038_/B _6037_/B vssd1 vssd1 vccd1 vccd1 _6039_/A sky130_fd_sc_hd__nor2_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7987_ _8023_/Q _8063_/Q _7990_/S vssd1 vssd1 vccd1 vccd1 _8063_/D sky130_fd_sc_hd__mux2_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6938_ _7445_/A vssd1 vssd1 vccd1 vccd1 _6938_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6869_ _7027_/A _6842_/B _6842_/C vssd1 vssd1 vccd1 vccd1 _6870_/B sky130_fd_sc_hd__o21ai_1
XFILLER_22_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4220_ _4209_/X _4217_/Y _4218_/Y _4230_/C vssd1 vssd1 vccd1 vccd1 _4244_/A sky130_fd_sc_hd__a211o_2
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4151_ _4175_/B _4147_/B _4147_/C _4168_/B1 vssd1 vssd1 vccd1 vccd1 _4152_/B sky130_fd_sc_hd__o31a_2
XFILLER_68_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4082_ _4088_/A _8052_/Q _4096_/A vssd1 vssd1 vccd1 vccd1 _4083_/B sky130_fd_sc_hd__o21ai_4
XFILLER_83_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7910_ _7887_/A _7887_/B _7910_/C _7910_/D vssd1 vssd1 vccd1 vccd1 _7911_/B sky130_fd_sc_hd__and4bb_2
X_7841_ _6636_/Y _7617_/A _7823_/A _7773_/X vssd1 vssd1 vccd1 vccd1 _7842_/B sky130_fd_sc_hd__a31o_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7772_ _7765_/X _7795_/B _7771_/Y vssd1 vssd1 vccd1 vccd1 _7772_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4984_ _4984_/A _4984_/B _4984_/C vssd1 vssd1 vccd1 vccd1 _5018_/A sky130_fd_sc_hd__nand3_1
X_6723_ _6616_/C _6616_/B _6733_/S vssd1 vssd1 vccd1 vccd1 _6723_/X sky130_fd_sc_hd__mux2_1
X_6654_ _6695_/S _6654_/B vssd1 vssd1 vccd1 vccd1 _6655_/B sky130_fd_sc_hd__or2_1
X_5605_ _5616_/A _5605_/B vssd1 vssd1 vccd1 vccd1 _5660_/B sky130_fd_sc_hd__nand2_1
X_6585_ _6521_/A _6524_/B _6709_/A vssd1 vssd1 vccd1 vccd1 _6585_/X sky130_fd_sc_hd__o21a_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5536_ _5537_/A _5537_/B vssd1 vssd1 vccd1 vccd1 _5536_/Y sky130_fd_sc_hd__nor2_1
X_5467_ _5467_/A _5467_/B vssd1 vssd1 vccd1 vccd1 _5468_/B sky130_fd_sc_hd__nand2_2
X_7206_ _7281_/A _7281_/C vssd1 vssd1 vccd1 vccd1 _7206_/Y sky130_fd_sc_hd__nand2_1
X_4418_ _4412_/A _4412_/B _4377_/A vssd1 vssd1 vccd1 vccd1 _4418_/X sky130_fd_sc_hd__a21o_1
X_5398_ _5399_/A _5399_/B vssd1 vssd1 vccd1 vccd1 _5398_/X sky130_fd_sc_hd__and2_1
XFILLER_113_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7137_ _7025_/Y _7187_/A _7087_/B vssd1 vssd1 vccd1 vccd1 _7182_/A sky130_fd_sc_hd__o21a_2
X_4349_ _4430_/B _4430_/C _4430_/A vssd1 vssd1 vccd1 vccd1 _4349_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7068_ _7068_/A _7306_/B vssd1 vssd1 vccd1 vccd1 _7127_/B sky130_fd_sc_hd__nand2_2
XFILLER_100_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6019_ _6021_/A0 _6018_/B _6030_/B vssd1 vssd1 vccd1 vccd1 _6020_/A sky130_fd_sc_hd__o21a_2
XFILLER_74_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6370_ _6492_/B _6353_/Y _6451_/A _6369_/Y vssd1 vssd1 vccd1 vccd1 _6371_/B sky130_fd_sc_hd__o22a_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5321_ _5325_/A _5325_/B vssd1 vssd1 vccd1 vccd1 _5321_/X sky130_fd_sc_hd__or2_1
XFILLER_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8040_ _8065_/CLK _8040_/D vssd1 vssd1 vccd1 vccd1 _8040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5252_ _5745_/A _5722_/A _5722_/B _5723_/A _6951_/D vssd1 vssd1 vccd1 vccd1 _5252_/X
+ sky130_fd_sc_hd__a32o_1
X_4203_ _8069_/Q _4204_/B vssd1 vssd1 vccd1 vccd1 _4216_/C sky130_fd_sc_hd__xor2_4
XFILLER_68_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5183_ _5183_/A _5183_/B vssd1 vssd1 vccd1 vccd1 _5215_/A sky130_fd_sc_hd__nand2_4
XFILLER_110_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4134_ _4303_/B _4133_/X _4131_/X vssd1 vssd1 vccd1 vccd1 _5066_/B sky130_fd_sc_hd__a21o_1
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4065_ _4081_/A vssd1 vssd1 vccd1 vccd1 _4080_/C sky130_fd_sc_hd__clkinv_2
XFILLER_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7824_ _7649_/A _7793_/Y _7823_/Y vssd1 vssd1 vccd1 vccd1 _7824_/Y sky130_fd_sc_hd__o21ai_2
X_7755_ _7755_/A _7831_/A vssd1 vssd1 vccd1 vccd1 _7908_/A sky130_fd_sc_hd__nor2_8
X_4967_ _5090_/A _5033_/B vssd1 vssd1 vccd1 vccd1 _4968_/B sky130_fd_sc_hd__or2_4
X_6706_ _6706_/A vssd1 vssd1 vccd1 vccd1 _6707_/B sky130_fd_sc_hd__inv_2
X_7686_ _7544_/B _7889_/B _7889_/A vssd1 vssd1 vccd1 vccd1 _7687_/C sky130_fd_sc_hd__mux2_2
X_4898_ _4874_/A _4947_/C _4892_/A _4892_/B vssd1 vssd1 vccd1 vccd1 _4900_/A sky130_fd_sc_hd__o2bb2a_4
XFILLER_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6637_ _6753_/S _6749_/S vssd1 vssd1 vccd1 vccd1 _6638_/A sky130_fd_sc_hd__or2_2
X_6568_ _6530_/Y _6539_/C _6525_/B vssd1 vssd1 vccd1 vccd1 _6568_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_22_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5519_ _5672_/A _6971_/B vssd1 vssd1 vccd1 vccd1 _5521_/B sky130_fd_sc_hd__nor2_4
X_6499_ _6549_/A _6548_/B vssd1 vssd1 vccd1 vccd1 _6550_/D sky130_fd_sc_hd__nor2_2
Xfanout131 _4111_/X vssd1 vssd1 vccd1 vccd1 _6021_/A0 sky130_fd_sc_hd__buf_2
Xfanout120 _4350_/X vssd1 vssd1 vccd1 vccd1 _4456_/B sky130_fd_sc_hd__buf_4
Xfanout153 _7068_/A vssd1 vssd1 vccd1 vccd1 _7123_/A sky130_fd_sc_hd__clkbuf_16
Xfanout142 _7057_/A vssd1 vssd1 vccd1 vccd1 _7116_/A sky130_fd_sc_hd__buf_8
Xfanout164 _7027_/A vssd1 vssd1 vccd1 vccd1 _4360_/A sky130_fd_sc_hd__buf_6
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout197 _5107_/X vssd1 vssd1 vccd1 vccd1 _6951_/D sky130_fd_sc_hd__clkbuf_16
Xfanout186 _4260_/C vssd1 vssd1 vccd1 vccd1 _4259_/B sky130_fd_sc_hd__buf_4
XFILLER_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout175 _7311_/A vssd1 vssd1 vccd1 vccd1 _7214_/A sky130_fd_sc_hd__buf_8
XFILLER_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5870_ _6873_/B _5927_/B vssd1 vssd1 vccd1 vccd1 _5877_/A sky130_fd_sc_hd__nand2_1
X_4821_ _4820_/S _4798_/A _4926_/A vssd1 vssd1 vccd1 vccd1 _4894_/A sky130_fd_sc_hd__a21o_2
X_7540_ _7766_/B _7797_/B _7539_/X vssd1 vssd1 vccd1 vccd1 _7554_/B sky130_fd_sc_hd__o21ai_4
X_4752_ _4757_/B vssd1 vssd1 vccd1 vccd1 _4752_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4683_ _4665_/A _4665_/B _4665_/C vssd1 vssd1 vccd1 vccd1 _4685_/C sky130_fd_sc_hd__a21o_1
X_7471_ _7471_/A _7471_/B vssd1 vssd1 vccd1 vccd1 _7471_/X sky130_fd_sc_hd__xor2_2
X_6422_ _6451_/A _6422_/B vssd1 vssd1 vccd1 vccd1 _6422_/X sky130_fd_sc_hd__or2_1
X_6353_ _6354_/A _6431_/S vssd1 vssd1 vccd1 vccd1 _6353_/Y sky130_fd_sc_hd__nand2_1
X_6284_ _4053_/Y _4178_/X _4180_/Y _4055_/B _6283_/X vssd1 vssd1 vccd1 vccd1 _6284_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5304_ _5666_/A _5432_/A vssd1 vssd1 vccd1 vccd1 _5306_/S sky130_fd_sc_hd__nand2_2
XFILLER_115_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8023_ _8077_/CLK _8023_/D vssd1 vssd1 vccd1 vccd1 _8023_/Q sky130_fd_sc_hd__dfxtp_1
X_5235_ _5236_/A _5236_/B vssd1 vssd1 vccd1 vccd1 _5961_/A sky130_fd_sc_hd__or2_2
X_5166_ _5541_/A _5166_/B _5166_/C vssd1 vssd1 vccd1 vccd1 _5166_/X sky130_fd_sc_hd__and3_1
XFILLER_68_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4117_ _4117_/A _4117_/B _4117_/C vssd1 vssd1 vccd1 vccd1 _4117_/Y sky130_fd_sc_hd__nor3_4
XFILLER_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5097_ _5098_/B vssd1 vssd1 vccd1 vccd1 _5097_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4048_ _4096_/A _4080_/B vssd1 vssd1 vccd1 vccd1 _4050_/B sky130_fd_sc_hd__nand2_4
XFILLER_44_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7807_ _7759_/Y _7760_/X _7787_/B _7728_/A vssd1 vssd1 vccd1 vccd1 _7887_/A sky130_fd_sc_hd__o31a_4
X_5999_ _6000_/A _6000_/B vssd1 vssd1 vccd1 vccd1 _6320_/A sky130_fd_sc_hd__nor2_4
XFILLER_52_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7738_ _7738_/A _7738_/B vssd1 vssd1 vccd1 vccd1 _7739_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7669_ _7831_/A _6226_/X _7668_/X vssd1 vssd1 vccd1 vccd1 _7731_/A sky130_fd_sc_hd__a21oi_4
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5020_/A _5020_/B vssd1 vssd1 vccd1 vccd1 _5022_/B sky130_fd_sc_hd__nand2_4
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6971_ _7027_/A _6971_/B _6970_/X vssd1 vssd1 vccd1 vccd1 _7024_/A sky130_fd_sc_hd__or3b_1
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5922_ _5922_/A _5922_/B vssd1 vssd1 vccd1 vccd1 _5924_/A sky130_fd_sc_hd__or2_1
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5853_ _5925_/A _5853_/B vssd1 vssd1 vccd1 vccd1 _5921_/A sky130_fd_sc_hd__nor2_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4804_ _4806_/A _4806_/B vssd1 vssd1 vccd1 vccd1 _4804_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_34_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5784_ _5786_/A _5786_/B vssd1 vssd1 vccd1 vccd1 _5787_/A sky130_fd_sc_hd__nor2_8
X_7523_ _7513_/S _7512_/Y _7517_/Y _7522_/X vssd1 vssd1 vccd1 vccd1 _7523_/X sky130_fd_sc_hd__a211o_1
X_4735_ _4580_/X _4735_/B vssd1 vssd1 vccd1 vccd1 _4848_/B sky130_fd_sc_hd__and2b_2
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7454_ _7454_/A _7454_/B vssd1 vssd1 vccd1 vccd1 _7454_/X sky130_fd_sc_hd__or2_1
X_4666_ _4665_/B _4665_/C _4665_/A vssd1 vssd1 vccd1 vccd1 _4668_/B sky130_fd_sc_hd__a21bo_1
X_6405_ _7057_/A _6839_/B _6445_/S vssd1 vssd1 vccd1 vccd1 _6407_/B sky130_fd_sc_hd__mux2_2
X_7385_ _7442_/A _7442_/B _6989_/X vssd1 vssd1 vccd1 vccd1 _7445_/B sky130_fd_sc_hd__o21bai_2
X_4597_ _4596_/A _4596_/B _4596_/C _4588_/X vssd1 vssd1 vccd1 vccd1 _4599_/B sky130_fd_sc_hd__a31o_2
X_6336_ _6336_/A _6336_/B vssd1 vssd1 vccd1 vccd1 _6338_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6267_ _7611_/D _6267_/B _7568_/B vssd1 vssd1 vccd1 vccd1 _6267_/X sky130_fd_sc_hd__and3_1
X_8006_ _8081_/Q _8025_/Q _8007_/S vssd1 vssd1 vccd1 vccd1 _8081_/D sky130_fd_sc_hd__mux2_1
X_6198_ _6225_/S _6196_/X _6197_/X vssd1 vssd1 vccd1 vccd1 _6255_/A sky130_fd_sc_hd__o21ai_2
X_5218_ _5220_/A _5220_/B vssd1 vssd1 vccd1 vccd1 _5218_/Y sky130_fd_sc_hd__nor2_1
X_5149_ _5207_/A _5715_/A vssd1 vssd1 vccd1 vccd1 _6783_/A sky130_fd_sc_hd__nor2_4
XFILLER_28_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4520_ _7247_/A _4496_/B _4494_/X vssd1 vssd1 vccd1 vccd1 _4546_/A sky130_fd_sc_hd__o21ai_4
X_4451_ _4451_/A _4451_/B _4451_/C vssd1 vssd1 vccd1 vccd1 _4453_/B sky130_fd_sc_hd__nand3_2
X_7170_ _7213_/A _7170_/B _7213_/B vssd1 vssd1 vccd1 vccd1 _7173_/B sky130_fd_sc_hd__and3_2
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6121_ _7358_/B _6174_/A _6177_/A _6115_/X _6120_/X vssd1 vssd1 vccd1 vccd1 _6121_/Y
+ sky130_fd_sc_hd__a221oi_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4382_ _4348_/X _4365_/Y _4429_/B _4494_/A vssd1 vssd1 vccd1 vccd1 _4382_/X sky130_fd_sc_hd__o31a_1
XFILLER_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6052_ _6054_/A _6054_/B vssd1 vssd1 vccd1 vccd1 _6067_/A sky130_fd_sc_hd__and2b_1
XFILLER_58_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5003_/A _5003_/B vssd1 vssd1 vccd1 vccd1 _5005_/B sky130_fd_sc_hd__xnor2_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6954_ _6957_/B _6954_/B vssd1 vssd1 vccd1 vccd1 _7006_/B sky130_fd_sc_hd__nor2_4
XFILLER_81_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5905_ _5921_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _5922_/A sky130_fd_sc_hd__and2_1
X_6885_ _6857_/C _6882_/Y _6897_/B _6947_/C vssd1 vssd1 vccd1 vccd1 _6896_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5836_ _5836_/A _5836_/B vssd1 vssd1 vccd1 vccd1 _5837_/B sky130_fd_sc_hd__or2_1
X_5767_ _5767_/A _5767_/B vssd1 vssd1 vccd1 vccd1 _5804_/A sky130_fd_sc_hd__xor2_4
XFILLER_108_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7506_ _7490_/X _7473_/X _7527_/S vssd1 vssd1 vccd1 vccd1 _7506_/X sky130_fd_sc_hd__mux2_1
X_4718_ _7281_/A _5034_/A _4718_/C vssd1 vssd1 vccd1 vccd1 _4726_/B sky130_fd_sc_hd__and3_1
X_5698_ _5700_/B _5700_/A vssd1 vssd1 vccd1 vccd1 _5698_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_107_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7437_ _7438_/B _7524_/B vssd1 vssd1 vccd1 vccd1 _7437_/Y sky130_fd_sc_hd__nor2_1
X_4649_ _4648_/B _4648_/C _4648_/A vssd1 vssd1 vccd1 vccd1 _4650_/C sky130_fd_sc_hd__a21o_1
XFILLER_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7368_ _7370_/A _7369_/B vssd1 vssd1 vccd1 vccd1 _7516_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6319_ _7400_/A _6322_/B _6577_/A _6006_/X vssd1 vssd1 vccd1 vccd1 _6320_/B sky130_fd_sc_hd__o2bb2ai_4
X_7299_ _7299_/A _7299_/B vssd1 vssd1 vccd1 vccd1 _7324_/A sky130_fd_sc_hd__nand2_1
XFILLER_103_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6670_ _6669_/Y _6662_/X _6713_/S vssd1 vssd1 vccd1 vccd1 _6670_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5621_ _5621_/A _5880_/A vssd1 vssd1 vccd1 vccd1 _5621_/Y sky130_fd_sc_hd__nor2_1
X_5552_ _5554_/B _5554_/A vssd1 vssd1 vccd1 vccd1 _5558_/A sky130_fd_sc_hd__nand2b_1
X_4503_ _4503_/A _4503_/B vssd1 vssd1 vccd1 vccd1 _4505_/B sky130_fd_sc_hd__xor2_4
X_5483_ _5471_/A _5471_/B _5461_/X vssd1 vssd1 vccd1 vccd1 _5485_/B sky130_fd_sc_hd__a21oi_2
XFILLER_104_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4434_ _4494_/A _4429_/X _4431_/X _4433_/X vssd1 vssd1 vccd1 vccd1 _4558_/B sky130_fd_sc_hd__a2bb2o_4
X_7222_ _7220_/A _7220_/B _7243_/A vssd1 vssd1 vccd1 vccd1 _7229_/B sky130_fd_sc_hd__o21ba_2
X_4365_ _4430_/B _4430_/C vssd1 vssd1 vccd1 vccd1 _4365_/Y sky130_fd_sc_hd__nor2_1
X_7153_ _7154_/A _7154_/B vssd1 vssd1 vccd1 vccd1 _7155_/A sky130_fd_sc_hd__nor2_1
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6104_ _6104_/A _6104_/B vssd1 vssd1 vccd1 vccd1 _6192_/B sky130_fd_sc_hd__xnor2_4
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7084_ _7084_/A _7084_/B vssd1 vssd1 vccd1 vccd1 _7087_/A sky130_fd_sc_hd__nand2_4
XFILLER_100_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6035_ _6035_/A0 _6034_/Y _6035_/S vssd1 vssd1 vccd1 vccd1 _6037_/B sky130_fd_sc_hd__mux2_4
X_4296_ _4296_/A _4296_/B vssd1 vssd1 vccd1 vccd1 _4296_/Y sky130_fd_sc_hd__nand2_4
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7986_ _8022_/Q _8062_/Q _7986_/S vssd1 vssd1 vccd1 vccd1 _8062_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6937_ _6937_/A _6937_/B vssd1 vssd1 vccd1 vccd1 _7445_/A sky130_fd_sc_hd__or2_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6868_ _6884_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _6881_/A sky130_fd_sc_hd__xnor2_4
X_5819_ _5919_/A _5858_/B vssd1 vssd1 vccd1 vccd1 _5821_/B sky130_fd_sc_hd__nand2_1
X_6799_ _6804_/A _6799_/B vssd1 vssd1 vccd1 vccd1 _6800_/C sky130_fd_sc_hd__nand2_1
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4150_ _6326_/B vssd1 vssd1 vccd1 vccd1 _6272_/B sky130_fd_sc_hd__inv_6
XFILLER_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4081_ _4081_/A _4081_/B _4080_/B vssd1 vssd1 vccd1 vccd1 _4081_/X sky130_fd_sc_hd__or3b_4
XFILLER_68_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7840_ _6636_/Y _7617_/A _7823_/A vssd1 vssd1 vccd1 vccd1 _7895_/A sky130_fd_sc_hd__a21oi_2
XFILLER_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7771_ _7765_/X _7795_/B _7802_/B2 vssd1 vssd1 vccd1 vccd1 _7771_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4983_ _5013_/A _5013_/C _5034_/A _4947_/C vssd1 vssd1 vccd1 vccd1 _4984_/C sky130_fd_sc_hd__a2bb2o_2
XFILLER_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6722_ _6721_/X _6616_/D _6733_/S vssd1 vssd1 vccd1 vccd1 _6722_/X sky130_fd_sc_hd__mux2_1
X_6653_ _6713_/S _6645_/Y _6651_/Y _6652_/Y vssd1 vssd1 vccd1 vccd1 _6653_/X sky130_fd_sc_hd__a22o_1
X_5604_ _5604_/A _5604_/B vssd1 vssd1 vccd1 vccd1 _5605_/B sky130_fd_sc_hd__nand2_1
X_6584_ _6584_/A _6584_/B vssd1 vssd1 vccd1 vccd1 _6584_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_11_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5535_ _5537_/A _5537_/B vssd1 vssd1 vccd1 vccd1 _5535_/Y sky130_fd_sc_hd__nand2_1
X_5466_ _5466_/A _5466_/B vssd1 vssd1 vccd1 vccd1 _5467_/B sky130_fd_sc_hd__nor2_2
XFILLER_117_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4417_ _4483_/A _7311_/A _4441_/A vssd1 vssd1 vccd1 vccd1 _4472_/B sky130_fd_sc_hd__mux2_2
X_7205_ _7205_/A _7205_/B vssd1 vssd1 vccd1 vccd1 _7220_/A sky130_fd_sc_hd__xnor2_2
X_5397_ _5298_/A _5298_/B _5347_/B _5358_/A _5358_/B vssd1 vssd1 vccd1 vccd1 _5414_/A
+ sky130_fd_sc_hd__a32oi_4
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7136_ _7136_/A _7210_/B vssd1 vssd1 vccd1 vccd1 _7187_/A sky130_fd_sc_hd__nor2_2
X_4348_ _4430_/B _4430_/C vssd1 vssd1 vccd1 vccd1 _4348_/X sky130_fd_sc_hd__and2_1
XFILLER_100_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4279_ _4354_/A _4483_/A _4275_/X _6035_/A0 _4278_/Y vssd1 vssd1 vccd1 vccd1 _6315_/A
+ sky130_fd_sc_hd__a221oi_4
XFILLER_59_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7067_ _7067_/A _7067_/B vssd1 vssd1 vccd1 vccd1 _7127_/A sky130_fd_sc_hd__xor2_4
XFILLER_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6018_ _6018_/A _6018_/B vssd1 vssd1 vccd1 vccd1 _6030_/B sky130_fd_sc_hd__nand2_4
XFILLER_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7969_ _8048_/Q _7970_/C _8049_/Q vssd1 vssd1 vccd1 vccd1 _7971_/C sky130_fd_sc_hd__a21o_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5320_ _5352_/A _5352_/B _7319_/B vssd1 vssd1 vccd1 vccd1 _5325_/B sky130_fd_sc_hd__nand3_4
X_5251_ _5367_/A _5672_/A vssd1 vssd1 vccd1 vccd1 _5431_/A sky130_fd_sc_hd__or2_2
X_4202_ _6278_/B _4200_/Y _4201_/X _4193_/B _4193_/A vssd1 vssd1 vccd1 vccd1 _4227_/S
+ sky130_fd_sc_hd__a2111o_4
X_5182_ _5182_/A _5182_/B _5182_/C vssd1 vssd1 vccd1 vccd1 _5183_/B sky130_fd_sc_hd__or3_2
X_4133_ _6274_/A _5993_/B _4132_/X vssd1 vssd1 vccd1 vccd1 _4133_/X sky130_fd_sc_hd__a21o_1
XFILLER_68_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4064_ _4064_/A _4064_/B vssd1 vssd1 vccd1 vccd1 _4081_/A sky130_fd_sc_hd__nand2_4
XFILLER_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7823_ _7823_/A _7823_/B vssd1 vssd1 vccd1 vccd1 _7823_/Y sky130_fd_sc_hd__nand2_2
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7754_ _7928_/A _7754_/B vssd1 vssd1 vccd1 vccd1 _8034_/D sky130_fd_sc_hd__nor2_1
XFILLER_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6705_ _6733_/S _6670_/X _6704_/Y vssd1 vssd1 vccd1 vccd1 _6706_/A sky130_fd_sc_hd__o21a_1
X_4966_ _4959_/A _4959_/B _4956_/X vssd1 vssd1 vccd1 vccd1 _4968_/A sky130_fd_sc_hd__o21a_4
X_7685_ _7657_/B _7504_/X _7657_/Y vssd1 vssd1 vccd1 vccd1 _7889_/B sky130_fd_sc_hd__o21a_2
X_4897_ _4897_/A _4897_/B vssd1 vssd1 vccd1 vccd1 _5034_/B sky130_fd_sc_hd__and2_4
X_6636_ _7894_/A vssd1 vssd1 vccd1 vccd1 _6636_/Y sky130_fd_sc_hd__clkinv_2
X_6567_ _6578_/A _6567_/B vssd1 vssd1 vccd1 vccd1 _6605_/A sky130_fd_sc_hd__xnor2_1
XFILLER_22_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5518_ _5518_/A _5518_/B vssd1 vssd1 vccd1 vccd1 _5521_/A sky130_fd_sc_hd__xnor2_4
X_6498_ _6571_/B _6572_/A _6570_/A vssd1 vssd1 vccd1 vccd1 _6548_/B sky130_fd_sc_hd__nand3b_4
X_5449_ _5449_/A _5449_/B vssd1 vssd1 vccd1 vccd1 _5450_/B sky130_fd_sc_hd__xnor2_4
XFILLER_59_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout121 _7284_/A vssd1 vssd1 vccd1 vccd1 _4654_/A sky130_fd_sc_hd__buf_8
Xfanout110 _5316_/Y vssd1 vssd1 vccd1 vccd1 _5797_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout132 _4110_/Y vssd1 vssd1 vccd1 vccd1 _4303_/B sky130_fd_sc_hd__clkbuf_8
Xfanout143 _4340_/Y vssd1 vssd1 vccd1 vccd1 _7057_/A sky130_fd_sc_hd__buf_6
Xfanout154 _4501_/A vssd1 vssd1 vccd1 vccd1 _4430_/A sky130_fd_sc_hd__buf_4
Xfanout165 _4325_/Y vssd1 vssd1 vccd1 vccd1 _7027_/A sky130_fd_sc_hd__clkbuf_16
X_7119_ _7119_/A _7119_/B vssd1 vssd1 vccd1 vccd1 _7120_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout187 _4234_/X vssd1 vssd1 vccd1 vccd1 _4260_/C sky130_fd_sc_hd__buf_4
Xfanout198 _6800_/B vssd1 vssd1 vccd1 vccd1 _7046_/B sky130_fd_sc_hd__buf_8
Xfanout176 _4342_/X vssd1 vssd1 vccd1 vccd1 _7311_/A sky130_fd_sc_hd__buf_8
XFILLER_103_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4820_ _4923_/B _4923_/C _4820_/S vssd1 vssd1 vccd1 vccd1 _4927_/A sky130_fd_sc_hd__mux2_8
XFILLER_33_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4773_/A _4988_/A _4751_/C _4991_/A vssd1 vssd1 vccd1 vccd1 _4757_/B sky130_fd_sc_hd__or4b_4
XFILLER_119_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7470_ _7537_/C vssd1 vssd1 vccd1 vccd1 _7470_/Y sky130_fd_sc_hd__inv_2
X_4682_ _4714_/A _4714_/B vssd1 vssd1 vccd1 vccd1 _4727_/A sky130_fd_sc_hd__and2_2
X_6421_ _6408_/X _6420_/X _6431_/S vssd1 vssd1 vccd1 vccd1 _6422_/B sky130_fd_sc_hd__mux2_1
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6352_ _6359_/A _7402_/A vssd1 vssd1 vccd1 vccd1 _6483_/A sky130_fd_sc_hd__and2_2
XFILLER_115_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6283_ _4053_/Y _4178_/X _6274_/Y _6282_/Y vssd1 vssd1 vccd1 vccd1 _6283_/X sky130_fd_sc_hd__o22a_1
X_5303_ _6800_/B _5880_/A vssd1 vssd1 vccd1 vccd1 _5303_/Y sky130_fd_sc_hd__nor2_4
X_8022_ _8063_/CLK _8022_/D vssd1 vssd1 vccd1 vccd1 _8022_/Q sky130_fd_sc_hd__dfxtp_1
X_5234_ _5179_/A _5179_/B _5177_/X vssd1 vssd1 vccd1 vccd1 _5236_/B sky130_fd_sc_hd__a21oi_1
X_5165_ _5956_/A _5165_/B _5166_/C vssd1 vssd1 vccd1 vccd1 _5165_/X sky130_fd_sc_hd__and3b_1
X_4116_ _4095_/A _4115_/Y _4081_/A vssd1 vssd1 vccd1 vccd1 _4116_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5096_ _5095_/A _5095_/B _5095_/C vssd1 vssd1 vccd1 vccd1 _5098_/B sky130_fd_sc_hd__a21oi_2
X_4047_ _6272_/A vssd1 vssd1 vccd1 vccd1 _6060_/A sky130_fd_sc_hd__clkinv_8
XFILLER_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7806_ _7856_/A _7806_/B vssd1 vssd1 vccd1 vccd1 _8036_/D sky130_fd_sc_hd__nor2_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _6017_/B _6027_/A vssd1 vssd1 vccd1 vccd1 _6000_/B sky130_fd_sc_hd__nor2_4
XFILLER_33_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7737_ _7738_/A _7738_/B vssd1 vssd1 vccd1 vccd1 _7789_/A sky130_fd_sc_hd__and2_1
X_4949_ _4949_/A _4949_/B vssd1 vssd1 vccd1 vccd1 _4986_/B sky130_fd_sc_hd__xnor2_4
X_7668_ _7639_/B _6170_/X _7639_/Y _7784_/A vssd1 vssd1 vccd1 vccd1 _7668_/X sky130_fd_sc_hd__o211a_1
XFILLER_20_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6619_ _6621_/B vssd1 vssd1 vccd1 vccd1 _6619_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7599_ _7939_/A _7623_/A _7623_/B vssd1 vssd1 vccd1 vccd1 _7600_/C sky130_fd_sc_hd__a21oi_1
XFILLER_118_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6970_ _6970_/A _6970_/B vssd1 vssd1 vccd1 vccd1 _6970_/X sky130_fd_sc_hd__xor2_1
XFILLER_80_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5921_ _5921_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _5922_/B sky130_fd_sc_hd__nor2_1
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5852_ _5834_/A _5834_/B _5834_/C vssd1 vssd1 vccd1 vccd1 _5866_/B sky130_fd_sc_hd__a21oi_2
X_4803_ _4851_/A _4818_/B _4805_/B vssd1 vssd1 vccd1 vccd1 _4806_/B sky130_fd_sc_hd__a21bo_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5783_ _5781_/A _5781_/B _5782_/X vssd1 vssd1 vccd1 vccd1 _5786_/B sky130_fd_sc_hd__a21oi_4
X_7522_ _7516_/C _7518_/Y _7521_/Y vssd1 vssd1 vccd1 vccd1 _7522_/X sky130_fd_sc_hd__a21o_1
X_4734_ _4846_/A _4846_/B _4613_/X vssd1 vssd1 vccd1 vccd1 _4848_/A sky130_fd_sc_hd__a21oi_4
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7453_ _7448_/Y _7452_/X _7479_/S vssd1 vssd1 vccd1 vccd1 _7453_/X sky130_fd_sc_hd__mux2_1
X_4665_ _4665_/A _4665_/B _4665_/C vssd1 vssd1 vccd1 vccd1 _4685_/A sky130_fd_sc_hd__nand3_1
X_6404_ _6443_/A _6404_/B vssd1 vssd1 vccd1 vccd1 _6407_/A sky130_fd_sc_hd__nand2_1
X_7384_ _7440_/A _7440_/B _7049_/A vssd1 vssd1 vccd1 vccd1 _7442_/B sky130_fd_sc_hd__a21oi_2
X_4596_ _4596_/A _4596_/B _4596_/C vssd1 vssd1 vccd1 vccd1 _4646_/C sky130_fd_sc_hd__nand3_2
XFILLER_115_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6335_ _6308_/A _6334_/Y _6343_/B _7416_/A vssd1 vssd1 vccd1 vccd1 _6341_/B sky130_fd_sc_hd__a2bb2o_2
XFILLER_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6266_ _7831_/A _6264_/X _6265_/X vssd1 vssd1 vccd1 vccd1 _7568_/B sky130_fd_sc_hd__o21a_1
X_8005_ _8080_/Q _8024_/Q _8007_/S vssd1 vssd1 vccd1 vccd1 _8080_/D sky130_fd_sc_hd__mux2_1
X_6197_ _6112_/X _6190_/X _6193_/X _6226_/S vssd1 vssd1 vccd1 vccd1 _6197_/X sky130_fd_sc_hd__a211o_1
XFILLER_69_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5217_ _5215_/A _5215_/B _5216_/Y vssd1 vssd1 vccd1 vccd1 _5220_/B sky130_fd_sc_hd__o21a_2
XFILLER_57_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5148_ _5386_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _5465_/A sky130_fd_sc_hd__or2_2
XFILLER_28_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5079_ _5174_/A _5200_/A vssd1 vssd1 vccd1 vccd1 _5182_/A sky130_fd_sc_hd__and2b_2
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4450_ _4455_/A _5040_/A _4448_/Y vssd1 vssd1 vccd1 vccd1 _4451_/C sky130_fd_sc_hd__a21o_2
XFILLER_116_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4381_ _4602_/A _4407_/B _7136_/A vssd1 vssd1 vccd1 vccd1 _4429_/B sky130_fd_sc_hd__a21o_1
X_6120_ _6242_/S _6120_/B vssd1 vssd1 vccd1 vccd1 _6120_/X sky130_fd_sc_hd__and2b_1
XFILLER_86_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6051_ _4080_/X _6050_/Y _6051_/S vssd1 vssd1 vccd1 vccd1 _6054_/B sky130_fd_sc_hd__mux2_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5002_ _5010_/A _5010_/B _4996_/Y vssd1 vssd1 vccd1 vccd1 _5005_/A sky130_fd_sc_hd__a21boi_4
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6953_ _6902_/A _7150_/B _7046_/B _7284_/A vssd1 vssd1 vccd1 vccd1 _6954_/B sky130_fd_sc_hd__o22a_1
Xclkbuf_3_5__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _8057_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6884_ _6884_/A _6884_/B vssd1 vssd1 vccd1 vccd1 _6897_/B sky130_fd_sc_hd__nand2_1
X_5904_ _5904_/A _5904_/B vssd1 vssd1 vccd1 vccd1 _5921_/B sky130_fd_sc_hd__and2_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5835_ _5826_/A _5826_/B _5826_/C _5866_/A vssd1 vssd1 vccd1 vccd1 _5838_/A sky130_fd_sc_hd__a31o_4
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5766_ _5767_/A _5767_/B vssd1 vssd1 vccd1 vccd1 _5766_/Y sky130_fd_sc_hd__nand2b_1
X_7505_ _7485_/X _7504_/X _7657_/B vssd1 vssd1 vccd1 vccd1 _7797_/B sky130_fd_sc_hd__mux2_2
X_4717_ _4717_/A _4717_/B vssd1 vssd1 vccd1 vccd1 _4718_/C sky130_fd_sc_hd__and2_1
X_5697_ _5697_/A _5697_/B vssd1 vssd1 vccd1 vccd1 _5700_/B sky130_fd_sc_hd__xnor2_4
X_7436_ _7436_/A _7436_/B vssd1 vssd1 vccd1 vccd1 _7524_/B sky130_fd_sc_hd__xor2_2
X_4648_ _4648_/A _4648_/B _4648_/C vssd1 vssd1 vccd1 vccd1 _4650_/B sky130_fd_sc_hd__nand3_4
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7367_ _7367_/A _7367_/B vssd1 vssd1 vccd1 vccd1 _7369_/B sky130_fd_sc_hd__nor2_1
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4579_ _4569_/X _4571_/Y _4577_/A _4578_/X vssd1 vssd1 vccd1 vccd1 _4583_/A sky130_fd_sc_hd__o211a_2
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6318_ _6007_/A _6766_/S _6317_/Y vssd1 vssd1 vccd1 vccd1 _6577_/A sky130_fd_sc_hd__a21oi_4
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7298_ _7371_/A _7294_/B _7294_/C vssd1 vssd1 vccd1 vccd1 _7299_/B sky130_fd_sc_hd__o21ai_1
XFILLER_103_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6249_ _6193_/A _6131_/X _6225_/S _6248_/X _6245_/X vssd1 vssd1 vccd1 vccd1 _6249_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5620_ _5714_/A _7195_/B _5714_/C vssd1 vssd1 vccd1 vccd1 _5666_/B sky130_fd_sc_hd__and3_2
X_5551_ _5551_/A _5551_/B vssd1 vssd1 vccd1 vccd1 _5554_/B sky130_fd_sc_hd__xnor2_1
X_4502_ _7165_/A _4585_/B vssd1 vssd1 vccd1 vccd1 _4503_/B sky130_fd_sc_hd__nand2_4
XFILLER_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5482_ _5482_/A _5482_/B vssd1 vssd1 vccd1 vccd1 _5485_/A sky130_fd_sc_hd__xnor2_2
X_7221_ _7242_/A _7242_/B vssd1 vssd1 vccd1 vccd1 _7243_/A sky130_fd_sc_hd__nor2_1
X_4433_ _4366_/X _4396_/Y _4432_/Y _4360_/Y vssd1 vssd1 vccd1 vccd1 _4433_/X sky130_fd_sc_hd__o22a_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4364_ _4334_/A _4334_/B _4376_/B _4376_/C vssd1 vssd1 vccd1 vccd1 _4407_/B sky130_fd_sc_hd__o2bb2a_4
X_7152_ _7371_/A _7150_/B _7156_/B _7149_/Y vssd1 vssd1 vccd1 vccd1 _7154_/B sky130_fd_sc_hd__o31a_1
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6103_ _6104_/A _6104_/B vssd1 vssd1 vccd1 vccd1 _6111_/B sky130_fd_sc_hd__xor2_4
X_4295_ _6278_/A _5134_/A2 _4292_/X _5135_/C1 vssd1 vssd1 vccd1 vccd1 _4296_/B sky130_fd_sc_hd__a211o_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7083_ _7027_/A _7344_/B _7027_/C vssd1 vssd1 vccd1 vccd1 _7084_/B sky130_fd_sc_hd__o21ai_2
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6034_ _6034_/A _6296_/A vssd1 vssd1 vccd1 vccd1 _6034_/Y sky130_fd_sc_hd__xnor2_4
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7985_ _8021_/Q _8061_/Q _7986_/S vssd1 vssd1 vccd1 vccd1 _8061_/D sky130_fd_sc_hd__mux2_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6936_ _6936_/A _6988_/A vssd1 vssd1 vccd1 vccd1 _6937_/B sky130_fd_sc_hd__and2_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6867_ _6884_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _6887_/A sky130_fd_sc_hd__nand2b_1
XFILLER_22_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6798_ _6798_/A _6798_/B vssd1 vssd1 vccd1 vccd1 _6799_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5818_ _5794_/A _5794_/B _5794_/C vssd1 vssd1 vccd1 vccd1 _5826_/B sky130_fd_sc_hd__a21o_1
X_5749_ _5750_/A _5750_/B _5750_/C vssd1 vssd1 vccd1 vccd1 _5749_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7419_ _7419_/A _7419_/B _7438_/A _7436_/B vssd1 vssd1 vccd1 vccd1 _7424_/A sky130_fd_sc_hd__or4b_4
XFILLER_104_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4080_ _4081_/B _4080_/B _4080_/C vssd1 vssd1 vccd1 vccd1 _4080_/X sky130_fd_sc_hd__and3b_4
XFILLER_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7770_ _7798_/A _7770_/B vssd1 vssd1 vccd1 vccd1 _7795_/B sky130_fd_sc_hd__nand2_2
XFILLER_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4982_ _5040_/A _5040_/B vssd1 vssd1 vccd1 vccd1 _4984_/B sky130_fd_sc_hd__and2_2
X_6721_ _6712_/X _6720_/X _6739_/S vssd1 vssd1 vccd1 vccd1 _6721_/X sky130_fd_sc_hd__mux2_1
X_6652_ _6713_/S _6697_/S vssd1 vssd1 vccd1 vccd1 _6652_/Y sky130_fd_sc_hd__nor2_1
X_5603_ _5597_/A _5597_/B _5598_/Y vssd1 vssd1 vccd1 vccd1 _5660_/A sky130_fd_sc_hd__a21bo_2
XFILLER_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6583_ _7886_/A _6583_/B vssd1 vssd1 vccd1 vccd1 _6584_/B sky130_fd_sc_hd__nor2_1
X_5534_ _5534_/A _5534_/B vssd1 vssd1 vccd1 vccd1 _5537_/B sky130_fd_sc_hd__xnor2_4
X_5465_ _5465_/A _6871_/B vssd1 vssd1 vccd1 vccd1 _5467_/A sky130_fd_sc_hd__nand2_2
X_7204_ _7204_/A _7204_/B vssd1 vssd1 vccd1 vccd1 _7229_/A sky130_fd_sc_hd__xnor2_4
X_4416_ _4413_/X _4414_/X _4377_/A _4455_/A vssd1 vssd1 vccd1 vccd1 _4416_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5396_ _5551_/A _5551_/B _5359_/Y vssd1 vssd1 vccd1 vccd1 _5426_/A sky130_fd_sc_hd__a21oi_4
X_7135_ _7135_/A _7135_/B vssd1 vssd1 vccd1 vccd1 _7158_/A sky130_fd_sc_hd__xnor2_4
X_4347_ _4340_/A _4340_/B _4551_/A _4406_/A vssd1 vssd1 vccd1 vccd1 _4430_/C sky130_fd_sc_hd__a22o_4
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4278_ _4219_/Y _4276_/X _4277_/X vssd1 vssd1 vccd1 vccd1 _4278_/Y sky130_fd_sc_hd__a21oi_2
X_7066_ _7067_/A _7067_/B vssd1 vssd1 vccd1 vccd1 _7066_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6017_ _6017_/A _6017_/B vssd1 vssd1 vccd1 vccd1 _6024_/A sky130_fd_sc_hd__xnor2_2
XFILLER_67_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7968_ _8048_/Q _7970_/C _7967_/Y vssd1 vssd1 vccd1 vccd1 _8048_/D sky130_fd_sc_hd__a21oi_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7899_ _7649_/A _7869_/A _7869_/B vssd1 vssd1 vccd1 vccd1 _7900_/B sky130_fd_sc_hd__o21ai_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6919_ _6919_/A _6919_/B vssd1 vssd1 vccd1 vccd1 _6968_/B sky130_fd_sc_hd__nor2_4
XFILLER_52_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5250_ _5259_/A _5399_/A vssd1 vssd1 vccd1 vccd1 _5250_/Y sky130_fd_sc_hd__nor2_1
X_4201_ _4216_/B _4200_/B _4199_/X vssd1 vssd1 vccd1 vccd1 _4201_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5181_ _5181_/A _5181_/B vssd1 vssd1 vccd1 vccd1 _5220_/A sky130_fd_sc_hd__nand2_4
X_4132_ _4074_/Y _4118_/X _4056_/S _4071_/Y vssd1 vssd1 vccd1 vccd1 _4132_/X sky130_fd_sc_hd__o211a_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4063_ _4063_/A _4117_/C vssd1 vssd1 vccd1 vccd1 _4064_/B sky130_fd_sc_hd__nor2_4
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7822_ _7822_/A _7822_/B vssd1 vssd1 vccd1 vccd1 _7823_/B sky130_fd_sc_hd__or2_1
XFILLER_91_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7753_ _7562_/B _7751_/X _7752_/X vssd1 vssd1 vccd1 vccd1 _7754_/B sky130_fd_sc_hd__o21ba_1
X_4965_ _4965_/A _4965_/B vssd1 vssd1 vccd1 vccd1 _5003_/A sky130_fd_sc_hd__xnor2_4
X_6704_ _6751_/S _6704_/B vssd1 vssd1 vccd1 vccd1 _6704_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7684_ _7684_/A _7684_/B vssd1 vssd1 vccd1 vccd1 _7707_/A sky130_fd_sc_hd__nor2_1
X_4896_ _4929_/A _5041_/D1 _4844_/X _4732_/X vssd1 vssd1 vccd1 vccd1 _4897_/B sky130_fd_sc_hd__o211ai_1
XFILLER_20_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6635_ _6635_/A _6635_/B vssd1 vssd1 vccd1 vccd1 _6635_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_22_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6566_ _6578_/A _6567_/B vssd1 vssd1 vccd1 vccd1 _6617_/B sky130_fd_sc_hd__and2b_1
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5517_ _7281_/C _5723_/A vssd1 vssd1 vccd1 vccd1 _5575_/A sky130_fd_sc_hd__nand2_2
XFILLER_118_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6497_ _6443_/A _6394_/B _6496_/X vssd1 vssd1 vccd1 vccd1 _6570_/A sky130_fd_sc_hd__o21ai_4
X_5448_ _5449_/A _5449_/B vssd1 vssd1 vccd1 vccd1 _5448_/Y sky130_fd_sc_hd__nand2b_1
Xfanout100 _6448_/S vssd1 vssd1 vccd1 vccd1 _6445_/S sky130_fd_sc_hd__buf_6
Xfanout122 _4356_/Y vssd1 vssd1 vccd1 vccd1 _7284_/A sky130_fd_sc_hd__clkbuf_16
X_5379_ _5379_/A _5379_/B vssd1 vssd1 vccd1 vccd1 _5689_/B sky130_fd_sc_hd__or2_4
Xfanout111 _7281_/D vssd1 vssd1 vccd1 vccd1 _5919_/A sky130_fd_sc_hd__buf_6
XFILLER_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout144 _6999_/A vssd1 vssd1 vccd1 vccd1 _7165_/A sky130_fd_sc_hd__buf_6
Xfanout155 _6878_/C vssd1 vssd1 vccd1 vccd1 _4501_/A sky130_fd_sc_hd__clkbuf_8
Xfanout133 _7247_/A vssd1 vssd1 vccd1 vccd1 _7334_/A sky130_fd_sc_hd__buf_6
X_7118_ _7119_/A _7119_/B vssd1 vssd1 vccd1 vccd1 _7134_/B sky130_fd_sc_hd__or2_2
XFILLER_101_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout199 _6800_/B vssd1 vssd1 vccd1 vccd1 _6805_/B sky130_fd_sc_hd__buf_12
XFILLER_86_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout166 _5087_/B vssd1 vssd1 vccd1 vccd1 _5977_/B sky130_fd_sc_hd__buf_12
Xfanout188 _5990_/B vssd1 vssd1 vccd1 vccd1 _5989_/B sky130_fd_sc_hd__buf_8
XFILLER_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7049_ _7049_/A _7049_/B vssd1 vssd1 vccd1 vccd1 _7440_/A sky130_fd_sc_hd__nor2_1
Xfanout177 _4342_/X vssd1 vssd1 vccd1 vccd1 _6902_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _5019_/A _4751_/C _5090_/B _5020_/A vssd1 vssd1 vccd1 vccd1 _4750_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4681_ _4687_/A _4681_/B vssd1 vssd1 vccd1 vccd1 _4714_/B sky130_fd_sc_hd__nor2_1
X_6420_ _7319_/B _6951_/A _6456_/S vssd1 vssd1 vccd1 vccd1 _6420_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6351_ _7402_/A vssd1 vssd1 vccd1 vccd1 _6368_/A sky130_fd_sc_hd__inv_2
XFILLER_108_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5302_ _6800_/B _5755_/A vssd1 vssd1 vccd1 vccd1 _5432_/A sky130_fd_sc_hd__nor2_8
X_6282_ _6274_/A _6274_/B _6281_/X vssd1 vssd1 vccd1 vccd1 _6282_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_5_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8021_ _8077_/CLK _8021_/D vssd1 vssd1 vccd1 vccd1 _8021_/Q sky130_fd_sc_hd__dfxtp_1
X_5233_ _5959_/B _5233_/B vssd1 vssd1 vccd1 vccd1 _5236_/A sky130_fd_sc_hd__nand2_1
X_5164_ _6806_/A _5207_/A vssd1 vssd1 vccd1 vccd1 _5164_/X sky130_fd_sc_hd__or2_1
XFILLER_96_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4115_ _4102_/A _4114_/Y _4095_/B vssd1 vssd1 vccd1 vccd1 _4115_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_69_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5095_ _5095_/A _5095_/B _5095_/C vssd1 vssd1 vccd1 vccd1 _5098_/A sky130_fd_sc_hd__and3_1
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4046_ _8065_/Q _4046_/B vssd1 vssd1 vccd1 vccd1 _4046_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_83_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7805_ _8036_/Q _7944_/B _7803_/X _7804_/X vssd1 vssd1 vccd1 vccd1 _7806_/B sky130_fd_sc_hd__a22oi_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5997_ _6017_/B _6027_/A vssd1 vssd1 vccd1 vccd1 _5997_/Y sky130_fd_sc_hd__nand2_1
X_7736_ _7894_/A _6732_/C _6634_/Y vssd1 vssd1 vccd1 vccd1 _7738_/B sky130_fd_sc_hd__o21a_1
X_4948_ _5014_/A _5013_/C vssd1 vssd1 vccd1 vccd1 _4986_/A sky130_fd_sc_hd__nor2_4
X_7667_ _7639_/B _6170_/X _7639_/Y vssd1 vssd1 vccd1 vccd1 _7667_/Y sky130_fd_sc_hd__o21ai_2
X_4879_ _4879_/A _4879_/B vssd1 vssd1 vccd1 vccd1 _4880_/B sky130_fd_sc_hd__nand2_1
X_6618_ _6626_/C _6618_/B vssd1 vssd1 vccd1 vccd1 _6621_/B sky130_fd_sc_hd__or2_2
X_7598_ _7939_/A _7623_/A _7623_/B vssd1 vssd1 vccd1 vccd1 _7600_/B sky130_fd_sc_hd__and3_1
XFILLER_106_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6549_ _6549_/A _6549_/B vssd1 vssd1 vccd1 vccd1 _6581_/A sky130_fd_sc_hd__xnor2_4
XFILLER_4_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5920_ _5919_/A _5927_/B _5919_/C vssd1 vssd1 vccd1 vccd1 _6236_/B sky130_fd_sc_hd__a21oi_1
XFILLER_80_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5851_ _5851_/A _5851_/B vssd1 vssd1 vccd1 vccd1 _5871_/A sky130_fd_sc_hd__xor2_4
X_4802_ _4851_/A _4818_/B vssd1 vssd1 vccd1 vccd1 _4805_/C sky130_fd_sc_hd__nand2_1
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5782_ _5782_/A _5927_/B _5813_/B vssd1 vssd1 vccd1 vccd1 _5782_/X sky130_fd_sc_hd__and3_1
X_7521_ _7370_/B _7519_/X _7520_/Y vssd1 vssd1 vccd1 vccd1 _7521_/Y sky130_fd_sc_hd__o21ai_1
X_4733_ _4692_/Y _4836_/A _4708_/X _4710_/Y vssd1 vssd1 vccd1 vccd1 _4846_/B sky130_fd_sc_hd__o31ai_4
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7452_ _7452_/A _7452_/B vssd1 vssd1 vccd1 vccd1 _7452_/X sky130_fd_sc_hd__xor2_1
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6403_ _6488_/A _6362_/Y _6402_/X _6441_/S vssd1 vssd1 vccd1 vccd1 _6404_/B sky130_fd_sc_hd__a2bb2o_2
X_4664_ _4664_/A _4664_/B vssd1 vssd1 vccd1 vccd1 _4665_/C sky130_fd_sc_hd__xnor2_2
X_7383_ _7439_/A _7439_/B _7106_/A vssd1 vssd1 vccd1 vccd1 _7440_/B sky130_fd_sc_hd__o21ai_2
X_4595_ _4594_/B _4594_/C _4594_/A vssd1 vssd1 vccd1 vccd1 _4596_/C sky130_fd_sc_hd__a21o_1
X_6334_ _6338_/A _6336_/B vssd1 vssd1 vccd1 vccd1 _6334_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_115_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6265_ _6211_/X _6212_/X _7784_/A vssd1 vssd1 vccd1 vccd1 _6265_/X sky130_fd_sc_hd__a21o_1
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8004_ _8079_/Q _8023_/Q _8004_/S vssd1 vssd1 vccd1 vccd1 _8079_/D sky130_fd_sc_hd__mux2_1
X_5216_ _5240_/A _5240_/B vssd1 vssd1 vccd1 vccd1 _5216_/Y sky130_fd_sc_hd__nand2_1
X_6196_ _6194_/X _6195_/X _7570_/B vssd1 vssd1 vccd1 vccd1 _6196_/X sky130_fd_sc_hd__mux2_2
XFILLER_111_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5147_ _5087_/B _4296_/Y _5145_/X _5322_/A vssd1 vssd1 vccd1 vccd1 _5147_/X sky130_fd_sc_hd__a211o_1
XFILLER_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5078_ _5582_/A _5367_/A vssd1 vssd1 vccd1 vccd1 _5103_/B sky130_fd_sc_hd__nor2_4
X_4029_ _8018_/Q _8019_/Q _7955_/S vssd1 vssd1 vccd1 vccd1 _8019_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7719_ _7720_/A _7720_/B vssd1 vssd1 vccd1 vccd1 _7738_/A sky130_fd_sc_hd__and2b_1
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4380_ _4359_/Y _4424_/A _4378_/X _4379_/Y _7085_/A vssd1 vssd1 vccd1 vccd1 _4380_/X
+ sky130_fd_sc_hd__a2111o_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _6326_/A _6274_/A _4080_/X vssd1 vssd1 vccd1 vccd1 _6050_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_86_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5001_ _5001_/A _5001_/B vssd1 vssd1 vccd1 vccd1 _5010_/B sky130_fd_sc_hd__xor2_4
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6952_ _7123_/A _7269_/B vssd1 vssd1 vccd1 vccd1 _7006_/A sky130_fd_sc_hd__nand2_2
X_6883_ _7123_/A _7114_/B _6903_/B vssd1 vssd1 vccd1 vccd1 _6884_/B sky130_fd_sc_hd__a21o_1
XFILLER_34_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5903_ _5884_/B _5884_/C _5927_/C vssd1 vssd1 vccd1 vccd1 _5904_/B sky130_fd_sc_hd__o21ai_1
XFILLER_62_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5834_ _5834_/A _5834_/B _5834_/C vssd1 vssd1 vccd1 vccd1 _5866_/A sky130_fd_sc_hd__and3_2
XFILLER_14_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5765_ _5765_/A _5765_/B vssd1 vssd1 vccd1 vccd1 _5767_/B sky130_fd_sc_hd__xor2_4
X_7504_ _7503_/Y _7467_/X _7624_/S vssd1 vssd1 vccd1 vccd1 _7504_/X sky130_fd_sc_hd__mux2_1
X_4716_ _4716_/A _4716_/B vssd1 vssd1 vccd1 vccd1 _4717_/B sky130_fd_sc_hd__or2_1
X_5696_ _5740_/A _5740_/B _5687_/Y vssd1 vssd1 vccd1 vccd1 _5700_/A sky130_fd_sc_hd__a21bo_4
X_7435_ _7438_/A _7436_/B _7430_/A _7889_/A _7657_/B vssd1 vssd1 vccd1 vccd1 _7554_/A
+ sky130_fd_sc_hd__a32o_1
X_4647_ _4646_/C _4646_/B _4636_/B vssd1 vssd1 vccd1 vccd1 _4648_/C sky130_fd_sc_hd__a21bo_2
X_7366_ _7366_/A _7366_/B _7366_/C _7365_/X vssd1 vssd1 vccd1 vccd1 _7367_/B sky130_fd_sc_hd__or4b_1
XFILLER_89_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6317_ _6317_/A _6766_/S vssd1 vssd1 vccd1 vccd1 _6317_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4578_ _4498_/B _4575_/Y _4573_/Y _4574_/A vssd1 vssd1 vccd1 vccd1 _4578_/X sky130_fd_sc_hd__a211o_2
XFILLER_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7297_ _7297_/A _7297_/B vssd1 vssd1 vccd1 vccd1 _7488_/A sky130_fd_sc_hd__xnor2_4
XFILLER_89_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6248_ _6248_/A _6248_/B vssd1 vssd1 vccd1 vccd1 _6248_/X sky130_fd_sc_hd__or2_1
X_6179_ _6178_/X _6176_/X _6199_/S vssd1 vssd1 vccd1 vccd1 _6179_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5550_ _5560_/A _5560_/B _5540_/Y vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__a21o_1
XFILLER_31_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5481_ _5468_/A _5467_/A _5467_/B _5469_/X vssd1 vssd1 vccd1 vccd1 _5487_/A sky130_fd_sc_hd__a31o_4
X_4501_ _4501_/A _4551_/B vssd1 vssd1 vccd1 vccd1 _4505_/A sky130_fd_sc_hd__nand2_4
X_7220_ _7220_/A _7220_/B vssd1 vssd1 vccd1 vccd1 _7242_/B sky130_fd_sc_hd__xnor2_1
X_4432_ _7245_/A _4407_/A _7215_/A vssd1 vssd1 vccd1 vccd1 _4432_/Y sky130_fd_sc_hd__a21oi_1
X_7151_ _7151_/A _7151_/B vssd1 vssd1 vccd1 vccd1 _7156_/B sky130_fd_sc_hd__xor2_4
X_4363_ _4430_/B _4430_/C _7136_/A _4430_/A vssd1 vssd1 vccd1 vccd1 _4363_/X sky130_fd_sc_hd__a211o_1
XFILLER_112_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6102_ _6102_/A _6102_/B vssd1 vssd1 vccd1 vccd1 _6104_/B sky130_fd_sc_hd__xnor2_4
X_4294_ _4094_/B _5134_/A2 _4293_/X _4303_/B vssd1 vssd1 vccd1 vccd1 _4296_/A sky130_fd_sc_hd__a211o_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7082_ _7082_/A _7082_/B vssd1 vssd1 vccd1 vccd1 _7090_/A sky130_fd_sc_hd__or2_4
XFILLER_112_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6033_ _6326_/B _6033_/B vssd1 vssd1 vccd1 vccd1 _6296_/A sky130_fd_sc_hd__or2_4
XFILLER_58_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7984_ _8020_/Q _8060_/Q _7986_/S vssd1 vssd1 vccd1 vccd1 _8060_/D sky130_fd_sc_hd__mux2_1
XFILLER_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6935_ _6936_/A _6988_/A vssd1 vssd1 vccd1 vccd1 _6937_/A sky130_fd_sc_hd__nor2_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6866_ _6866_/A _6866_/B vssd1 vssd1 vccd1 vccd1 _6868_/B sky130_fd_sc_hd__xnor2_4
X_6797_ _6798_/A _6798_/B vssd1 vssd1 vccd1 vccd1 _6804_/A sky130_fd_sc_hd__or2_1
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5817_ _5817_/A _5817_/B vssd1 vssd1 vccd1 vccd1 _5848_/A sky130_fd_sc_hd__xor2_2
X_5748_ _5748_/A _5748_/B vssd1 vssd1 vccd1 vccd1 _5750_/C sky130_fd_sc_hd__xor2_2
X_5679_ _5679_/A _5679_/B vssd1 vssd1 vccd1 vccd1 _5681_/B sky130_fd_sc_hd__xnor2_4
X_7418_ _7421_/C _7418_/B vssd1 vssd1 vccd1 vccd1 _7419_/B sky130_fd_sc_hd__xnor2_1
XFILLER_116_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7349_ _7349_/A _7349_/B vssd1 vssd1 vccd1 vccd1 _7374_/A sky130_fd_sc_hd__xnor2_2
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4981_ _5013_/A _5013_/C _5013_/B _4947_/C vssd1 vssd1 vccd1 vccd1 _4984_/A sky130_fd_sc_hd__or4b_2
X_6720_ _6689_/S _6694_/X _6719_/Y _6645_/A vssd1 vssd1 vccd1 vccd1 _6720_/X sky130_fd_sc_hd__a211o_4
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6651_ _6651_/A vssd1 vssd1 vccd1 vccd1 _6651_/Y sky130_fd_sc_hd__inv_2
X_6582_ _6546_/A _6581_/Y _6547_/A vssd1 vssd1 vccd1 vccd1 _6582_/X sky130_fd_sc_hd__o21a_1
X_5602_ _5604_/A _5604_/B vssd1 vssd1 vccd1 vccd1 _5616_/A sky130_fd_sc_hd__or2_2
XFILLER_32_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5533_ _5518_/A _5574_/A _5520_/Y vssd1 vssd1 vccd1 vccd1 _5537_/A sky130_fd_sc_hd__o21ai_4
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5464_ _5275_/C _5464_/B _6783_/A vssd1 vssd1 vccd1 vccd1 _5466_/B sky130_fd_sc_hd__and3b_1
XFILLER_117_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4415_ _4413_/X _4414_/X _4455_/A vssd1 vssd1 vccd1 vccd1 _4488_/B sky130_fd_sc_hd__a21o_1
X_5395_ _5395_/A _5395_/B vssd1 vssd1 vccd1 vccd1 _5551_/B sky130_fd_sc_hd__xnor2_4
X_7203_ _7203_/A _7203_/B vssd1 vssd1 vccd1 vccd1 _7232_/A sky130_fd_sc_hd__xnor2_4
X_4346_ _4406_/A _4551_/A vssd1 vssd1 vccd1 vccd1 _4412_/A sky130_fd_sc_hd__nand2_4
X_7134_ _7135_/A _7134_/B _7160_/A vssd1 vssd1 vccd1 vccd1 _7134_/X sky130_fd_sc_hd__and3_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4277_ _4242_/A _6017_/A _4548_/C _6035_/A0 vssd1 vssd1 vccd1 vccd1 _4277_/X sky130_fd_sc_hd__a211o_1
X_7065_ _5977_/B _5133_/Y _5136_/Y _7284_/A _5322_/A vssd1 vssd1 vccd1 vccd1 _7173_/A
+ sky130_fd_sc_hd__a2111oi_4
X_6016_ _6077_/A vssd1 vssd1 vccd1 vccd1 _6078_/B sky130_fd_sc_hd__clkinv_4
XFILLER_39_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7967_ _8048_/Q _7970_/C _7971_/B vssd1 vssd1 vccd1 vccd1 _7967_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7898_ _7921_/A _7898_/B vssd1 vssd1 vccd1 vccd1 _7900_/A sky130_fd_sc_hd__nor2_1
X_6918_ _4320_/X _7306_/B _6916_/C vssd1 vssd1 vccd1 vccd1 _6919_/B sky130_fd_sc_hd__a21oi_2
X_6849_ _6849_/A _6849_/B vssd1 vssd1 vccd1 vccd1 _6850_/B sky130_fd_sc_hd__and2_1
XFILLER_10_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4200_ _4216_/B _4200_/B vssd1 vssd1 vccd1 vccd1 _4200_/Y sky130_fd_sc_hd__nand2_1
X_5180_ _5180_/A _5180_/B vssd1 vssd1 vccd1 vccd1 _5181_/B sky130_fd_sc_hd__or2_2
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4131_ _4050_/Y _4303_/C _4130_/X _6021_/A0 vssd1 vssd1 vccd1 vccd1 _4131_/X sky130_fd_sc_hd__o211a_1
XFILLER_110_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4062_ _6272_/A _4062_/B vssd1 vssd1 vccd1 vccd1 _4117_/C sky130_fd_sc_hd__xnor2_4
XFILLER_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7821_ _7822_/A _7822_/B vssd1 vssd1 vccd1 vccd1 _7823_/A sky130_fd_sc_hd__nand2_2
XFILLER_64_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7752_ _8033_/Q _4018_/X _7857_/B _8034_/Q vssd1 vssd1 vccd1 vccd1 _7752_/X sky130_fd_sc_hd__a22o_1
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4964_ _4965_/A _4965_/B vssd1 vssd1 vccd1 vccd1 _4964_/X sky130_fd_sc_hd__and2b_1
X_6703_ _6653_/X _6672_/A _6733_/S vssd1 vssd1 vccd1 vccd1 _6703_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7683_ _7923_/A _7683_/B _7721_/B vssd1 vssd1 vccd1 vccd1 _7683_/X sky130_fd_sc_hd__and3_1
X_4895_ _4903_/A _4903_/B vssd1 vssd1 vccd1 vccd1 _4905_/A sky130_fd_sc_hd__nand2b_2
X_6634_ _6635_/A _6635_/B vssd1 vssd1 vccd1 vccd1 _6634_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6565_ _6565_/A _6565_/B vssd1 vssd1 vccd1 vccd1 _6567_/B sky130_fd_sc_hd__and2_1
X_6496_ _6347_/Y _6432_/X _6495_/X _6488_/B vssd1 vssd1 vccd1 vccd1 _6496_/X sky130_fd_sc_hd__a211o_2
X_5516_ _5516_/A _5800_/A vssd1 vssd1 vccd1 vccd1 _5574_/A sky130_fd_sc_hd__or2_2
X_5447_ _5464_/B _5275_/C _5470_/A _5446_/X vssd1 vssd1 vccd1 vccd1 _5449_/B sky130_fd_sc_hd__o211a_4
Xfanout112 _5315_/X vssd1 vssd1 vccd1 vccd1 _7281_/D sky130_fd_sc_hd__buf_8
Xfanout101 _5969_/Y vssd1 vssd1 vccd1 vccd1 _6139_/B sky130_fd_sc_hd__clkbuf_8
X_5378_ _5378_/A _5908_/A _5378_/C vssd1 vssd1 vccd1 vccd1 _5379_/B sky130_fd_sc_hd__and3_1
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout123 _4355_/Y vssd1 vssd1 vccd1 vccd1 _7285_/A sky130_fd_sc_hd__buf_8
X_4329_ _6034_/A _4327_/X _4328_/Y _4266_/X vssd1 vssd1 vccd1 vccd1 _4329_/X sky130_fd_sc_hd__o2bb2a_4
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout134 _4354_/X vssd1 vssd1 vccd1 vccd1 _7247_/A sky130_fd_sc_hd__clkbuf_16
Xfanout156 _4330_/X vssd1 vssd1 vccd1 vccd1 _6878_/C sky130_fd_sc_hd__buf_6
Xfanout145 _4339_/Y vssd1 vssd1 vccd1 vccd1 _6999_/A sky130_fd_sc_hd__buf_8
X_7117_ _7161_/A _7161_/B vssd1 vssd1 vccd1 vccd1 _7119_/B sky130_fd_sc_hd__nand2_1
Xfanout167 _6030_/A vssd1 vssd1 vccd1 vccd1 _5087_/B sky130_fd_sc_hd__buf_8
Xfanout189 _6017_/A vssd1 vssd1 vccd1 vccd1 _4315_/B sky130_fd_sc_hd__buf_4
X_7048_ _7048_/A _7048_/B _7051_/A vssd1 vssd1 vccd1 vccd1 _7049_/B sky130_fd_sc_hd__and3_1
Xfanout178 _7213_/B vssd1 vssd1 vccd1 vccd1 _4551_/A sky130_fd_sc_hd__buf_8
XFILLER_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4680_ _4679_/C _4717_/A vssd1 vssd1 vccd1 vccd1 _4681_/B sky130_fd_sc_hd__and2b_1
XFILLER_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6350_ _6350_/A _6350_/B vssd1 vssd1 vccd1 vccd1 _7402_/A sky130_fd_sc_hd__or2_4
XFILLER_115_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5301_ _7235_/B _5880_/A vssd1 vssd1 vccd1 vccd1 _5666_/A sky130_fd_sc_hd__nor2_4
X_6281_ _4094_/B _4190_/Y _6279_/X _6280_/X vssd1 vssd1 vccd1 vccd1 _6281_/X sky130_fd_sc_hd__o22a_1
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8020_ _8077_/CLK _8020_/D vssd1 vssd1 vccd1 vccd1 _8020_/Q sky130_fd_sc_hd__dfxtp_1
X_5232_ _5232_/A _5232_/B _5232_/C vssd1 vssd1 vccd1 vccd1 _5233_/B sky130_fd_sc_hd__or3_1
X_5163_ _5541_/A _5386_/A vssd1 vssd1 vccd1 vccd1 _5956_/A sky130_fd_sc_hd__or2_4
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4114_ _4084_/X _4113_/X _4102_/B vssd1 vssd1 vccd1 vccd1 _4114_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5094_ _4746_/A _5093_/Y _4752_/Y vssd1 vssd1 vccd1 vccd1 _5095_/C sky130_fd_sc_hd__a21o_1
X_4045_ _8062_/Q _8061_/Q _4057_/B _5107_/C _4066_/A vssd1 vssd1 vccd1 vccd1 _4046_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7804_ _8035_/Q _7964_/C _7562_/B vssd1 vssd1 vccd1 vccd1 _7804_/X sky130_fd_sc_hd__a21bo_1
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _5996_/A _5996_/B vssd1 vssd1 vccd1 vccd1 _6000_/A sky130_fd_sc_hd__nor2_2
XFILLER_52_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7735_ _7728_/Y _7733_/X _7734_/Y vssd1 vssd1 vccd1 vccd1 _7735_/Y sky130_fd_sc_hd__o21ai_1
X_4947_ _4947_/A _4949_/A _4947_/C vssd1 vssd1 vccd1 vccd1 _4947_/X sky130_fd_sc_hd__and3_1
XFILLER_24_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7666_ _7664_/X _7665_/Y _7928_/A vssd1 vssd1 vccd1 vccd1 _8031_/D sky130_fd_sc_hd__a21oi_1
X_4878_ _4878_/A _4878_/B vssd1 vssd1 vccd1 vccd1 _4906_/A sky130_fd_sc_hd__xnor2_4
X_6617_ _6617_/A _6617_/B _6617_/C vssd1 vssd1 vccd1 vccd1 _6618_/B sky130_fd_sc_hd__nor3_1
X_7597_ _7597_/A _7597_/B vssd1 vssd1 vccd1 vccd1 _7623_/B sky130_fd_sc_hd__xnor2_2
XFILLER_20_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6548_ _7607_/A _6548_/B vssd1 vssd1 vccd1 vccd1 _6549_/B sky130_fd_sc_hd__and2_2
XFILLER_118_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6479_ _6479_/A _6479_/B vssd1 vssd1 vccd1 vccd1 _6543_/A sky130_fd_sc_hd__or2_4
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5850_ _5850_/A _5850_/B vssd1 vssd1 vccd1 vccd1 _5875_/A sky130_fd_sc_hd__xnor2_1
X_4801_ _4800_/A _4800_/B _4793_/X vssd1 vssd1 vccd1 vccd1 _4818_/B sky130_fd_sc_hd__a21oi_2
X_5781_ _5781_/A _5781_/B vssd1 vssd1 vccd1 vccd1 _5813_/B sky130_fd_sc_hd__xor2_2
X_7520_ _4355_/Y _7085_/B _7306_/C _7333_/Y _7365_/X vssd1 vssd1 vccd1 vccd1 _7520_/Y
+ sky130_fd_sc_hd__a2111oi_1
X_4732_ _4692_/Y _4836_/A _4708_/X _4709_/Y vssd1 vssd1 vccd1 vccd1 _4732_/X sky130_fd_sc_hd__o31a_2
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7451_ _7450_/X _7444_/X _7515_/S vssd1 vssd1 vccd1 vccd1 _7451_/X sky130_fd_sc_hd__mux2_1
X_4663_ _4663_/A _4663_/B _4664_/B vssd1 vssd1 vccd1 vccd1 _4670_/A sky130_fd_sc_hd__and3_1
XFILLER_119_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6402_ _6381_/B _6401_/X _6484_/S vssd1 vssd1 vccd1 vccd1 _6402_/X sky130_fd_sc_hd__mux2_1
X_7382_ _7477_/A _7477_/B _7155_/A vssd1 vssd1 vccd1 vccd1 _7439_/B sky130_fd_sc_hd__a21oi_2
X_4594_ _4594_/A _4594_/B _4594_/C vssd1 vssd1 vccd1 vccd1 _4596_/B sky130_fd_sc_hd__nand3_2
X_6333_ _6031_/B _6034_/Y _6767_/S vssd1 vssd1 vccd1 vccd1 _6336_/B sky130_fd_sc_hd__mux2_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6264_ _6196_/X _6263_/X _7639_/B vssd1 vssd1 vccd1 vccd1 _6264_/X sky130_fd_sc_hd__mux2_2
XFILLER_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8003_ _8078_/Q _8022_/Q _8004_/S vssd1 vssd1 vccd1 vccd1 _8078_/D sky130_fd_sc_hd__mux2_1
X_5215_ _5215_/A _5215_/B vssd1 vssd1 vccd1 vccd1 _5240_/B sky130_fd_sc_hd__xor2_4
X_6195_ _6176_/X _6182_/X _6199_/S vssd1 vssd1 vccd1 vccd1 _6195_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5146_ _5087_/B _4296_/Y _5145_/X _5322_/A vssd1 vssd1 vccd1 vccd1 _6873_/B sky130_fd_sc_hd__a211oi_4
XFILLER_57_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5077_ _5745_/A _5352_/A _5352_/B vssd1 vssd1 vccd1 vccd1 _5110_/A sky130_fd_sc_hd__nand3_4
X_4028_ _8017_/Q _8018_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _8018_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5979_ _6311_/A _6177_/A vssd1 vssd1 vccd1 vccd1 _6010_/B sky130_fd_sc_hd__xnor2_4
XFILLER_12_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7718_ _6757_/A _7717_/Y _7718_/S vssd1 vssd1 vccd1 vccd1 _7720_/B sky130_fd_sc_hd__mux2_2
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7649_ _7649_/A _7649_/B vssd1 vssd1 vccd1 vccd1 _7654_/A sky130_fd_sc_hd__or2_1
XFILLER_20_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5009_/A _5000_/B vssd1 vssd1 vccd1 vccd1 _5010_/A sky130_fd_sc_hd__nor2_4
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6951_ _6951_/A _7285_/A _7114_/B _6951_/D vssd1 vssd1 vccd1 vccd1 _6957_/B sky130_fd_sc_hd__and4_2
XFILLER_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6882_ _7057_/A _7046_/B _6903_/A vssd1 vssd1 vccd1 vccd1 _6882_/Y sky130_fd_sc_hd__o21ai_1
X_5902_ _5902_/A _5902_/B vssd1 vssd1 vccd1 vccd1 _5917_/A sky130_fd_sc_hd__xor2_2
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5833_ _5851_/A _5833_/B _5833_/C vssd1 vssd1 vccd1 vccd1 _5834_/C sky130_fd_sc_hd__and3_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7503_ _7403_/A _7766_/A _7438_/B _7502_/Y vssd1 vssd1 vccd1 vccd1 _7503_/Y sky130_fd_sc_hd__o31ai_1
X_5764_ _5788_/B _5788_/A vssd1 vssd1 vccd1 vccd1 _5767_/A sky130_fd_sc_hd__nand2b_4
X_5695_ _5695_/A _5695_/B vssd1 vssd1 vccd1 vccd1 _5740_/B sky130_fd_sc_hd__xnor2_4
X_4715_ _4727_/A _4727_/B vssd1 vssd1 vccd1 vccd1 _4726_/A sky130_fd_sc_hd__nor2_1
X_7434_ _7535_/A vssd1 vssd1 vccd1 vccd1 _7538_/S sky130_fd_sc_hd__clkinv_4
X_4646_ _4636_/B _4646_/B _4646_/C vssd1 vssd1 vccd1 vccd1 _4648_/B sky130_fd_sc_hd__nand3b_4
X_7365_ _7366_/C _7365_/B vssd1 vssd1 vccd1 vccd1 _7365_/X sky130_fd_sc_hd__xor2_1
X_4577_ _4577_/A vssd1 vssd1 vccd1 vccd1 _4581_/B sky130_fd_sc_hd__inv_2
XFILLER_30_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6316_ _6348_/B _6315_/Y _7401_/A vssd1 vssd1 vccd1 vccd1 _6322_/B sky130_fd_sc_hd__mux2_8
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7296_ _7297_/A _7297_/B vssd1 vssd1 vccd1 vccd1 _7296_/X sky130_fd_sc_hd__and2b_1
XFILLER_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6247_ _6232_/Y _6206_/X _6262_/S vssd1 vssd1 vccd1 vccd1 _6248_/B sky130_fd_sc_hd__mux2_1
X_6178_ _6878_/B _6139_/B _6175_/A _6242_/S _6177_/Y vssd1 vssd1 vccd1 vccd1 _6178_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5129_ _5207_/A _5198_/B vssd1 vssd1 vccd1 vccd1 _5151_/C sky130_fd_sc_hd__or2_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5480_ _5613_/A _5480_/B vssd1 vssd1 vccd1 vccd1 _6144_/A sky130_fd_sc_hd__xor2_2
X_4500_ _4455_/A _4551_/B _4458_/X _4457_/Y vssd1 vssd1 vccd1 vccd1 _4506_/A sky130_fd_sc_hd__a31o_4
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_1 _6590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4431_ _7136_/A _4349_/Y _4430_/X _4411_/A vssd1 vssd1 vccd1 vccd1 _4431_/X sky130_fd_sc_hd__o31a_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7150_ _7371_/A _7150_/B vssd1 vssd1 vccd1 vccd1 _7156_/A sky130_fd_sc_hd__nor2_1
X_4362_ _7215_/A _4441_/A _4407_/A _7261_/A _7136_/A vssd1 vssd1 vccd1 vccd1 _4362_/X
+ sky130_fd_sc_hd__o311a_1
X_6101_ _6059_/B _6096_/B _6059_/A vssd1 vssd1 vccd1 vccd1 _6102_/B sky130_fd_sc_hd__o21ba_2
X_4293_ _4074_/Y _4118_/X _6274_/A _4071_/Y vssd1 vssd1 vccd1 vccd1 _4293_/X sky130_fd_sc_hd__o211a_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7081_ _7081_/A _7081_/B _7081_/C vssd1 vssd1 vccd1 vccd1 _7082_/B sky130_fd_sc_hd__and3_1
XFILLER_100_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6032_ _6326_/B _6033_/B vssd1 vssd1 vccd1 vccd1 _6035_/S sky130_fd_sc_hd__nand2_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7983_ _8019_/Q _8059_/Q _7986_/S vssd1 vssd1 vccd1 vccd1 _8059_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6934_ _6987_/B _6987_/C _6987_/A vssd1 vssd1 vccd1 vccd1 _6988_/A sky130_fd_sc_hd__o21ai_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6865_ _7114_/B _6903_/B vssd1 vssd1 vccd1 vccd1 _6884_/A sky130_fd_sc_hd__nand2_4
XFILLER_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6796_ _6780_/A _6791_/B _6782_/B _6782_/A vssd1 vssd1 vccd1 vccd1 _6798_/B sky130_fd_sc_hd__o22a_1
X_5816_ _5816_/A vssd1 vssd1 vccd1 vccd1 _5847_/B sky130_fd_sc_hd__inv_2
XFILLER_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5747_ _5751_/A _5751_/B vssd1 vssd1 vccd1 vccd1 _5750_/B sky130_fd_sc_hd__and2_1
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7417_ _7421_/A _7421_/B _7657_/A vssd1 vssd1 vccd1 vccd1 _7418_/B sky130_fd_sc_hd__o21a_1
X_5678_ _5726_/A _5726_/B _5671_/A vssd1 vssd1 vccd1 vccd1 _5681_/A sky130_fd_sc_hd__a21oi_4
X_4629_ _4654_/A _5014_/A vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__nor2_1
X_7348_ _7348_/A _7348_/B vssd1 vssd1 vccd1 vccd1 _7508_/A sky130_fd_sc_hd__xnor2_2
XFILLER_103_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7279_ _7213_/A _7170_/B _7285_/A _7281_/D _7213_/B vssd1 vssd1 vccd1 vccd1 _7279_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_89_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4980_ _4980_/A _4980_/B vssd1 vssd1 vccd1 vccd1 _5008_/A sky130_fd_sc_hd__xor2_4
X_6650_ _6691_/A _6650_/B vssd1 vssd1 vccd1 vccd1 _6651_/A sky130_fd_sc_hd__or2_1
X_6581_ _6581_/A _6581_/B vssd1 vssd1 vccd1 vccd1 _6581_/Y sky130_fd_sc_hd__nor2_1
X_5601_ _5618_/A _5618_/B _5591_/Y vssd1 vssd1 vccd1 vccd1 _5604_/B sky130_fd_sc_hd__a21boi_2
XFILLER_118_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5532_ _5325_/A _5639_/A _5529_/Y _5585_/B vssd1 vssd1 vccd1 vccd1 _5538_/A sky130_fd_sc_hd__a2bb2oi_4
XFILLER_11_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5463_ _5440_/A _5440_/B _5438_/X vssd1 vssd1 vccd1 vccd1 _5468_/A sky130_fd_sc_hd__a21o_4
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5394_ _5394_/A _5394_/B vssd1 vssd1 vccd1 vccd1 _5395_/B sky130_fd_sc_hd__xnor2_4
X_7202_ _7202_/A _7202_/B vssd1 vssd1 vccd1 vccd1 _7234_/A sky130_fd_sc_hd__xnor2_4
X_4414_ _4412_/A _4412_/B _4441_/A vssd1 vssd1 vccd1 vccd1 _4414_/X sky130_fd_sc_hd__a21o_1
X_4345_ _4376_/A _7311_/A vssd1 vssd1 vccd1 vccd1 _4441_/B sky130_fd_sc_hd__nor2_1
X_7133_ _7135_/A _7135_/B vssd1 vssd1 vccd1 vccd1 _7133_/X sky130_fd_sc_hd__and2b_1
XFILLER_113_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4276_ _4172_/B _4169_/Y _5989_/B vssd1 vssd1 vccd1 vccd1 _4276_/X sky130_fd_sc_hd__mux2_2
X_7064_ _7091_/B _7064_/B vssd1 vssd1 vccd1 vccd1 _7111_/A sky130_fd_sc_hd__nand2_4
X_6015_ _6060_/A _6805_/B _6015_/C vssd1 vssd1 vccd1 vccd1 _6077_/A sky130_fd_sc_hd__or3_4
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7966_ _7970_/C _7966_/B _7971_/B vssd1 vssd1 vccd1 vccd1 _8047_/D sky130_fd_sc_hd__and3b_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7897_ _7867_/A _7895_/C _7773_/X vssd1 vssd1 vccd1 vccd1 _7898_/B sky130_fd_sc_hd__o21bai_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6917_ _7027_/A _6917_/B vssd1 vssd1 vccd1 vccd1 _6968_/A sky130_fd_sc_hd__nor2_4
X_6848_ _6849_/A _6849_/B vssd1 vssd1 vccd1 vccd1 _6862_/A sky130_fd_sc_hd__nor2_2
XFILLER_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6779_ _6916_/A _6878_/B vssd1 vssd1 vccd1 vccd1 _6791_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4130_ _4078_/A _4119_/Y _4062_/B _4111_/A vssd1 vssd1 vccd1 vccd1 _4130_/X sky130_fd_sc_hd__a211o_1
XFILLER_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4061_ _8060_/Q _4061_/B vssd1 vssd1 vccd1 vccd1 _4062_/B sky130_fd_sc_hd__xor2_4
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7820_ _7894_/A _7583_/X _7773_/X vssd1 vssd1 vccd1 vccd1 _7822_/B sky130_fd_sc_hd__o21ba_1
XFILLER_76_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7751_ _7802_/B2 _7750_/X _7743_/Y _7735_/Y vssd1 vssd1 vccd1 vccd1 _7751_/X sky130_fd_sc_hd__o211a_2
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4963_ _4963_/A _4963_/B vssd1 vssd1 vccd1 vccd1 _4965_/B sky130_fd_sc_hd__nor2_4
X_6702_ _6638_/Y _6657_/X _6675_/X _7616_/S _6701_/X vssd1 vssd1 vccd1 vccd1 _6732_/A
+ sky130_fd_sc_hd__a221o_1
X_7682_ _7682_/A _7682_/B vssd1 vssd1 vccd1 vccd1 _7721_/B sky130_fd_sc_hd__or2_1
X_6633_ _7616_/S _6632_/X _6631_/X vssd1 vssd1 vccd1 vccd1 _6635_/B sky130_fd_sc_hd__a21o_1
X_4894_ _4894_/A _4894_/B vssd1 vssd1 vccd1 vccd1 _4903_/B sky130_fd_sc_hd__xnor2_2
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6564_ _6564_/A _6697_/S vssd1 vssd1 vccd1 vccd1 _6565_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6495_ _6450_/Y _6495_/B vssd1 vssd1 vccd1 vccd1 _6495_/X sky130_fd_sc_hd__and2b_1
X_5515_ _5722_/A _5722_/B _7281_/C vssd1 vssd1 vccd1 vccd1 _5518_/B sky130_fd_sc_hd__and3_2
X_5446_ _6871_/B _5446_/B _6916_/C vssd1 vssd1 vccd1 vccd1 _5446_/X sky130_fd_sc_hd__or3_1
Xfanout102 _7366_/B vssd1 vssd1 vccd1 vccd1 _7371_/B sky130_fd_sc_hd__buf_8
X_5377_ _5377_/A _5377_/B vssd1 vssd1 vccd1 vccd1 _5545_/A sky130_fd_sc_hd__xor2_4
Xfanout113 _4558_/B vssd1 vssd1 vccd1 vccd1 _4988_/A sky130_fd_sc_hd__buf_8
X_4328_ _4548_/A _4356_/A vssd1 vssd1 vccd1 vccd1 _4328_/Y sky130_fd_sc_hd__nand2_1
Xfanout135 _7306_/A vssd1 vssd1 vccd1 vccd1 _7281_/A sky130_fd_sc_hd__buf_6
Xfanout146 _4642_/A vssd1 vssd1 vccd1 vccd1 _4436_/A sky130_fd_sc_hd__buf_6
X_7116_ _7116_/A _7247_/D vssd1 vssd1 vccd1 vccd1 _7161_/B sky130_fd_sc_hd__nor2_4
Xfanout124 _4411_/A vssd1 vssd1 vccd1 vccd1 _4494_/A sky130_fd_sc_hd__buf_6
XFILLER_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4259_ _6017_/A _4259_/B vssd1 vssd1 vccd1 vccd1 _6033_/B sky130_fd_sc_hd__nand2_1
Xfanout168 _4081_/X vssd1 vssd1 vccd1 vccd1 _7213_/A sky130_fd_sc_hd__buf_12
X_7047_ _7048_/B _7051_/A _7048_/A vssd1 vssd1 vccd1 vccd1 _7049_/A sky130_fd_sc_hd__a21oi_2
Xfanout157 _4602_/A vssd1 vssd1 vccd1 vccd1 _4377_/A sky130_fd_sc_hd__clkbuf_8
Xfanout179 _6951_/A vssd1 vssd1 vccd1 vccd1 _7213_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7949_ _7949_/A _7949_/B vssd1 vssd1 vccd1 vccd1 _7949_/Y sky130_fd_sc_hd__nand2_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5300_ _5029_/X _5299_/X _5703_/B vssd1 vssd1 vccd1 vccd1 _5881_/A sky130_fd_sc_hd__a21bo_2
XFILLER_115_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6280_ _4094_/B _4190_/Y _4200_/B _4098_/B vssd1 vssd1 vccd1 vccd1 _6280_/X sky130_fd_sc_hd__a22o_1
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5231_ _5232_/A _5232_/B _5232_/C vssd1 vssd1 vccd1 vccd1 _5959_/B sky130_fd_sc_hd__o21ai_2
XFILLER_69_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5162_ _5180_/A _5180_/B vssd1 vssd1 vccd1 vccd1 _5181_/A sky130_fd_sc_hd__nand2_2
X_4113_ _4112_/Y _4087_/B _6326_/A vssd1 vssd1 vccd1 vccd1 _4113_/X sky130_fd_sc_hd__mux2_1
X_5093_ _5093_/A _5093_/B vssd1 vssd1 vccd1 vccd1 _5093_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_110_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4044_ _8064_/Q _8063_/Q vssd1 vssd1 vccd1 vccd1 _5107_/C sky130_fd_sc_hd__or2_2
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7803_ _6268_/X _7787_/X _7802_/Y _7903_/B1 vssd1 vssd1 vccd1 vccd1 _7803_/X sky130_fd_sc_hd__a211o_4
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7734_ _7728_/Y _7733_/X _6269_/X vssd1 vssd1 vccd1 vccd1 _7734_/Y sky130_fd_sc_hd__a21oi_1
X_5995_ _5995_/A _6021_/S vssd1 vssd1 vccd1 vccd1 _5996_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4946_ _4847_/X _4848_/Y _4773_/A _5013_/A vssd1 vssd1 vccd1 vccd1 _4949_/B sky130_fd_sc_hd__a211o_4
X_7665_ _8030_/Q _4018_/X _7857_/B _8031_/Q vssd1 vssd1 vccd1 vccd1 _7665_/Y sky130_fd_sc_hd__a22oi_1
X_4877_ _4878_/A _4878_/B vssd1 vssd1 vccd1 vccd1 _4877_/X sky130_fd_sc_hd__and2b_1
XFILLER_20_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6616_ _6621_/A _6616_/B _6616_/C _6616_/D vssd1 vssd1 vccd1 vccd1 _6616_/X sky130_fd_sc_hd__or4_1
X_7596_ _7597_/A _7597_/B vssd1 vssd1 vccd1 vccd1 _7629_/A sky130_fd_sc_hd__nand2b_2
X_6547_ _6547_/A _6547_/B vssd1 vssd1 vccd1 vccd1 _6555_/A sky130_fd_sc_hd__nand2_4
XFILLER_20_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6478_ _6437_/A _6478_/B vssd1 vssd1 vccd1 vccd1 _6478_/X sky130_fd_sc_hd__and2b_1
XFILLER_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5429_ _5423_/A _5423_/B _5413_/Y vssd1 vssd1 vccd1 vccd1 _5453_/A sky130_fd_sc_hd__a21o_1
XFILLER_101_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8079_ _8079_/CLK _8079_/D vssd1 vssd1 vccd1 vccd1 _8079_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4800_ _4800_/A _4800_/B vssd1 vssd1 vccd1 vccd1 _4805_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5780_ _5782_/A _5927_/B vssd1 vssd1 vccd1 vccd1 _5813_/A sky130_fd_sc_hd__nand2_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _4691_/A _4730_/A _4730_/B _4690_/A _4691_/X vssd1 vssd1 vccd1 vccd1 _4836_/B
+ sky130_fd_sc_hd__a311o_4
XFILLER_14_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7450_ _7446_/X _7449_/X _7502_/B vssd1 vssd1 vccd1 vccd1 _7450_/X sky130_fd_sc_hd__mux2_1
X_4662_ _4662_/A _5013_/B vssd1 vssd1 vccd1 vccd1 _4664_/B sky130_fd_sc_hd__nor2_2
X_6401_ _6388_/X _6400_/X _6431_/S vssd1 vssd1 vccd1 vccd1 _6401_/X sky130_fd_sc_hd__mux2_1
X_4593_ _4662_/A _5014_/A _4616_/C vssd1 vssd1 vccd1 vccd1 _4594_/C sky130_fd_sc_hd__or3_2
X_7381_ _7474_/A _7474_/B _7199_/A vssd1 vssd1 vccd1 vccd1 _7477_/B sky130_fd_sc_hd__o21ai_4
X_6332_ _6327_/B _6329_/Y _6336_/A vssd1 vssd1 vccd1 vccd1 _6338_/A sky130_fd_sc_hd__o21ba_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6263_ _6214_/X _6262_/X _7570_/B vssd1 vssd1 vccd1 vccd1 _6263_/X sky130_fd_sc_hd__mux2_1
X_8002_ _8077_/Q _8021_/Q _8007_/S vssd1 vssd1 vccd1 vccd1 _8077_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5214_ _5265_/A _5214_/B vssd1 vssd1 vccd1 vccd1 _5240_/A sky130_fd_sc_hd__xnor2_4
X_6194_ _6161_/Y _6178_/X _6199_/S vssd1 vssd1 vccd1 vccd1 _6194_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5145_ _5268_/A _5145_/B _5145_/C vssd1 vssd1 vccd1 vccd1 _5145_/X sky130_fd_sc_hd__and3_2
X_5076_ _5782_/A _5352_/A _5352_/B vssd1 vssd1 vccd1 vccd1 _5200_/A sky130_fd_sc_hd__and3_4
X_4027_ _8016_/Q _8017_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _8017_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5978_ _5973_/Y _5976_/Y _5977_/Y vssd1 vssd1 vccd1 vccd1 _6349_/B sky130_fd_sc_hd__o21ai_4
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7717_ _7717_/A vssd1 vssd1 vccd1 vccd1 _7717_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4929_ _4929_/A _5020_/B vssd1 vssd1 vccd1 vccd1 _4930_/B sky130_fd_sc_hd__and2_1
X_7648_ _7648_/A _7648_/B _7648_/C vssd1 vssd1 vccd1 vccd1 _7649_/B sky130_fd_sc_hd__and3_1
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7579_ _7579_/A _7579_/B vssd1 vssd1 vccd1 vccd1 _7648_/A sky130_fd_sc_hd__and2_2
XFILLER_109_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6950_ _7285_/A _7114_/B vssd1 vssd1 vccd1 vccd1 _7067_/B sky130_fd_sc_hd__nand2_2
XFILLER_93_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5901_ _5901_/A _5901_/B vssd1 vssd1 vccd1 vccd1 _5909_/A sky130_fd_sc_hd__or2_1
XFILLER_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6881_ _6881_/A _6881_/B vssd1 vssd1 vccd1 vccd1 _6896_/A sky130_fd_sc_hd__xnor2_2
X_5832_ _6971_/B _7285_/B _5855_/B _5855_/C vssd1 vssd1 vccd1 vccd1 _5833_/C sky130_fd_sc_hd__or4_1
X_5763_ _5763_/A _5763_/B vssd1 vssd1 vccd1 vccd1 _5788_/B sky130_fd_sc_hd__xnor2_4
X_7502_ _7766_/A _7502_/B vssd1 vssd1 vccd1 vccd1 _7502_/Y sky130_fd_sc_hd__nand2_1
X_4714_ _4714_/A _4714_/B vssd1 vssd1 vccd1 vccd1 _4727_/B sky130_fd_sc_hd__nor2_1
X_5694_ _5694_/A _5694_/B vssd1 vssd1 vccd1 vccd1 _5695_/B sky130_fd_sc_hd__xnor2_4
XFILLER_107_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7433_ _7424_/A _7431_/X _7438_/B vssd1 vssd1 vccd1 vccd1 _7433_/X sky130_fd_sc_hd__a21o_1
X_4645_ _4596_/B _4596_/C _4596_/A vssd1 vssd1 vccd1 vccd1 _4646_/B sky130_fd_sc_hd__a21o_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7364_ _7364_/A _7364_/B vssd1 vssd1 vccd1 vccd1 _7516_/A sky130_fd_sc_hd__or2_1
X_4576_ _4574_/A _4573_/Y _4575_/Y _4498_/B vssd1 vssd1 vccd1 vccd1 _4577_/A sky130_fd_sc_hd__o211ai_4
X_6315_ _6315_/A _6766_/S vssd1 vssd1 vccd1 vccd1 _6315_/Y sky130_fd_sc_hd__xnor2_2
X_7295_ _7293_/A _7293_/B _7299_/A vssd1 vssd1 vccd1 vccd1 _7297_/B sky130_fd_sc_hd__a21bo_2
X_6246_ _6156_/A _6205_/X _6231_/A _6242_/S vssd1 vssd1 vccd1 vccd1 _6248_/A sky130_fd_sc_hd__a22o_1
XFILLER_39_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6177_ _6177_/A _6177_/B vssd1 vssd1 vccd1 vccd1 _6177_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5128_ _5207_/A _5198_/B vssd1 vssd1 vccd1 vccd1 _5128_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5059_ _5247_/B _5247_/C _5058_/X _4831_/X vssd1 vssd1 vccd1 vccd1 _5062_/A sky130_fd_sc_hd__a211o_2
XFILLER_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_2 _4326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4430_ _4430_/A _4430_/B _4430_/C vssd1 vssd1 vccd1 vccd1 _4430_/X sky130_fd_sc_hd__and3_1
XFILLER_98_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6100_ _6088_/Y _6092_/B _6095_/X _7639_/A vssd1 vssd1 vccd1 vccd1 _6104_/A sky130_fd_sc_hd__o31a_4
X_4361_ _4430_/B _6999_/A _4412_/B _7085_/A vssd1 vssd1 vccd1 vccd1 _4361_/X sky130_fd_sc_hd__a31o_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4292_ _4074_/Y _4118_/X _4098_/B _4071_/Y vssd1 vssd1 vccd1 vccd1 _4292_/X sky130_fd_sc_hd__o211a_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7080_ _7081_/A _7081_/B _7081_/C vssd1 vssd1 vccd1 vccd1 _7082_/A sky130_fd_sc_hd__a21oi_1
X_6031_ _6031_/A _6031_/B vssd1 vssd1 vccd1 vccd1 _6038_/B sky130_fd_sc_hd__xnor2_2
XFILLER_79_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7982_ _8018_/Q _8058_/Q _7986_/S vssd1 vssd1 vccd1 vccd1 _8058_/D sky130_fd_sc_hd__mux2_1
XFILLER_81_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6933_ _6939_/B _6939_/A vssd1 vssd1 vccd1 vccd1 _6987_/C sky130_fd_sc_hd__and2b_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6864_ _7123_/A _6951_/A _7195_/B _6951_/D vssd1 vssd1 vccd1 vccd1 _6903_/B sky130_fd_sc_hd__and4_4
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5815_ _5815_/A _5815_/B _5815_/C vssd1 vssd1 vccd1 vccd1 _5816_/A sky130_fd_sc_hd__and3_1
X_6795_ _6795_/A _6795_/B vssd1 vssd1 vccd1 vccd1 _6798_/A sky130_fd_sc_hd__xnor2_1
XFILLER_22_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5746_ _5746_/A _5746_/B vssd1 vssd1 vccd1 vccd1 _5751_/B sky130_fd_sc_hd__xnor2_4
XFILLER_108_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5677_ _5677_/A _5677_/B vssd1 vssd1 vccd1 vccd1 _5726_/B sky130_fd_sc_hd__xnor2_4
X_7416_ _7416_/A _7416_/B vssd1 vssd1 vccd1 vccd1 _7421_/C sky130_fd_sc_hd__xnor2_4
X_4628_ _4662_/A _5033_/A vssd1 vssd1 vccd1 vccd1 _4632_/A sky130_fd_sc_hd__nor2_2
XFILLER_116_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7347_ _7348_/B _7348_/A vssd1 vssd1 vccd1 vccd1 _7347_/X sky130_fd_sc_hd__and2b_1
X_4559_ _7116_/A _4630_/B _4630_/C vssd1 vssd1 vccd1 vccd1 _4561_/B sky130_fd_sc_hd__or3_2
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7278_ _7278_/A _7278_/B vssd1 vssd1 vccd1 vccd1 _7302_/A sky130_fd_sc_hd__xnor2_4
XFILLER_103_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6229_ _5847_/Y _6228_/X _6174_/A vssd1 vssd1 vccd1 vccd1 _6229_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6580_ _6580_/A _6580_/B vssd1 vssd1 vccd1 vccd1 _6592_/A sky130_fd_sc_hd__xor2_4
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5600_ _5600_/A _5600_/B vssd1 vssd1 vccd1 vccd1 _5618_/B sky130_fd_sc_hd__xnor2_4
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5531_ _5531_/A _5531_/B vssd1 vssd1 vccd1 vccd1 _5585_/B sky130_fd_sc_hd__xnor2_4
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5462_ _5462_/A _5462_/B vssd1 vssd1 vccd1 vccd1 _5471_/A sky130_fd_sc_hd__xnor2_4
X_7201_ _7201_/A _7201_/B vssd1 vssd1 vccd1 vccd1 _7238_/A sky130_fd_sc_hd__nor2_4
X_5393_ _5394_/A _5394_/B vssd1 vssd1 vccd1 vccd1 _5393_/Y sky130_fd_sc_hd__nand2_1
X_4413_ _4441_/B _4413_/B vssd1 vssd1 vccd1 vccd1 _4413_/X sky130_fd_sc_hd__or2_2
X_4344_ _4356_/A _4406_/A vssd1 vssd1 vccd1 vccd1 _7294_/A sky130_fd_sc_hd__nand2_8
X_7132_ _7134_/B _7160_/A vssd1 vssd1 vccd1 vccd1 _7135_/B sky130_fd_sc_hd__nand2_2
XFILLER_113_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7063_ _7063_/A _7063_/B vssd1 vssd1 vccd1 vccd1 _7064_/B sky130_fd_sc_hd__or2_2
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6014_ _6272_/B _7949_/B vssd1 vssd1 vccd1 vccd1 _6015_/C sky130_fd_sc_hd__nor2_2
X_4275_ _4356_/A _4275_/B _4275_/C vssd1 vssd1 vccd1 vccd1 _4275_/X sky130_fd_sc_hd__and3_1
XFILLER_86_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7965_ _8046_/Q _7964_/C _8047_/Q vssd1 vssd1 vccd1 vccd1 _7966_/B sky130_fd_sc_hd__a21o_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7896_ _7921_/A vssd1 vssd1 vccd1 vccd1 _7920_/A sky130_fd_sc_hd__inv_2
X_6916_ _6916_/A _7306_/B _6916_/C vssd1 vssd1 vccd1 vccd1 _6919_/A sky130_fd_sc_hd__and3_2
X_6847_ _6845_/A _6845_/B _6866_/A _6846_/Y vssd1 vssd1 vccd1 vccd1 _6849_/B sky130_fd_sc_hd__o2bb2a_1
X_6778_ _6969_/A _6778_/B vssd1 vssd1 vccd1 vccd1 _6783_/B sky130_fd_sc_hd__or2_4
X_5729_ _5765_/A _5765_/B _5727_/X vssd1 vssd1 vccd1 vccd1 _5732_/A sky130_fd_sc_hd__a21oi_4
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4060_ _8059_/Q _4080_/B _4096_/A vssd1 vssd1 vccd1 vccd1 _4061_/B sky130_fd_sc_hd__o21a_2
XFILLER_49_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7750_ _7750_/A _7764_/B vssd1 vssd1 vccd1 vccd1 _7750_/X sky130_fd_sc_hd__xor2_1
XFILLER_91_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4962_ _4931_/B _4925_/B _4925_/C vssd1 vssd1 vccd1 vccd1 _4963_/B sky130_fd_sc_hd__a21oi_2
X_6701_ _6749_/S _6701_/B vssd1 vssd1 vccd1 vccd1 _6701_/X sky130_fd_sc_hd__and2_1
X_7681_ _7682_/A _7682_/B vssd1 vssd1 vccd1 vccd1 _7683_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4893_ _4894_/A _4927_/B _4926_/A vssd1 vssd1 vccd1 vccd1 _4903_/A sky130_fd_sc_hd__o21ba_1
X_6632_ _6610_/A _6619_/Y _6608_/X vssd1 vssd1 vccd1 vccd1 _6632_/X sky130_fd_sc_hd__a21o_1
XFILLER_32_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6563_ _6577_/A _6641_/B vssd1 vssd1 vccd1 vccd1 _6578_/A sky130_fd_sc_hd__or2_2
XFILLER_20_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6494_ _6443_/A _6404_/B _6493_/X vssd1 vssd1 vccd1 vccd1 _6572_/A sky130_fd_sc_hd__o21ai_4
X_5514_ _5522_/A _5522_/B vssd1 vssd1 vccd1 vccd1 _5523_/A sky130_fd_sc_hd__nor2_4
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5445_ _5445_/A _7281_/C _5446_/B _5797_/A vssd1 vssd1 vccd1 vccd1 _5470_/A sky130_fd_sc_hd__or4_4
XFILLER_87_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5376_ _5377_/A _5377_/B vssd1 vssd1 vccd1 vccd1 _5376_/Y sky130_fd_sc_hd__nor2_1
X_7115_ _7114_/C _7007_/B _7128_/A vssd1 vssd1 vccd1 vccd1 _7161_/A sky130_fd_sc_hd__o21ba_4
Xfanout103 _7366_/B vssd1 vssd1 vccd1 vccd1 _5925_/A sky130_fd_sc_hd__buf_8
XFILLER_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4327_ _4547_/C _4275_/B _4275_/C _4260_/X vssd1 vssd1 vccd1 vccd1 _4327_/X sky130_fd_sc_hd__a31o_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout136 _4353_/Y vssd1 vssd1 vccd1 vccd1 _7306_/A sky130_fd_sc_hd__buf_8
Xfanout147 _4642_/A vssd1 vssd1 vccd1 vccd1 _7215_/A sky130_fd_sc_hd__clkbuf_4
Xfanout114 _4383_/X vssd1 vssd1 vccd1 vccd1 _5019_/A sky130_fd_sc_hd__buf_8
Xfanout125 _7025_/A vssd1 vssd1 vccd1 vccd1 _4411_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4258_ _6007_/A _6317_/A vssd1 vssd1 vccd1 vccd1 _4258_/X sky130_fd_sc_hd__or2_2
Xfanout169 _4081_/X vssd1 vssd1 vccd1 vccd1 _5986_/S sky130_fd_sc_hd__clkbuf_8
Xfanout158 _7261_/A vssd1 vssd1 vccd1 vccd1 _4602_/A sky130_fd_sc_hd__buf_6
X_7046_ _7371_/A _7046_/B _7045_/Y vssd1 vssd1 vccd1 vccd1 _7051_/A sky130_fd_sc_hd__or3b_2
XFILLER_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4189_ _8072_/Q _4189_/B vssd1 vssd1 vccd1 vccd1 _4192_/B sky130_fd_sc_hd__xnor2_4
XFILLER_27_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7948_ _8010_/Q _8009_/Q vssd1 vssd1 vccd1 vccd1 _7948_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7879_ _8038_/Q _7879_/B vssd1 vssd1 vccd1 vccd1 _7879_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5230_ _5230_/A _5230_/B vssd1 vssd1 vccd1 vccd1 _5232_/C sky130_fd_sc_hd__xnor2_1
XFILLER_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5161_ _5169_/A _5161_/B vssd1 vssd1 vccd1 vccd1 _5180_/B sky130_fd_sc_hd__and2_1
XFILLER_110_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4112_ _4088_/A _8052_/Q vssd1 vssd1 vccd1 vccd1 _4112_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_69_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5092_ _5092_/A vssd1 vssd1 vccd1 vccd1 _5093_/B sky130_fd_sc_hd__inv_2
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4043_ _8062_/Q _8061_/Q _4057_/B vssd1 vssd1 vccd1 vccd1 _5107_/B sky130_fd_sc_hd__or3_4
XFILLER_96_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7802_ _7793_/Y _7794_/X _7801_/X _7802_/B2 vssd1 vssd1 vccd1 vccd1 _7802_/Y sky130_fd_sc_hd__o22ai_4
X_5994_ _5995_/A _6021_/S vssd1 vssd1 vccd1 vccd1 _6027_/A sky130_fd_sc_hd__and2_2
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7733_ _7702_/X _7731_/B _7758_/A vssd1 vssd1 vccd1 vccd1 _7733_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4945_ _4945_/A _4945_/B vssd1 vssd1 vccd1 vccd1 _5054_/B sky130_fd_sc_hd__xnor2_2
X_7664_ _7647_/Y _7655_/X _7663_/X _7903_/B1 vssd1 vssd1 vccd1 vccd1 _7664_/X sky130_fd_sc_hd__a31o_2
X_4876_ _4876_/A _4876_/B vssd1 vssd1 vccd1 vccd1 _4878_/B sky130_fd_sc_hd__xnor2_4
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6615_ _6615_/A _6615_/B vssd1 vssd1 vccd1 vccd1 _6616_/D sky130_fd_sc_hd__and2_1
X_7595_ _7544_/A _7594_/Y _7889_/A vssd1 vssd1 vccd1 vccd1 _7597_/B sky130_fd_sc_hd__mux2_4
XFILLER_20_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6546_ _6546_/A vssd1 vssd1 vccd1 vccd1 _6547_/B sky130_fd_sc_hd__inv_2
XFILLER_106_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6477_ _6536_/A vssd1 vssd1 vccd1 vccd1 _6477_/Y sky130_fd_sc_hd__inv_2
X_5428_ _5422_/A _5422_/B _5420_/Y vssd1 vssd1 vccd1 vccd1 _5455_/A sky130_fd_sc_hd__o21ai_2
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5359_ _5360_/A _5360_/B vssd1 vssd1 vccd1 vccd1 _5359_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8078_ _8079_/CLK _8078_/D vssd1 vssd1 vccd1 vccd1 _8078_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7029_ _7031_/B _7031_/A vssd1 vssd1 vccd1 vccd1 _7029_/X sky130_fd_sc_hd__and2b_1
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _4730_/A _4730_/B vssd1 vssd1 vccd1 vccd1 _4730_/Y sky130_fd_sc_hd__nand2_1
X_4661_ _4660_/A _4660_/B _4676_/A vssd1 vssd1 vccd1 vccd1 _4665_/B sky130_fd_sc_hd__o21bai_2
X_6400_ _7269_/B _6999_/A _6445_/S vssd1 vssd1 vccd1 vccd1 _6400_/X sky130_fd_sc_hd__mux2_1
X_7380_ _7472_/A _7472_/B _7237_/X vssd1 vssd1 vccd1 vccd1 _7474_/B sky130_fd_sc_hd__a21oi_4
X_6331_ _7413_/A _6342_/B _6330_/Y _6559_/A vssd1 vssd1 vccd1 vccd1 _6343_/B sky130_fd_sc_hd__a22o_1
X_4592_ _4662_/A _5014_/A _4616_/C vssd1 vssd1 vccd1 vccd1 _4594_/B sky130_fd_sc_hd__o21ai_4
XFILLER_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6262_ _6009_/X _7639_/A _6262_/S vssd1 vssd1 vccd1 vccd1 _6262_/X sky130_fd_sc_hd__mux2_1
X_8001_ _8076_/Q _8020_/Q _8004_/S vssd1 vssd1 vccd1 vccd1 _8076_/D sky130_fd_sc_hd__mux2_1
X_6193_ _6193_/A _6200_/B _6200_/C vssd1 vssd1 vccd1 vccd1 _6193_/X sky130_fd_sc_hd__and3_1
X_5213_ _5265_/A _5214_/B vssd1 vssd1 vccd1 vccd1 _5213_/X sky130_fd_sc_hd__and2b_1
X_5144_ _5165_/B _6807_/A _5208_/A _5143_/X vssd1 vssd1 vccd1 vccd1 _5152_/B sky130_fd_sc_hd__o31a_2
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5075_ _5352_/A _5352_/B vssd1 vssd1 vccd1 vccd1 _5683_/A sky130_fd_sc_hd__nand2_2
X_4026_ _8015_/Q _8016_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _8016_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5977_ _5977_/A _5977_/B _5977_/C _5977_/D vssd1 vssd1 vccd1 vccd1 _5977_/Y sky130_fd_sc_hd__nand4_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7716_ _7616_/S _7582_/A _6631_/X vssd1 vssd1 vccd1 vccd1 _7717_/A sky130_fd_sc_hd__a21o_1
X_4928_ _4936_/A _4936_/B vssd1 vssd1 vccd1 vccd1 _4928_/X sky130_fd_sc_hd__and2b_1
X_7647_ _7644_/Y _7645_/X _7646_/Y vssd1 vssd1 vccd1 vccd1 _7647_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _4865_/A _4865_/B vssd1 vssd1 vccd1 vccd1 _4860_/C sky130_fd_sc_hd__and2_1
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7578_ _7577_/A _7576_/Y _7577_/Y _6268_/X vssd1 vssd1 vccd1 vccd1 _7578_/X sky130_fd_sc_hd__o211a_2
Xclkbuf_3_0__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _8075_/CLK sky130_fd_sc_hd__clkbuf_16
X_6529_ _6529_/A _6529_/B vssd1 vssd1 vccd1 vccd1 _6539_/B sky130_fd_sc_hd__xor2_4
XFILLER_109_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5900_ _5900_/A _5900_/B vssd1 vssd1 vccd1 vccd1 _5901_/B sky130_fd_sc_hd__and2_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6880_ _6881_/B _6881_/A vssd1 vssd1 vccd1 vccd1 _6887_/B sky130_fd_sc_hd__nand2b_1
XFILLER_61_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5831_ _5797_/A _5855_/B _5800_/D vssd1 vssd1 vccd1 vccd1 _5833_/B sky130_fd_sc_hd__o21ai_1
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5762_ _5762_/A _5794_/A vssd1 vssd1 vccd1 vccd1 _5788_/A sky130_fd_sc_hd__nand2_4
X_7501_ _7493_/X _7500_/A _7535_/A vssd1 vssd1 vccd1 vccd1 _7542_/B sky130_fd_sc_hd__mux2_2
X_4713_ _4685_/X _4686_/Y _4687_/A vssd1 vssd1 vccd1 vccd1 _4720_/B sky130_fd_sc_hd__o21bai_2
X_5693_ _5694_/A _5694_/B vssd1 vssd1 vccd1 vccd1 _5693_/X sky130_fd_sc_hd__and2b_1
X_7432_ _7424_/A _7424_/B _7430_/B vssd1 vssd1 vccd1 vccd1 _7438_/B sky130_fd_sc_hd__o21bai_4
X_4644_ _4644_/A _4644_/B vssd1 vssd1 vccd1 vccd1 _4648_/A sky130_fd_sc_hd__xor2_4
X_7363_ _7363_/A _7363_/B vssd1 vssd1 vccd1 vccd1 _7364_/B sky130_fd_sc_hd__and2_1
X_4575_ _4497_/A _4497_/B _4497_/C vssd1 vssd1 vccd1 vccd1 _4575_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6314_ _6349_/B _6766_/S _6311_/Y _6350_/A vssd1 vssd1 vccd1 vccd1 _6348_/B sky130_fd_sc_hd__a211o_4
X_7294_ _7294_/A _7294_/B _7294_/C vssd1 vssd1 vccd1 vccd1 _7299_/A sky130_fd_sc_hd__or3_1
X_6245_ _6254_/S _6245_/B _6245_/C vssd1 vssd1 vccd1 vccd1 _6245_/X sky130_fd_sc_hd__or3_1
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6176_ _5782_/A _6139_/B _6127_/A _6172_/X _6175_/X vssd1 vssd1 vccd1 vccd1 _6176_/X
+ sky130_fd_sc_hd__o221a_1
X_5127_ _5207_/A _5367_/A vssd1 vssd1 vccd1 vccd1 _6807_/A sky130_fd_sc_hd__or2_4
XFILLER_57_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5058_ _5058_/A _5247_/A vssd1 vssd1 vccd1 vccd1 _5058_/X sky130_fd_sc_hd__or2_1
XFILLER_29_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4009_ _8012_/Q _8011_/Q _8014_/Q _8013_/Q vssd1 vssd1 vccd1 vccd1 _4009_/X sky130_fd_sc_hd__or4_1
XFILLER_53_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_3 _4342_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4360_ _4360_/A _7261_/A vssd1 vssd1 vccd1 vccd1 _4360_/Y sky130_fd_sc_hd__nand2_2
X_4291_ _6311_/A vssd1 vssd1 vccd1 vccd1 _6349_/A sky130_fd_sc_hd__inv_2
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _6030_/A _6030_/B vssd1 vssd1 vccd1 vccd1 _6031_/B sky130_fd_sc_hd__xnor2_4
XFILLER_86_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7981_ _8017_/Q _8057_/Q _7990_/S vssd1 vssd1 vccd1 vccd1 _8057_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6932_ _6987_/B _6932_/B vssd1 vssd1 vccd1 vccd1 _6939_/B sky130_fd_sc_hd__or2_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6863_ _6863_/A _6863_/B vssd1 vssd1 vccd1 vccd1 _6888_/A sky130_fd_sc_hd__xor2_4
XFILLER_34_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5814_ _5815_/A _5815_/B _5815_/C vssd1 vssd1 vccd1 vccd1 _5847_/A sky130_fd_sc_hd__a21o_1
X_6794_ _6795_/A _6795_/B vssd1 vssd1 vccd1 vccd1 _6812_/B sky130_fd_sc_hd__and2_1
XFILLER_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5745_ _5745_/A _5908_/A _5908_/C vssd1 vssd1 vccd1 vccd1 _5751_/A sky130_fd_sc_hd__and3_4
X_5676_ _5676_/A _5676_/B vssd1 vssd1 vccd1 vccd1 _5677_/B sky130_fd_sc_hd__xnor2_4
XFILLER_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7415_ _7421_/B _7415_/B vssd1 vssd1 vccd1 vccd1 _7436_/B sky130_fd_sc_hd__xnor2_4
X_4627_ _4627_/A _4627_/B vssd1 vssd1 vccd1 vccd1 _4634_/A sky130_fd_sc_hd__nor2_2
XFILLER_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7346_ _7349_/A _7349_/B _7343_/X vssd1 vssd1 vccd1 vccd1 _7348_/B sky130_fd_sc_hd__a21oi_2
X_4558_ _7214_/A _4558_/B vssd1 vssd1 vccd1 vccd1 _4630_/C sky130_fd_sc_hd__or2_2
X_7277_ _7277_/A _7277_/B vssd1 vssd1 vccd1 vccd1 _7290_/A sky130_fd_sc_hd__xnor2_4
X_4489_ _4472_/A _4414_/X _4483_/X _4485_/Y vssd1 vssd1 vccd1 vccd1 _4489_/X sky130_fd_sc_hd__a31o_1
XFILLER_103_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6228_ _6228_/A _6228_/B vssd1 vssd1 vccd1 vccd1 _6228_/X sky130_fd_sc_hd__and2_1
XFILLER_103_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6159_ _6159_/A _6159_/B vssd1 vssd1 vccd1 vccd1 _6177_/B sky130_fd_sc_hd__xnor2_4
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput5 _8044_/Q vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__buf_4
XFILLER_110_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5530_ _5530_/A _5683_/B vssd1 vssd1 vccd1 vccd1 _5585_/A sky130_fd_sc_hd__or2_4
X_5461_ _5462_/A _5462_/B vssd1 vssd1 vccd1 vccd1 _5461_/X sky130_fd_sc_hd__and2b_1
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4412_ _4412_/A _4412_/B vssd1 vssd1 vccd1 vccd1 _4424_/B sky130_fd_sc_hd__nand2_1
X_7200_ _7319_/A _7195_/B _7195_/C vssd1 vssd1 vccd1 vccd1 _7201_/B sky130_fd_sc_hd__a21oi_2
X_5392_ _5394_/A _5394_/B vssd1 vssd1 vccd1 vccd1 _5392_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4343_ _4354_/A _4376_/A vssd1 vssd1 vccd1 vccd1 _4343_/Y sky130_fd_sc_hd__nor2_8
X_7131_ _7159_/A _7159_/B vssd1 vssd1 vccd1 vccd1 _7160_/A sky130_fd_sc_hd__nand2_2
XFILLER_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4274_ _4187_/B _4259_/B _4270_/X _4315_/B vssd1 vssd1 vccd1 vccd1 _4275_/C sky130_fd_sc_hd__a211o_1
X_7062_ _7063_/A _7063_/B vssd1 vssd1 vccd1 vccd1 _7091_/B sky130_fd_sc_hd__nand2_4
X_6013_ _7398_/A _6003_/Y _6008_/Y _6012_/Y _6084_/A vssd1 vssd1 vccd1 vccd1 _6088_/A
+ sky130_fd_sc_hd__o2111a_4
XFILLER_86_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7964_ _8047_/Q _8046_/Q _7964_/C vssd1 vssd1 vccd1 vccd1 _7970_/C sky130_fd_sc_hd__and3_2
XFILLER_82_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6915_ _7025_/A _7344_/B vssd1 vssd1 vccd1 vccd1 _6970_/B sky130_fd_sc_hd__nor2_1
X_7895_ _7895_/A _7895_/B _7895_/C vssd1 vssd1 vccd1 vccd1 _7921_/A sky130_fd_sc_hd__and3_2
X_6846_ _6866_/B vssd1 vssd1 vccd1 vccd1 _6846_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6777_ _6873_/A _7114_/B vssd1 vssd1 vccd1 vccd1 _6782_/A sky130_fd_sc_hd__nand2_4
XFILLER_10_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5728_ _5728_/A _5728_/B vssd1 vssd1 vccd1 vccd1 _5765_/B sky130_fd_sc_hd__xor2_4
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5659_ _5657_/A _5657_/B _5658_/Y vssd1 vssd1 vccd1 vccd1 _5708_/A sky130_fd_sc_hd__o21ai_4
XFILLER_117_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7329_ _7329_/A _7329_/B vssd1 vssd1 vccd1 vccd1 _7350_/A sky130_fd_sc_hd__xnor2_2
XFILLER_117_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4961_ _4995_/A _4995_/B _4953_/X vssd1 vssd1 vccd1 vccd1 _4965_/A sky130_fd_sc_hd__a21oi_4
X_6700_ _6687_/X _6699_/X _6753_/S vssd1 vssd1 vccd1 vccd1 _6701_/B sky130_fd_sc_hd__mux2_1
X_7680_ _7649_/B _7654_/B _7649_/A vssd1 vssd1 vccd1 vccd1 _7682_/B sky130_fd_sc_hd__a21oi_1
X_4892_ _4892_/A _4892_/B vssd1 vssd1 vccd1 vccd1 _4927_/B sky130_fd_sc_hd__xnor2_4
X_6631_ _7773_/A _7583_/S vssd1 vssd1 vccd1 vccd1 _6631_/X sky130_fd_sc_hd__and2_1
XFILLER_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6562_ _6562_/A _6562_/B vssd1 vssd1 vccd1 vccd1 _6562_/Y sky130_fd_sc_hd__nor2_1
X_6493_ _6492_/A _6440_/X _6483_/Y _6495_/B _6488_/B vssd1 vssd1 vccd1 vccd1 _6493_/X
+ sky130_fd_sc_hd__a221o_2
X_5513_ _5303_/Y _5566_/A _5563_/A _5563_/B vssd1 vssd1 vccd1 vccd1 _5522_/B sky130_fd_sc_hd__a22oi_4
X_5444_ _5411_/A _5411_/B _5409_/Y vssd1 vssd1 vccd1 vccd1 _5449_/A sky130_fd_sc_hd__o21a_2
X_5375_ _5375_/A _5375_/B vssd1 vssd1 vccd1 vccd1 _5377_/B sky130_fd_sc_hd__xnor2_4
Xfanout104 _7366_/B vssd1 vssd1 vccd1 vccd1 _5683_/B sky130_fd_sc_hd__buf_4
X_7114_ _7281_/B _7114_/B _7114_/C vssd1 vssd1 vccd1 vccd1 _7128_/A sky130_fd_sc_hd__and3_2
XFILLER_87_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4326_ _4322_/X _4323_/X _4324_/X vssd1 vssd1 vccd1 vccd1 _4326_/X sky130_fd_sc_hd__o21a_4
Xfanout137 _7294_/A vssd1 vssd1 vccd1 vccd1 _7371_/A sky130_fd_sc_hd__buf_4
Xfanout126 _6969_/A vssd1 vssd1 vccd1 vccd1 _7025_/A sky130_fd_sc_hd__buf_6
Xfanout115 _4383_/X vssd1 vssd1 vccd1 vccd1 _4551_/B sky130_fd_sc_hd__buf_6
XFILLER_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4257_ _4239_/Y _4547_/C _4245_/X _4256_/Y vssd1 vssd1 vccd1 vccd1 _6317_/A sky130_fd_sc_hd__a31o_4
Xfanout159 _7030_/A vssd1 vssd1 vccd1 vccd1 _7261_/A sky130_fd_sc_hd__buf_6
Xfanout148 _7012_/A vssd1 vssd1 vccd1 vccd1 _4642_/A sky130_fd_sc_hd__buf_4
X_7045_ _7045_/A _7045_/B vssd1 vssd1 vccd1 vccd1 _7045_/Y sky130_fd_sc_hd__xnor2_1
X_4188_ _8071_/Q _4175_/B _4211_/B vssd1 vssd1 vccd1 vccd1 _4189_/B sky130_fd_sc_hd__o21ai_4
XFILLER_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7947_ _8010_/Q _8009_/Q _7947_/C vssd1 vssd1 vccd1 vccd1 _7947_/X sky130_fd_sc_hd__or3_1
XFILLER_82_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7878_ _7923_/A _7869_/X _7877_/X _7903_/B1 vssd1 vssd1 vccd1 vccd1 _7878_/X sky130_fd_sc_hd__a211o_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6829_ _6828_/B _7392_/B _6828_/A vssd1 vssd1 vccd1 vccd1 _6830_/B sky130_fd_sc_hd__o21a_1
XFILLER_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5160_ _5160_/A _5160_/B vssd1 vssd1 vccd1 vccd1 _5161_/B sky130_fd_sc_hd__or2_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4111_ _4111_/A _6018_/A vssd1 vssd1 vccd1 vccd1 _4111_/X sky130_fd_sc_hd__or2_1
XFILLER_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5091_ _4920_/A _4751_/C _5090_/X vssd1 vssd1 vccd1 vccd1 _5092_/A sky130_fd_sc_hd__a21o_1
XFILLER_110_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4042_ _8060_/Q _8059_/Q _8058_/Q _4052_/B vssd1 vssd1 vccd1 vccd1 _4057_/B sky130_fd_sc_hd__or4_4
XFILLER_84_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7801_ _7801_/A _7874_/B vssd1 vssd1 vccd1 vccd1 _7801_/X sky130_fd_sc_hd__xor2_4
X_5993_ _6272_/A _5993_/B vssd1 vssd1 vccd1 vccd1 _6021_/S sky130_fd_sc_hd__nand2_1
X_7732_ _7702_/A _7757_/B _7757_/D vssd1 vssd1 vccd1 vccd1 _7758_/A sky130_fd_sc_hd__and3b_1
XFILLER_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4944_ _4945_/A _4945_/B vssd1 vssd1 vccd1 vccd1 _4944_/X sky130_fd_sc_hd__or2_1
X_7663_ _7663_/A _7663_/B vssd1 vssd1 vccd1 vccd1 _7663_/X sky130_fd_sc_hd__or2_1
X_4875_ _4998_/A _4947_/C vssd1 vssd1 vccd1 vccd1 _4876_/B sky130_fd_sc_hd__nand2_2
X_6614_ _6614_/A _6614_/B vssd1 vssd1 vccd1 vccd1 _6615_/B sky130_fd_sc_hd__or2_1
X_7594_ _7594_/A vssd1 vssd1 vccd1 vccd1 _7594_/Y sky130_fd_sc_hd__inv_2
X_6545_ _6545_/A _6545_/B vssd1 vssd1 vccd1 vccd1 _6546_/A sky130_fd_sc_hd__xor2_4
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6476_ _6476_/A _6476_/B vssd1 vssd1 vccd1 vccd1 _6536_/A sky130_fd_sc_hd__nand2_4
XFILLER_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5427_ _5556_/A _5556_/B vssd1 vssd1 vccd1 vccd1 _5612_/B sky130_fd_sc_hd__nand2_1
XFILLER_114_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5358_ _5358_/A _5358_/B vssd1 vssd1 vccd1 vccd1 _5360_/B sky130_fd_sc_hd__xnor2_4
X_8077_ _8077_/CLK _8077_/D vssd1 vssd1 vccd1 vccd1 _8077_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4309_ _6806_/A vssd1 vssd1 vccd1 vccd1 _5745_/A sky130_fd_sc_hd__inv_8
XFILLER_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5289_ _5054_/B _5054_/C _5054_/D _4944_/X vssd1 vssd1 vccd1 vccd1 _5290_/B sky130_fd_sc_hd__o31a_2
X_7028_ _5445_/A _7366_/B _7086_/A _7084_/A vssd1 vssd1 vccd1 vccd1 _7031_/B sky130_fd_sc_hd__o31a_4
XFILLER_47_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _4660_/A _4660_/B _4676_/A vssd1 vssd1 vccd1 vccd1 _4665_/A sky130_fd_sc_hd__or3b_2
XFILLER_9_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6330_ _6330_/A _6330_/B vssd1 vssd1 vccd1 vccd1 _6330_/Y sky130_fd_sc_hd__xnor2_1
X_4591_ _7247_/A _4988_/A vssd1 vssd1 vccd1 vccd1 _4616_/C sky130_fd_sc_hd__or2_2
XFILLER_115_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6261_ _6258_/X _6260_/Y _6544_/S vssd1 vssd1 vccd1 vccd1 _6267_/B sky130_fd_sc_hd__a21o_1
XFILLER_115_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8000_ _8075_/Q _8019_/Q _8004_/S vssd1 vssd1 vccd1 vccd1 _8075_/D sky130_fd_sc_hd__mux2_1
X_6192_ _6259_/A _6192_/B _6192_/C _6192_/D vssd1 vssd1 vccd1 vccd1 _6200_/C sky130_fd_sc_hd__or4_1
X_5212_ _5212_/A _5212_/B vssd1 vssd1 vccd1 vccd1 _5214_/B sky130_fd_sc_hd__xor2_4
X_5143_ _5128_/Y _5264_/A _5369_/A vssd1 vssd1 vccd1 vccd1 _5143_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5074_ _5074_/A _5074_/B _5074_/C vssd1 vssd1 vccd1 vccd1 _5352_/B sky130_fd_sc_hd__nand3_4
X_4025_ _8014_/Q _8015_/Q _7955_/S vssd1 vssd1 vccd1 vccd1 _8015_/D sky130_fd_sc_hd__mux2_1
XFILLER_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5976_ _5268_/A _5974_/X _5975_/X _5986_/S vssd1 vssd1 vccd1 vccd1 _5976_/Y sky130_fd_sc_hd__o31ai_4
XFILLER_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7715_ _6187_/X _7744_/A _7744_/B _7714_/Y _7918_/B vssd1 vssd1 vccd1 vccd1 _7715_/X
+ sky130_fd_sc_hd__a311o_1
X_4927_ _4927_/A _4927_/B vssd1 vssd1 vccd1 vccd1 _4936_/B sky130_fd_sc_hd__xnor2_4
XFILLER_40_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7646_ _7644_/Y _7645_/X _6269_/X vssd1 vssd1 vccd1 vccd1 _7646_/Y sky130_fd_sc_hd__a21oi_1
X_4858_ _4860_/B _4858_/B vssd1 vssd1 vccd1 vccd1 _4865_/B sky130_fd_sc_hd__nor2_2
XFILLER_20_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7577_ _7577_/A _7611_/B vssd1 vssd1 vccd1 vccd1 _7577_/Y sky130_fd_sc_hd__nand2_1
X_4789_ _4789_/A _4789_/B vssd1 vssd1 vccd1 vccd1 _4813_/A sky130_fd_sc_hd__nor2_1
XFILLER_119_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6528_ _6462_/Y _6505_/X _6544_/S vssd1 vssd1 vccd1 vccd1 _6529_/B sky130_fd_sc_hd__mux2_4
XFILLER_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6459_ _6479_/A _6541_/B _6479_/B vssd1 vssd1 vccd1 vccd1 _6460_/A sky130_fd_sc_hd__o21bai_4
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5830_ _7319_/B _5855_/A _5855_/B _5855_/C vssd1 vssd1 vccd1 vccd1 _5851_/A sky130_fd_sc_hd__or4_4
XFILLER_62_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5761_ _5761_/A _5762_/A _5761_/C vssd1 vssd1 vccd1 vccd1 _5794_/A sky130_fd_sc_hd__nand3_4
X_7500_ _7500_/A vssd1 vssd1 vccd1 vccd1 _7500_/Y sky130_fd_sc_hd__inv_2
X_4712_ _4712_/A _4712_/B vssd1 vssd1 vccd1 vccd1 _4730_/A sky130_fd_sc_hd__nor2_2
X_7431_ _7436_/A _7436_/B _7419_/B vssd1 vssd1 vccd1 vccd1 _7431_/X sky130_fd_sc_hd__a21bo_1
X_5692_ _5692_/A _5692_/B vssd1 vssd1 vccd1 vccd1 _5694_/B sky130_fd_sc_hd__xnor2_4
X_4643_ _4644_/A _4644_/B vssd1 vssd1 vccd1 vccd1 _4697_/A sky130_fd_sc_hd__nand2_1
X_7362_ _7374_/A _7374_/B vssd1 vssd1 vccd1 vccd1 _7362_/X sky130_fd_sc_hd__and2b_1
X_4574_ _4574_/A _4574_/B _4574_/C vssd1 vssd1 vccd1 vccd1 _4574_/X sky130_fd_sc_hd__or3_4
Xfanout6 _6166_/S vssd1 vssd1 vccd1 vccd1 _7639_/B sky130_fd_sc_hd__buf_6
X_6313_ _5973_/Y _5976_/Y _5977_/Y _6311_/A vssd1 vssd1 vccd1 vccd1 _6350_/A sky130_fd_sc_hd__o211a_1
X_7293_ _7293_/A _7293_/B vssd1 vssd1 vccd1 vccd1 _7294_/C sky130_fd_sc_hd__xnor2_1
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6244_ _6262_/S _6232_/Y _6243_/X _6139_/B vssd1 vssd1 vccd1 vccd1 _6245_/C sky130_fd_sc_hd__a22o_1
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6175_ _6175_/A _6175_/B _5970_/B vssd1 vssd1 vccd1 vccd1 _6175_/X sky130_fd_sc_hd__or3b_1
XFILLER_69_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5126_ _5207_/A _5367_/A vssd1 vssd1 vccd1 vccd1 _5166_/C sky130_fd_sc_hd__nor2_2
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5057_ _5247_/B _5247_/C _5058_/A _5247_/A vssd1 vssd1 vccd1 vccd1 _5071_/A sky130_fd_sc_hd__a211o_1
X_4008_ _8016_/Q _8015_/Q _8018_/Q _8017_/Q vssd1 vssd1 vccd1 vccd1 _4008_/X sky130_fd_sc_hd__or4_1
XFILLER_84_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5959_ _5959_/A _5959_/B _5959_/C vssd1 vssd1 vccd1 vccd1 _5960_/B sky130_fd_sc_hd__nand3_1
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7629_ _7629_/A _7629_/B vssd1 vssd1 vccd1 vccd1 _7630_/B sky130_fd_sc_hd__and2_1
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_4 _7294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4290_ _4286_/Y _4354_/B _4354_/A vssd1 vssd1 vccd1 vccd1 _6311_/A sky130_fd_sc_hd__mux2_8
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7980_ _8016_/Q _8056_/Q _7990_/S vssd1 vssd1 vccd1 vccd1 _8056_/D sky130_fd_sc_hd__mux2_1
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6931_ _6931_/A _6931_/B _6931_/C vssd1 vssd1 vccd1 vccd1 _6932_/B sky130_fd_sc_hd__nor3_1
X_6862_ _6862_/A _6862_/B vssd1 vssd1 vccd1 vccd1 _6893_/A sky130_fd_sc_hd__xnor2_2
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5813_ _5813_/A _5813_/B vssd1 vssd1 vccd1 vccd1 _5815_/C sky130_fd_sc_hd__xor2_1
X_6793_ _6812_/A _6793_/B vssd1 vssd1 vccd1 vccd1 _6795_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5744_ _5746_/B _5746_/A vssd1 vssd1 vccd1 vccd1 _5750_/A sky130_fd_sc_hd__and2b_1
X_5675_ _5676_/A _5676_/B vssd1 vssd1 vccd1 vccd1 _5675_/X sky130_fd_sc_hd__or2_1
X_7414_ _7419_/A _7766_/A vssd1 vssd1 vccd1 vccd1 _7415_/B sky130_fd_sc_hd__or2_4
X_4626_ _4585_/B _7281_/B _4989_/A _7247_/A vssd1 vssd1 vccd1 vccd1 _4627_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_116_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7345_ _7345_/A _7345_/B vssd1 vssd1 vccd1 vccd1 _7349_/B sky130_fd_sc_hd__xnor2_4
X_4557_ _4642_/A _5033_/A vssd1 vssd1 vccd1 vccd1 _4561_/A sky130_fd_sc_hd__nor2_2
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4488_ _4501_/A _4488_/B _4488_/C vssd1 vssd1 vccd1 vccd1 _4488_/X sky130_fd_sc_hd__and3_1
X_7276_ _7276_/A _7276_/B vssd1 vssd1 vccd1 vccd1 _7300_/A sky130_fd_sc_hd__xnor2_4
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6227_ _6227_/A _6227_/B vssd1 vssd1 vccd1 vccd1 _6240_/A sky130_fd_sc_hd__xnor2_4
XFILLER_106_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6158_ _6155_/A _6155_/B _5496_/Y vssd1 vssd1 vccd1 vccd1 _6159_/B sky130_fd_sc_hd__o21a_2
XFILLER_58_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _5683_/A _7046_/B vssd1 vssd1 vccd1 vccd1 _5111_/B sky130_fd_sc_hd__or2_4
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _6088_/A _6088_/B _6078_/C _6078_/B vssd1 vssd1 vccd1 vccd1 _6092_/A sky130_fd_sc_hd__o2bb2a_4
XFILLER_85_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5460_ _5441_/A _5441_/B _5434_/A vssd1 vssd1 vccd1 vccd1 _5462_/B sky130_fd_sc_hd__a21o_2
XFILLER_117_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4411_ _4411_/A _4411_/B vssd1 vssd1 vccd1 vccd1 _4509_/A sky130_fd_sc_hd__or2_4
X_5391_ _5391_/A _5391_/B vssd1 vssd1 vccd1 vccd1 _5394_/B sky130_fd_sc_hd__xnor2_4
XFILLER_113_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4342_ _6034_/A _4266_/A _4266_/B _4267_/X _4354_/A vssd1 vssd1 vccd1 vccd1 _4342_/X
+ sky130_fd_sc_hd__a311o_4
X_7130_ _7130_/A _7130_/B vssd1 vssd1 vccd1 vccd1 _7159_/B sky130_fd_sc_hd__xnor2_1
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4273_ _4180_/Y _4259_/B _4271_/X _4219_/Y vssd1 vssd1 vccd1 vccd1 _4275_/B sky130_fd_sc_hd__a211o_1
X_7061_ _7112_/A _7112_/B vssd1 vssd1 vccd1 vccd1 _7063_/B sky130_fd_sc_hd__and2_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6012_ _6012_/A _6012_/B vssd1 vssd1 vccd1 vccd1 _6012_/Y sky130_fd_sc_hd__nor2_1
.ends

