magic
tech sky130B
magscale 1 2
timestamp 1680008312
<< viali >>
rect 12173 21573 12207 21607
rect 15301 21573 15335 21607
rect 20453 21573 20487 21607
rect 15209 21505 15243 21539
rect 15485 21505 15519 21539
rect 19625 21505 19659 21539
rect 19809 21437 19843 21471
rect 12357 21369 12391 21403
rect 15485 21301 15519 21335
rect 19441 21301 19475 21335
rect 20361 21301 20395 21335
rect 2789 21097 2823 21131
rect 16129 21097 16163 21131
rect 4353 21029 4387 21063
rect 10241 21029 10275 21063
rect 13645 21029 13679 21063
rect 16497 21029 16531 21063
rect 17325 21029 17359 21063
rect 11529 20961 11563 20995
rect 17969 20961 18003 20995
rect 2053 20893 2087 20927
rect 2145 20893 2179 20927
rect 5466 20893 5500 20927
rect 5733 20893 5767 20927
rect 8585 20893 8619 20927
rect 11805 20893 11839 20927
rect 12265 20893 12299 20927
rect 15301 20893 15335 20927
rect 15485 20893 15519 20927
rect 15669 20893 15703 20927
rect 16313 20893 16347 20927
rect 16589 20893 16623 20927
rect 17049 20893 17083 20927
rect 18245 20893 18279 20927
rect 19717 20893 19751 20927
rect 20085 20893 20119 20927
rect 2973 20825 3007 20859
rect 3157 20825 3191 20859
rect 8340 20825 8374 20859
rect 9137 20825 9171 20859
rect 9321 20825 9355 20859
rect 12532 20825 12566 20859
rect 17325 20825 17359 20859
rect 2329 20757 2363 20791
rect 7205 20757 7239 20791
rect 9505 20757 9539 20791
rect 17141 20757 17175 20791
rect 18889 20757 18923 20791
rect 1869 20553 1903 20587
rect 4353 20553 4387 20587
rect 8401 20553 8435 20587
rect 13829 20553 13863 20587
rect 18061 20553 18095 20587
rect 18705 20553 18739 20587
rect 2053 20485 2087 20519
rect 9956 20485 9990 20519
rect 12716 20485 12750 20519
rect 15761 20485 15795 20519
rect 1777 20417 1811 20451
rect 2697 20417 2731 20451
rect 5466 20417 5500 20451
rect 7021 20417 7055 20451
rect 7277 20417 7311 20451
rect 14473 20417 14507 20451
rect 15301 20417 15335 20451
rect 15945 20417 15979 20451
rect 16221 20417 16255 20451
rect 17049 20417 17083 20451
rect 17233 20417 17267 20451
rect 18889 20417 18923 20451
rect 19165 20417 19199 20451
rect 2513 20349 2547 20383
rect 5733 20349 5767 20383
rect 9689 20349 9723 20383
rect 12449 20349 12483 20383
rect 18981 20349 19015 20383
rect 19073 20349 19107 20383
rect 2053 20213 2087 20247
rect 2881 20213 2915 20247
rect 11069 20213 11103 20247
rect 16129 20213 16163 20247
rect 3065 20009 3099 20043
rect 16037 20009 16071 20043
rect 2053 19941 2087 19975
rect 4445 19941 4479 19975
rect 13553 19941 13587 19975
rect 1961 19873 1995 19907
rect 14657 19873 14691 19907
rect 2237 19805 2271 19839
rect 5558 19805 5592 19839
rect 5825 19805 5859 19839
rect 12173 19805 12207 19839
rect 15577 19805 15611 19839
rect 3249 19737 3283 19771
rect 3433 19737 3467 19771
rect 12440 19737 12474 19771
rect 14381 19737 14415 19771
rect 15209 19737 15243 19771
rect 15393 19737 15427 19771
rect 16221 19737 16255 19771
rect 16405 19737 16439 19771
rect 2421 19669 2455 19703
rect 2513 19465 2547 19499
rect 10885 19465 10919 19499
rect 16865 19465 16899 19499
rect 12348 19397 12382 19431
rect 14657 19397 14691 19431
rect 18889 19397 18923 19431
rect 2145 19329 2179 19363
rect 2329 19329 2363 19363
rect 5742 19329 5776 19363
rect 6009 19329 6043 19363
rect 6929 19329 6963 19363
rect 7185 19329 7219 19363
rect 9772 19329 9806 19363
rect 14841 19329 14875 19363
rect 16129 19329 16163 19363
rect 16313 19329 16347 19363
rect 17233 19329 17267 19363
rect 19073 19329 19107 19363
rect 19533 19329 19567 19363
rect 19717 19329 19751 19363
rect 9505 19261 9539 19295
rect 12081 19261 12115 19295
rect 15025 19261 15059 19295
rect 17049 19261 17083 19295
rect 17141 19261 17175 19295
rect 17325 19261 17359 19295
rect 13461 19193 13495 19227
rect 16129 19193 16163 19227
rect 4629 19125 4663 19159
rect 8309 19125 8343 19159
rect 18705 19125 18739 19159
rect 19625 19125 19659 19159
rect 4537 18921 4571 18955
rect 8401 18921 8435 18955
rect 10701 18921 10735 18955
rect 16589 18921 16623 18955
rect 5917 18785 5951 18819
rect 20361 18785 20395 18819
rect 3065 18717 3099 18751
rect 3249 18717 3283 18751
rect 8125 18717 8159 18751
rect 8217 18717 8251 18751
rect 9321 18717 9355 18751
rect 9588 18717 9622 18751
rect 12081 18717 12115 18751
rect 12357 18717 12391 18751
rect 16865 18717 16899 18751
rect 18705 18717 18739 18751
rect 18889 18717 18923 18751
rect 19441 18717 19475 18751
rect 19625 18717 19659 18751
rect 5650 18649 5684 18683
rect 16589 18649 16623 18683
rect 20913 18649 20947 18683
rect 3433 18581 3467 18615
rect 13645 18581 13679 18615
rect 16773 18581 16807 18615
rect 18521 18581 18555 18615
rect 19625 18581 19659 18615
rect 4077 18377 4111 18411
rect 15301 18377 15335 18411
rect 5650 18309 5684 18343
rect 7634 18309 7668 18343
rect 18521 18309 18555 18343
rect 18705 18309 18739 18343
rect 19441 18309 19475 18343
rect 1777 18241 1811 18275
rect 1961 18241 1995 18275
rect 2421 18241 2455 18275
rect 3709 18241 3743 18275
rect 3893 18241 3927 18275
rect 5917 18241 5951 18275
rect 7389 18241 7423 18275
rect 15485 18241 15519 18275
rect 15761 18241 15795 18275
rect 19349 18241 19383 18275
rect 19533 18241 19567 18275
rect 1869 18173 1903 18207
rect 18797 18173 18831 18207
rect 4537 18105 4571 18139
rect 8769 18105 8803 18139
rect 2513 18037 2547 18071
rect 15669 18037 15703 18071
rect 18245 18037 18279 18071
rect 2973 17833 3007 17867
rect 5733 17833 5767 17867
rect 11713 17833 11747 17867
rect 15485 17833 15519 17867
rect 1961 17629 1995 17663
rect 2237 17629 2271 17663
rect 3065 17629 3099 17663
rect 14841 17629 14875 17663
rect 15025 17629 15059 17663
rect 15761 17629 15795 17663
rect 16221 17629 16255 17663
rect 19441 17629 19475 17663
rect 2053 17561 2087 17595
rect 7021 17561 7055 17595
rect 10425 17561 10459 17595
rect 15485 17561 15519 17595
rect 19625 17561 19659 17595
rect 19809 17561 19843 17595
rect 2421 17493 2455 17527
rect 14933 17493 14967 17527
rect 15669 17493 15703 17527
rect 16313 17493 16347 17527
rect 1961 17289 1995 17323
rect 9934 17221 9968 17255
rect 14289 17221 14323 17255
rect 18521 17221 18555 17255
rect 19349 17221 19383 17255
rect 2329 17153 2363 17187
rect 3065 17153 3099 17187
rect 3249 17153 3283 17187
rect 5742 17153 5776 17187
rect 6009 17153 6043 17187
rect 7389 17153 7423 17187
rect 7645 17153 7679 17187
rect 12633 17153 12667 17187
rect 12909 17153 12943 17187
rect 16865 17153 16899 17187
rect 17601 17153 17635 17187
rect 18981 17153 19015 17187
rect 19441 17153 19475 17187
rect 20177 17153 20211 17187
rect 20361 17153 20395 17187
rect 20821 17153 20855 17187
rect 21005 17153 21039 17187
rect 2421 17085 2455 17119
rect 2605 17085 2639 17119
rect 9689 17085 9723 17119
rect 17693 17085 17727 17119
rect 19717 17085 19751 17119
rect 20269 17085 20303 17119
rect 11069 17017 11103 17051
rect 16957 17017 16991 17051
rect 3157 16949 3191 16983
rect 4629 16949 4663 16983
rect 8769 16949 8803 16983
rect 20913 16949 20947 16983
rect 16497 16745 16531 16779
rect 18705 16745 18739 16779
rect 11161 16677 11195 16711
rect 19993 16677 20027 16711
rect 3433 16609 3467 16643
rect 4537 16609 4571 16643
rect 7021 16609 7055 16643
rect 9781 16609 9815 16643
rect 12081 16609 12115 16643
rect 16129 16609 16163 16643
rect 16221 16609 16255 16643
rect 17509 16609 17543 16643
rect 17693 16609 17727 16643
rect 18429 16609 18463 16643
rect 2237 16541 2271 16575
rect 2421 16541 2455 16575
rect 3065 16541 3099 16575
rect 3249 16541 3283 16575
rect 7277 16541 7311 16575
rect 15209 16541 15243 16575
rect 15301 16541 15335 16575
rect 15853 16541 15887 16575
rect 16037 16541 16071 16575
rect 16313 16541 16347 16575
rect 17141 16541 17175 16575
rect 17417 16541 17451 16575
rect 18245 16541 18279 16575
rect 18337 16541 18371 16575
rect 18521 16541 18555 16575
rect 19441 16541 19475 16575
rect 19533 16541 19567 16575
rect 19717 16541 19751 16575
rect 19809 16541 19843 16575
rect 4782 16473 4816 16507
rect 10048 16473 10082 16507
rect 12326 16473 12360 16507
rect 2421 16405 2455 16439
rect 5917 16405 5951 16439
rect 8401 16405 8435 16439
rect 13461 16405 13495 16439
rect 1777 16201 1811 16235
rect 9321 16133 9355 16167
rect 19073 16133 19107 16167
rect 1869 16065 1903 16099
rect 2053 16065 2087 16099
rect 2881 16065 2915 16099
rect 3433 16065 3467 16099
rect 3617 16065 3651 16099
rect 16957 16065 16991 16099
rect 17141 16065 17175 16099
rect 17233 16065 17267 16099
rect 17417 16065 17451 16099
rect 18705 16065 18739 16099
rect 19441 16065 19475 16099
rect 19533 16065 19567 16099
rect 19901 16065 19935 16099
rect 1593 15997 1627 16031
rect 12633 15997 12667 16031
rect 12909 15997 12943 16031
rect 18521 15997 18555 16031
rect 2697 15929 2731 15963
rect 17049 15929 17083 15963
rect 3525 15861 3559 15895
rect 10609 15861 10643 15895
rect 14197 15861 14231 15895
rect 2145 15657 2179 15691
rect 17049 15657 17083 15691
rect 17233 15657 17267 15691
rect 19717 15589 19751 15623
rect 2329 15521 2363 15555
rect 2421 15521 2455 15555
rect 2605 15521 2639 15555
rect 2513 15453 2547 15487
rect 9597 15453 9631 15487
rect 9853 15453 9887 15487
rect 12357 15453 12391 15487
rect 15945 15453 15979 15487
rect 19441 15453 19475 15487
rect 12624 15385 12658 15419
rect 16497 15385 16531 15419
rect 17417 15385 17451 15419
rect 19717 15385 19751 15419
rect 10977 15317 11011 15351
rect 13737 15317 13771 15351
rect 17217 15317 17251 15351
rect 19533 15317 19567 15351
rect 3801 15113 3835 15147
rect 15301 15113 15335 15147
rect 17233 15113 17267 15147
rect 18797 15113 18831 15147
rect 20085 15113 20119 15147
rect 2973 15045 3007 15079
rect 7910 15045 7944 15079
rect 2329 14977 2363 15011
rect 2513 14977 2547 15011
rect 2789 14977 2823 15011
rect 3525 14977 3559 15011
rect 4701 14977 4735 15011
rect 12624 14977 12658 15011
rect 15485 14977 15519 15011
rect 15577 14977 15611 15011
rect 15761 14977 15795 15011
rect 15853 14977 15887 15011
rect 16865 14977 16899 15011
rect 18521 14977 18555 15011
rect 19349 14977 19383 15011
rect 20085 14977 20119 15011
rect 4445 14909 4479 14943
rect 7665 14909 7699 14943
rect 12357 14909 12391 14943
rect 16957 14909 16991 14943
rect 19257 14909 19291 14943
rect 20361 14909 20395 14943
rect 20177 14841 20211 14875
rect 5825 14773 5859 14807
rect 9045 14773 9079 14807
rect 13737 14773 13771 14807
rect 16865 14773 16899 14807
rect 2237 14569 2271 14603
rect 2329 14569 2363 14603
rect 19625 14569 19659 14603
rect 19809 14569 19843 14603
rect 15853 14501 15887 14535
rect 2421 14433 2455 14467
rect 16865 14433 16899 14467
rect 2145 14365 2179 14399
rect 5641 14365 5675 14399
rect 8125 14365 8159 14399
rect 9505 14365 9539 14399
rect 9781 14365 9815 14399
rect 12357 14365 12391 14399
rect 12624 14365 12658 14399
rect 16129 14365 16163 14399
rect 16773 14365 16807 14399
rect 16957 14365 16991 14399
rect 17049 14365 17083 14399
rect 17601 14365 17635 14399
rect 17785 14365 17819 14399
rect 18429 14365 18463 14399
rect 18613 14365 18647 14399
rect 5374 14297 5408 14331
rect 7858 14297 7892 14331
rect 15853 14297 15887 14331
rect 19441 14297 19475 14331
rect 4261 14229 4295 14263
rect 6745 14229 6779 14263
rect 11069 14229 11103 14263
rect 13737 14229 13771 14263
rect 16037 14229 16071 14263
rect 16589 14229 16623 14263
rect 17601 14229 17635 14263
rect 18521 14229 18555 14263
rect 19651 14229 19685 14263
rect 2421 14025 2455 14059
rect 15485 14025 15519 14059
rect 2329 13889 2363 13923
rect 4261 13889 4295 13923
rect 4528 13889 4562 13923
rect 7297 13889 7331 13923
rect 7553 13889 7587 13923
rect 10048 13889 10082 13923
rect 12808 13889 12842 13923
rect 14657 13889 14691 13923
rect 14749 13889 14783 13923
rect 14933 13889 14967 13923
rect 15577 13889 15611 13923
rect 15853 13889 15887 13923
rect 17049 13889 17083 13923
rect 18705 13889 18739 13923
rect 19901 13889 19935 13923
rect 9781 13821 9815 13855
rect 12541 13821 12575 13855
rect 15393 13821 15427 13855
rect 16221 13821 16255 13855
rect 16957 13821 16991 13855
rect 18889 13821 18923 13855
rect 18981 13821 19015 13855
rect 19625 13821 19659 13855
rect 13921 13753 13955 13787
rect 14933 13753 14967 13787
rect 5641 13685 5675 13719
rect 8677 13685 8711 13719
rect 11161 13685 11195 13719
rect 18521 13685 18555 13719
rect 5733 13481 5767 13515
rect 19717 13413 19751 13447
rect 18245 13345 18279 13379
rect 19993 13345 20027 13379
rect 7021 13277 7055 13311
rect 10425 13277 10459 13311
rect 16405 13277 16439 13311
rect 16497 13277 16531 13311
rect 18061 13277 18095 13311
rect 18613 13277 18647 13311
rect 12173 13209 12207 13243
rect 16773 13209 16807 13243
rect 18797 13209 18831 13243
rect 16221 13141 16255 13175
rect 16589 13141 16623 13175
rect 18705 13141 18739 13175
rect 19533 13141 19567 13175
rect 16037 12937 16071 12971
rect 19901 12937 19935 12971
rect 8208 12869 8242 12903
rect 12900 12869 12934 12903
rect 19809 12869 19843 12903
rect 5282 12801 5316 12835
rect 5549 12801 5583 12835
rect 10048 12801 10082 12835
rect 16037 12801 16071 12835
rect 19257 12801 19291 12835
rect 7941 12733 7975 12767
rect 9781 12733 9815 12767
rect 12633 12733 12667 12767
rect 15761 12733 15795 12767
rect 18889 12733 18923 12767
rect 15945 12665 15979 12699
rect 19092 12665 19126 12699
rect 4169 12597 4203 12631
rect 9321 12597 9355 12631
rect 11161 12597 11195 12631
rect 14013 12597 14047 12631
rect 18613 12597 18647 12631
rect 18981 12597 19015 12631
rect 15669 12393 15703 12427
rect 16221 12325 16255 12359
rect 11345 12257 11379 12291
rect 18613 12257 18647 12291
rect 19441 12257 19475 12291
rect 19625 12257 19659 12291
rect 19901 12257 19935 12291
rect 2237 12189 2271 12223
rect 2421 12189 2455 12223
rect 2513 12189 2547 12223
rect 2605 12189 2639 12223
rect 5641 12189 5675 12223
rect 6377 12189 6411 12223
rect 9229 12189 9263 12223
rect 9505 12189 9539 12223
rect 14289 12189 14323 12223
rect 16129 12189 16163 12223
rect 16405 12189 16439 12223
rect 18153 12189 18187 12223
rect 18705 12189 18739 12223
rect 19993 12189 20027 12223
rect 2881 12121 2915 12155
rect 5374 12121 5408 12155
rect 6644 12121 6678 12155
rect 11590 12121 11624 12155
rect 14534 12121 14568 12155
rect 16865 12121 16899 12155
rect 4261 12053 4295 12087
rect 7757 12053 7791 12087
rect 10609 12053 10643 12087
rect 12725 12053 12759 12087
rect 18337 12053 18371 12087
rect 2513 11849 2547 11883
rect 2973 11849 3007 11883
rect 16865 11849 16899 11883
rect 19533 11849 19567 11883
rect 2329 11713 2363 11747
rect 2973 11713 3007 11747
rect 3157 11713 3191 11747
rect 4261 11713 4295 11747
rect 4517 11713 4551 11747
rect 8309 11713 8343 11747
rect 8576 11713 8610 11747
rect 12633 11713 12667 11747
rect 12900 11713 12934 11747
rect 15669 11713 15703 11747
rect 16129 11713 16163 11747
rect 17049 11713 17083 11747
rect 17233 11713 17267 11747
rect 18337 11713 18371 11747
rect 18981 11713 19015 11747
rect 19165 11713 19199 11747
rect 19625 11713 19659 11747
rect 2145 11645 2179 11679
rect 17325 11645 17359 11679
rect 15761 11577 15795 11611
rect 5641 11509 5675 11543
rect 9689 11509 9723 11543
rect 14013 11509 14047 11543
rect 7665 11237 7699 11271
rect 16037 11237 16071 11271
rect 6285 11169 6319 11203
rect 15761 11169 15795 11203
rect 16221 11169 16255 11203
rect 18183 11101 18217 11135
rect 18337 11101 18371 11135
rect 6530 11033 6564 11067
rect 17969 11033 18003 11067
rect 2145 10761 2179 10795
rect 2973 10761 3007 10795
rect 3525 10761 3559 10795
rect 8401 10761 8435 10795
rect 13369 10761 13403 10795
rect 1869 10693 1903 10727
rect 7297 10693 7331 10727
rect 2145 10625 2179 10659
rect 2789 10625 2823 10659
rect 3065 10625 3099 10659
rect 3525 10625 3559 10659
rect 5733 10625 5767 10659
rect 6561 10625 6595 10659
rect 6745 10625 6779 10659
rect 7205 10625 7239 10659
rect 7573 10625 7607 10659
rect 8309 10625 8343 10659
rect 8493 10625 8527 10659
rect 13093 10625 13127 10659
rect 14013 10625 14047 10659
rect 15853 10625 15887 10659
rect 16129 10625 16163 10659
rect 18245 10625 18279 10659
rect 18429 10625 18463 10659
rect 18613 10625 18647 10659
rect 18705 10625 18739 10659
rect 19809 10625 19843 10659
rect 3801 10557 3835 10591
rect 6009 10557 6043 10591
rect 7389 10557 7423 10591
rect 13369 10557 13403 10591
rect 15945 10557 15979 10591
rect 19717 10557 19751 10591
rect 2053 10489 2087 10523
rect 2789 10489 2823 10523
rect 3617 10489 3651 10523
rect 5825 10489 5859 10523
rect 13921 10489 13955 10523
rect 18521 10489 18555 10523
rect 19441 10489 19475 10523
rect 5917 10421 5951 10455
rect 6653 10421 6687 10455
rect 7573 10421 7607 10455
rect 13185 10421 13219 10455
rect 15669 10421 15703 10455
rect 16129 10421 16163 10455
rect 18981 10421 19015 10455
rect 2145 10217 2179 10251
rect 2329 10217 2363 10251
rect 4169 10217 4203 10251
rect 6377 10217 6411 10251
rect 9137 10217 9171 10251
rect 10333 10217 10367 10251
rect 11253 10217 11287 10251
rect 11621 10217 11655 10251
rect 12081 10217 12115 10251
rect 12265 10217 12299 10251
rect 13185 10217 13219 10251
rect 14289 10217 14323 10251
rect 18337 10217 18371 10251
rect 20085 10217 20119 10251
rect 3341 10149 3375 10183
rect 4353 10149 4387 10183
rect 17233 10149 17267 10183
rect 17969 10149 18003 10183
rect 18429 10149 18463 10183
rect 2789 10081 2823 10115
rect 7481 10081 7515 10115
rect 8033 10081 8067 10115
rect 9689 10081 9723 10115
rect 10425 10081 10459 10115
rect 11529 10081 11563 10115
rect 13737 10081 13771 10115
rect 14933 10081 14967 10115
rect 15853 10081 15887 10115
rect 16589 10081 16623 10115
rect 16773 10081 16807 10115
rect 18521 10081 18555 10115
rect 18613 10081 18647 10115
rect 3065 10013 3099 10047
rect 4077 10013 4111 10047
rect 4261 10013 4295 10047
rect 4445 10013 4479 10047
rect 5733 10013 5767 10047
rect 5917 10013 5951 10047
rect 6009 10013 6043 10047
rect 6101 10013 6135 10047
rect 6929 10013 6963 10047
rect 7021 10013 7055 10047
rect 7665 10013 7699 10047
rect 9597 10013 9631 10047
rect 10517 10013 10551 10047
rect 11621 10013 11655 10047
rect 13461 10013 13495 10047
rect 13553 10013 13587 10047
rect 14470 10013 14504 10047
rect 14841 10013 14875 10047
rect 15485 10013 15519 10047
rect 15761 10013 15795 10047
rect 19441 10013 19475 10047
rect 19625 10013 19659 10047
rect 19717 10013 19751 10047
rect 19809 10013 19843 10047
rect 1961 9945 1995 9979
rect 2973 9945 3007 9979
rect 4721 9945 4755 9979
rect 7849 9945 7883 9979
rect 10793 9945 10827 9979
rect 12249 9945 12283 9979
rect 12449 9945 12483 9979
rect 13369 9945 13403 9979
rect 16865 9945 16899 9979
rect 2171 9877 2205 9911
rect 3157 9877 3191 9911
rect 7757 9877 7791 9911
rect 9505 9877 9539 9911
rect 10701 9877 10735 9911
rect 14473 9877 14507 9911
rect 15945 9877 15979 9911
rect 1869 9673 1903 9707
rect 6729 9673 6763 9707
rect 8217 9673 8251 9707
rect 9229 9673 9263 9707
rect 2053 9605 2087 9639
rect 5641 9605 5675 9639
rect 6929 9605 6963 9639
rect 7941 9605 7975 9639
rect 8309 9605 8343 9639
rect 10609 9605 10643 9639
rect 11897 9605 11931 9639
rect 13553 9605 13587 9639
rect 16313 9605 16347 9639
rect 1777 9537 1811 9571
rect 5825 9537 5859 9571
rect 8033 9537 8067 9571
rect 9137 9537 9171 9571
rect 9321 9537 9355 9571
rect 10793 9537 10827 9571
rect 10885 9537 10919 9571
rect 11713 9537 11747 9571
rect 11989 9537 12023 9571
rect 13277 9537 13311 9571
rect 13737 9537 13771 9571
rect 15945 9537 15979 9571
rect 16221 9537 16255 9571
rect 18797 9537 18831 9571
rect 18981 9537 19015 9571
rect 8125 9469 8159 9503
rect 15853 9469 15887 9503
rect 18521 9469 18555 9503
rect 2053 9401 2087 9435
rect 6009 9401 6043 9435
rect 10609 9401 10643 9435
rect 11713 9401 11747 9435
rect 6561 9333 6595 9367
rect 6745 9333 6779 9367
rect 15669 9333 15703 9367
rect 2053 9129 2087 9163
rect 7665 9129 7699 9163
rect 13185 9129 13219 9163
rect 13369 9129 13403 9163
rect 15761 9129 15795 9163
rect 16129 9129 16163 9163
rect 18889 9129 18923 9163
rect 2421 8993 2455 9027
rect 4445 8993 4479 9027
rect 7297 8993 7331 9027
rect 18429 8993 18463 9027
rect 2237 8925 2271 8959
rect 4261 8925 4295 8959
rect 7481 8925 7515 8959
rect 12449 8925 12483 8959
rect 12633 8925 12667 8959
rect 15945 8925 15979 8959
rect 16313 8925 16347 8959
rect 18521 8925 18555 8959
rect 18705 8925 18739 8959
rect 13353 8857 13387 8891
rect 13553 8857 13587 8891
rect 4077 8789 4111 8823
rect 12541 8789 12575 8823
rect 4261 8585 4295 8619
rect 6830 8585 6864 8619
rect 8493 8585 8527 8619
rect 10701 8585 10735 8619
rect 11897 8585 11931 8619
rect 12081 8585 12115 8619
rect 17877 8585 17911 8619
rect 11161 8517 11195 8551
rect 2973 8449 3007 8483
rect 3617 8449 3651 8483
rect 3801 8449 3835 8483
rect 3893 8449 3927 8483
rect 3985 8449 4019 8483
rect 4905 8449 4939 8483
rect 6653 8449 6687 8483
rect 6745 8449 6779 8483
rect 6929 8449 6963 8483
rect 7481 8449 7515 8483
rect 7573 8449 7607 8483
rect 7757 8449 7791 8483
rect 8769 8449 8803 8483
rect 9689 8449 9723 8483
rect 12909 8449 12943 8483
rect 13093 8449 13127 8483
rect 13829 8449 13863 8483
rect 14473 8449 14507 8483
rect 14657 8449 14691 8483
rect 15669 8449 15703 8483
rect 16129 8449 16163 8483
rect 17785 8449 17819 8483
rect 17969 8449 18003 8483
rect 18429 8449 18463 8483
rect 3065 8381 3099 8415
rect 4721 8381 4755 8415
rect 9321 8381 9355 8415
rect 9413 8381 9447 8415
rect 9781 8381 9815 8415
rect 14565 8381 14599 8415
rect 15761 8381 15795 8415
rect 19165 8381 19199 8415
rect 19625 8381 19659 8415
rect 7665 8313 7699 8347
rect 7941 8313 7975 8347
rect 10793 8313 10827 8347
rect 12449 8313 12483 8347
rect 13001 8313 13035 8347
rect 18613 8313 18647 8347
rect 19349 8313 19383 8347
rect 5089 8245 5123 8279
rect 9965 8245 9999 8279
rect 12081 8245 12115 8279
rect 13921 8245 13955 8279
rect 3249 8041 3283 8075
rect 3433 8041 3467 8075
rect 4077 8041 4111 8075
rect 7389 8041 7423 8075
rect 7573 8041 7607 8075
rect 8493 8041 8527 8075
rect 9781 8041 9815 8075
rect 10977 8041 11011 8075
rect 13645 8041 13679 8075
rect 15669 8041 15703 8075
rect 18613 8041 18647 8075
rect 19625 8041 19659 8075
rect 8401 7973 8435 8007
rect 13553 7973 13587 8007
rect 7021 7905 7055 7939
rect 9873 7905 9907 7939
rect 12541 7905 12575 7939
rect 13461 7905 13495 7939
rect 4445 7837 4479 7871
rect 5273 7837 5307 7871
rect 5457 7837 5491 7871
rect 5549 7837 5583 7871
rect 6009 7837 6043 7871
rect 6285 7837 6319 7871
rect 6377 7837 6411 7871
rect 8033 7837 8067 7871
rect 9652 7837 9686 7871
rect 10885 7837 10919 7871
rect 11253 7837 11287 7871
rect 13737 7837 13771 7871
rect 14473 7837 14507 7871
rect 14565 7837 14599 7871
rect 16313 7837 16347 7871
rect 16497 7837 16531 7871
rect 16957 7837 16991 7871
rect 17141 7837 17175 7871
rect 17417 7837 17451 7871
rect 18061 7837 18095 7871
rect 18429 7837 18463 7871
rect 19625 7837 19659 7871
rect 19809 7837 19843 7871
rect 3065 7769 3099 7803
rect 3281 7769 3315 7803
rect 4261 7769 4295 7803
rect 4353 7769 4387 7803
rect 4629 7769 4663 7803
rect 6193 7769 6227 7803
rect 9505 7769 9539 7803
rect 12265 7769 12299 7803
rect 14289 7769 14323 7803
rect 14657 7769 14691 7803
rect 15025 7769 15059 7803
rect 15853 7769 15887 7803
rect 17601 7769 17635 7803
rect 18245 7769 18279 7803
rect 18337 7769 18371 7803
rect 5089 7701 5123 7735
rect 6561 7701 6595 7735
rect 7389 7701 7423 7735
rect 10149 7701 10183 7735
rect 10701 7701 10735 7735
rect 15485 7701 15519 7735
rect 15653 7701 15687 7735
rect 16313 7701 16347 7735
rect 19441 7701 19475 7735
rect 4445 7497 4479 7531
rect 6561 7497 6595 7531
rect 7389 7497 7423 7531
rect 9413 7497 9447 7531
rect 10149 7497 10183 7531
rect 17601 7497 17635 7531
rect 18429 7497 18463 7531
rect 4261 7429 4295 7463
rect 10333 7429 10367 7463
rect 11713 7429 11747 7463
rect 12081 7429 12115 7463
rect 16005 7429 16039 7463
rect 16221 7429 16255 7463
rect 3893 7361 3927 7395
rect 6745 7361 6779 7395
rect 7665 7361 7699 7395
rect 8125 7361 8159 7395
rect 8953 7361 8987 7395
rect 9413 7361 9447 7395
rect 11897 7361 11931 7395
rect 12173 7361 12207 7395
rect 14289 7361 14323 7395
rect 17233 7361 17267 7395
rect 17325 7361 17359 7395
rect 17417 7361 17451 7395
rect 18613 7361 18647 7395
rect 18705 7361 18739 7395
rect 18797 7361 18831 7395
rect 6929 7293 6963 7327
rect 7389 7293 7423 7327
rect 7573 7293 7607 7327
rect 14013 7293 14047 7327
rect 8217 7225 8251 7259
rect 10701 7225 10735 7259
rect 15853 7225 15887 7259
rect 4261 7157 4295 7191
rect 9091 7157 9125 7191
rect 9229 7157 9263 7191
rect 10333 7157 10367 7191
rect 13737 7157 13771 7191
rect 14197 7157 14231 7191
rect 16037 7157 16071 7191
rect 15853 6953 15887 6987
rect 16037 6749 16071 6783
rect 16221 6749 16255 6783
rect 2237 2397 2271 2431
rect 5181 2397 5215 2431
rect 8125 2397 8159 2431
rect 10609 2397 10643 2431
rect 14289 2397 14323 2431
rect 16865 2397 16899 2431
rect 19441 2397 19475 2431
rect 21005 2397 21039 2431
rect 1961 2329 1995 2363
rect 4905 2329 4939 2363
rect 7849 2329 7883 2363
rect 10885 2329 10919 2363
rect 14565 2329 14599 2363
rect 17141 2329 17175 2363
rect 19717 2329 19751 2363
rect 21281 2329 21315 2363
<< metal1 >>
rect 1104 21786 22976 21808
rect 1104 21734 6378 21786
rect 6430 21734 6442 21786
rect 6494 21734 6506 21786
rect 6558 21734 6570 21786
rect 6622 21734 6634 21786
rect 6686 21734 11806 21786
rect 11858 21734 11870 21786
rect 11922 21734 11934 21786
rect 11986 21734 11998 21786
rect 12050 21734 12062 21786
rect 12114 21734 17234 21786
rect 17286 21734 17298 21786
rect 17350 21734 17362 21786
rect 17414 21734 17426 21786
rect 17478 21734 17490 21786
rect 17542 21734 22662 21786
rect 22714 21734 22726 21786
rect 22778 21734 22790 21786
rect 22842 21734 22854 21786
rect 22906 21734 22918 21786
rect 22970 21734 22976 21786
rect 1104 21712 22976 21734
rect 12158 21564 12164 21616
rect 12216 21564 12222 21616
rect 15289 21607 15347 21613
rect 15289 21604 15301 21607
rect 12406 21576 15301 21604
rect 12406 21468 12434 21576
rect 15289 21573 15301 21576
rect 15335 21604 15347 21607
rect 16482 21604 16488 21616
rect 15335 21576 16488 21604
rect 15335 21573 15347 21576
rect 15289 21567 15347 21573
rect 16482 21564 16488 21576
rect 16540 21564 16546 21616
rect 19978 21564 19984 21616
rect 20036 21604 20042 21616
rect 20441 21607 20499 21613
rect 20441 21604 20453 21607
rect 20036 21576 20453 21604
rect 20036 21564 20042 21576
rect 20441 21573 20453 21576
rect 20487 21573 20499 21607
rect 20441 21567 20499 21573
rect 15197 21539 15255 21545
rect 15197 21505 15209 21539
rect 15243 21505 15255 21539
rect 15197 21499 15255 21505
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21536 15531 21539
rect 16390 21536 16396 21548
rect 15519 21508 16396 21536
rect 15519 21505 15531 21508
rect 15473 21499 15531 21505
rect 10244 21440 12434 21468
rect 15212 21468 15240 21499
rect 16390 21496 16396 21508
rect 16448 21496 16454 21548
rect 19613 21539 19671 21545
rect 19613 21505 19625 21539
rect 19659 21505 19671 21539
rect 19613 21499 19671 21505
rect 16114 21468 16120 21480
rect 15212 21440 16120 21468
rect 10244 21344 10272 21440
rect 16114 21428 16120 21440
rect 16172 21428 16178 21480
rect 12345 21403 12403 21409
rect 12345 21369 12357 21403
rect 12391 21400 12403 21403
rect 15378 21400 15384 21412
rect 12391 21372 15384 21400
rect 12391 21369 12403 21372
rect 12345 21363 12403 21369
rect 15378 21360 15384 21372
rect 15436 21360 15442 21412
rect 17126 21360 17132 21412
rect 17184 21400 17190 21412
rect 19628 21400 19656 21499
rect 19702 21428 19708 21480
rect 19760 21468 19766 21480
rect 19797 21471 19855 21477
rect 19797 21468 19809 21471
rect 19760 21440 19809 21468
rect 19760 21428 19766 21440
rect 19797 21437 19809 21440
rect 19843 21437 19855 21471
rect 19797 21431 19855 21437
rect 17184 21372 19840 21400
rect 17184 21360 17190 21372
rect 19812 21344 19840 21372
rect 1854 21292 1860 21344
rect 1912 21332 1918 21344
rect 10226 21332 10232 21344
rect 1912 21304 10232 21332
rect 1912 21292 1918 21304
rect 10226 21292 10232 21304
rect 10284 21292 10290 21344
rect 15473 21335 15531 21341
rect 15473 21301 15485 21335
rect 15519 21332 15531 21335
rect 15930 21332 15936 21344
rect 15519 21304 15936 21332
rect 15519 21301 15531 21304
rect 15473 21295 15531 21301
rect 15930 21292 15936 21304
rect 15988 21292 15994 21344
rect 19426 21292 19432 21344
rect 19484 21292 19490 21344
rect 19794 21292 19800 21344
rect 19852 21292 19858 21344
rect 20346 21292 20352 21344
rect 20404 21292 20410 21344
rect 1104 21242 22816 21264
rect 1104 21190 3664 21242
rect 3716 21190 3728 21242
rect 3780 21190 3792 21242
rect 3844 21190 3856 21242
rect 3908 21190 3920 21242
rect 3972 21190 9092 21242
rect 9144 21190 9156 21242
rect 9208 21190 9220 21242
rect 9272 21190 9284 21242
rect 9336 21190 9348 21242
rect 9400 21190 14520 21242
rect 14572 21190 14584 21242
rect 14636 21190 14648 21242
rect 14700 21190 14712 21242
rect 14764 21190 14776 21242
rect 14828 21190 19948 21242
rect 20000 21190 20012 21242
rect 20064 21190 20076 21242
rect 20128 21190 20140 21242
rect 20192 21190 20204 21242
rect 20256 21190 22816 21242
rect 1104 21168 22816 21190
rect 2777 21131 2835 21137
rect 2777 21097 2789 21131
rect 2823 21128 2835 21131
rect 16117 21131 16175 21137
rect 16117 21128 16129 21131
rect 2823 21100 4568 21128
rect 2823 21097 2835 21100
rect 2777 21091 2835 21097
rect 4341 21063 4399 21069
rect 4341 21060 4353 21063
rect 2746 21032 4353 21060
rect 2746 20992 2774 21032
rect 4341 21029 4353 21032
rect 4387 21029 4399 21063
rect 4341 21023 4399 21029
rect 2148 20964 2774 20992
rect 2148 20933 2176 20964
rect 2958 20952 2964 21004
rect 3016 20992 3022 21004
rect 3016 20964 4476 20992
rect 3016 20952 3022 20964
rect 2041 20927 2099 20933
rect 2041 20893 2053 20927
rect 2087 20893 2099 20927
rect 2041 20887 2099 20893
rect 2133 20927 2191 20933
rect 2133 20893 2145 20927
rect 2179 20893 2191 20927
rect 2133 20887 2191 20893
rect 2056 20856 2084 20887
rect 2682 20856 2688 20868
rect 2056 20828 2688 20856
rect 2682 20816 2688 20828
rect 2740 20816 2746 20868
rect 2958 20816 2964 20868
rect 3016 20816 3022 20868
rect 3145 20859 3203 20865
rect 3145 20825 3157 20859
rect 3191 20856 3203 20859
rect 4246 20856 4252 20868
rect 3191 20828 4252 20856
rect 3191 20825 3203 20828
rect 3145 20819 3203 20825
rect 4246 20816 4252 20828
rect 4304 20816 4310 20868
rect 4448 20856 4476 20964
rect 4540 20924 4568 21100
rect 9048 21100 16129 21128
rect 5454 20927 5512 20933
rect 5454 20924 5466 20927
rect 4540 20896 5466 20924
rect 5454 20893 5466 20896
rect 5500 20893 5512 20927
rect 5454 20887 5512 20893
rect 5721 20927 5779 20933
rect 5721 20893 5733 20927
rect 5767 20924 5779 20927
rect 5994 20924 6000 20936
rect 5767 20896 6000 20924
rect 5767 20893 5779 20896
rect 5721 20887 5779 20893
rect 5994 20884 6000 20896
rect 6052 20884 6058 20936
rect 7006 20884 7012 20936
rect 7064 20924 7070 20936
rect 8573 20927 8631 20933
rect 8573 20924 8585 20927
rect 7064 20896 8585 20924
rect 7064 20884 7070 20896
rect 8573 20893 8585 20896
rect 8619 20893 8631 20927
rect 8573 20887 8631 20893
rect 8328 20859 8386 20865
rect 4448 20828 7328 20856
rect 2317 20791 2375 20797
rect 2317 20757 2329 20791
rect 2363 20788 2375 20791
rect 3970 20788 3976 20800
rect 2363 20760 3976 20788
rect 2363 20757 2375 20760
rect 2317 20751 2375 20757
rect 3970 20748 3976 20760
rect 4028 20748 4034 20800
rect 6914 20748 6920 20800
rect 6972 20788 6978 20800
rect 7193 20791 7251 20797
rect 7193 20788 7205 20791
rect 6972 20760 7205 20788
rect 6972 20748 6978 20760
rect 7193 20757 7205 20760
rect 7239 20757 7251 20791
rect 7300 20788 7328 20828
rect 8328 20825 8340 20859
rect 8374 20856 8386 20859
rect 9048 20856 9076 21100
rect 16117 21097 16129 21100
rect 16163 21097 16175 21131
rect 16117 21091 16175 21097
rect 16390 21088 16396 21140
rect 16448 21128 16454 21140
rect 17218 21128 17224 21140
rect 16448 21100 17224 21128
rect 16448 21088 16454 21100
rect 17218 21088 17224 21100
rect 17276 21088 17282 21140
rect 10226 21020 10232 21072
rect 10284 21020 10290 21072
rect 13633 21063 13691 21069
rect 13633 21029 13645 21063
rect 13679 21029 13691 21063
rect 13633 21023 13691 21029
rect 11517 20995 11575 21001
rect 11517 20961 11529 20995
rect 11563 20992 11575 20995
rect 13648 20992 13676 21023
rect 13814 21020 13820 21072
rect 13872 21060 13878 21072
rect 16485 21063 16543 21069
rect 16485 21060 16497 21063
rect 13872 21032 16497 21060
rect 13872 21020 13878 21032
rect 16485 21029 16497 21032
rect 16531 21060 16543 21063
rect 16531 21032 17080 21060
rect 16531 21029 16543 21032
rect 16485 21023 16543 21029
rect 11563 20964 12388 20992
rect 13648 20964 15700 20992
rect 11563 20961 11575 20964
rect 11517 20955 11575 20961
rect 11793 20927 11851 20933
rect 11793 20893 11805 20927
rect 11839 20924 11851 20927
rect 12158 20924 12164 20936
rect 11839 20896 12164 20924
rect 11839 20893 11851 20896
rect 11793 20887 11851 20893
rect 12158 20884 12164 20896
rect 12216 20924 12222 20936
rect 12253 20927 12311 20933
rect 12253 20924 12265 20927
rect 12216 20896 12265 20924
rect 12216 20884 12222 20896
rect 12253 20893 12265 20896
rect 12299 20893 12311 20927
rect 12360 20924 12388 20964
rect 15289 20927 15347 20933
rect 15289 20924 15301 20927
rect 12360 20896 15301 20924
rect 12253 20887 12311 20893
rect 15289 20893 15301 20896
rect 15335 20893 15347 20927
rect 15289 20887 15347 20893
rect 15470 20884 15476 20936
rect 15528 20884 15534 20936
rect 15672 20933 15700 20964
rect 15657 20927 15715 20933
rect 15657 20893 15669 20927
rect 15703 20924 15715 20927
rect 15703 20896 16252 20924
rect 15703 20893 15715 20896
rect 15657 20887 15715 20893
rect 8374 20828 9076 20856
rect 8374 20825 8386 20828
rect 8328 20819 8386 20825
rect 9122 20816 9128 20868
rect 9180 20816 9186 20868
rect 9306 20816 9312 20868
rect 9364 20816 9370 20868
rect 12520 20859 12578 20865
rect 12520 20825 12532 20859
rect 12566 20856 12578 20859
rect 16022 20856 16028 20868
rect 12566 20828 16028 20856
rect 12566 20825 12578 20828
rect 12520 20819 12578 20825
rect 16022 20816 16028 20828
rect 16080 20816 16086 20868
rect 16224 20856 16252 20896
rect 16298 20884 16304 20936
rect 16356 20884 16362 20936
rect 16482 20884 16488 20936
rect 16540 20924 16546 20936
rect 17052 20933 17080 21032
rect 17310 21020 17316 21072
rect 17368 21020 17374 21072
rect 17954 20952 17960 21004
rect 18012 20952 18018 21004
rect 16577 20927 16635 20933
rect 16577 20924 16589 20927
rect 16540 20896 16589 20924
rect 16540 20884 16546 20896
rect 16577 20893 16589 20896
rect 16623 20893 16635 20927
rect 16577 20887 16635 20893
rect 17037 20927 17095 20933
rect 17037 20893 17049 20927
rect 17083 20893 17095 20927
rect 17037 20887 17095 20893
rect 17144 20896 17448 20924
rect 17144 20856 17172 20896
rect 16224 20828 17172 20856
rect 17218 20816 17224 20868
rect 17276 20856 17282 20868
rect 17313 20859 17371 20865
rect 17313 20856 17325 20859
rect 17276 20828 17325 20856
rect 17276 20816 17282 20828
rect 17313 20825 17325 20828
rect 17359 20825 17371 20859
rect 17420 20856 17448 20896
rect 18230 20884 18236 20936
rect 18288 20884 18294 20936
rect 19702 20884 19708 20936
rect 19760 20884 19766 20936
rect 19886 20884 19892 20936
rect 19944 20924 19950 20936
rect 20073 20927 20131 20933
rect 20073 20924 20085 20927
rect 19944 20896 20085 20924
rect 19944 20884 19950 20896
rect 20073 20893 20085 20896
rect 20119 20893 20131 20927
rect 20073 20887 20131 20893
rect 19720 20856 19748 20884
rect 17420 20828 19748 20856
rect 20444 20868 20496 20874
rect 17313 20819 17371 20825
rect 9324 20788 9352 20816
rect 20444 20810 20496 20816
rect 7300 20760 9352 20788
rect 9493 20791 9551 20797
rect 7193 20751 7251 20757
rect 9493 20757 9505 20791
rect 9539 20788 9551 20791
rect 9950 20788 9956 20800
rect 9539 20760 9956 20788
rect 9539 20757 9551 20760
rect 9493 20751 9551 20757
rect 9950 20748 9956 20760
rect 10008 20748 10014 20800
rect 16482 20748 16488 20800
rect 16540 20788 16546 20800
rect 17129 20791 17187 20797
rect 17129 20788 17141 20791
rect 16540 20760 17141 20788
rect 16540 20748 16546 20760
rect 17129 20757 17141 20760
rect 17175 20788 17187 20791
rect 18690 20788 18696 20800
rect 17175 20760 18696 20788
rect 17175 20757 17187 20760
rect 17129 20751 17187 20757
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 18782 20748 18788 20800
rect 18840 20788 18846 20800
rect 18877 20791 18935 20797
rect 18877 20788 18889 20791
rect 18840 20760 18889 20788
rect 18840 20748 18846 20760
rect 18877 20757 18889 20760
rect 18923 20757 18935 20791
rect 18877 20751 18935 20757
rect 1104 20698 22976 20720
rect 1104 20646 6378 20698
rect 6430 20646 6442 20698
rect 6494 20646 6506 20698
rect 6558 20646 6570 20698
rect 6622 20646 6634 20698
rect 6686 20646 11806 20698
rect 11858 20646 11870 20698
rect 11922 20646 11934 20698
rect 11986 20646 11998 20698
rect 12050 20646 12062 20698
rect 12114 20646 17234 20698
rect 17286 20646 17298 20698
rect 17350 20646 17362 20698
rect 17414 20646 17426 20698
rect 17478 20646 17490 20698
rect 17542 20646 22662 20698
rect 22714 20646 22726 20698
rect 22778 20646 22790 20698
rect 22842 20646 22854 20698
rect 22906 20646 22918 20698
rect 22970 20646 22976 20698
rect 1104 20624 22976 20646
rect 1854 20544 1860 20596
rect 1912 20544 1918 20596
rect 2958 20584 2964 20596
rect 2056 20556 2964 20584
rect 2056 20525 2084 20556
rect 2958 20544 2964 20556
rect 3016 20544 3022 20596
rect 4246 20544 4252 20596
rect 4304 20584 4310 20596
rect 4341 20587 4399 20593
rect 4341 20584 4353 20587
rect 4304 20556 4353 20584
rect 4304 20544 4310 20556
rect 4341 20553 4353 20556
rect 4387 20553 4399 20587
rect 4341 20547 4399 20553
rect 8389 20587 8447 20593
rect 8389 20553 8401 20587
rect 8435 20584 8447 20587
rect 9122 20584 9128 20596
rect 8435 20556 9128 20584
rect 8435 20553 8447 20556
rect 8389 20547 8447 20553
rect 9122 20544 9128 20556
rect 9180 20544 9186 20596
rect 13814 20544 13820 20596
rect 13872 20544 13878 20596
rect 17954 20544 17960 20596
rect 18012 20584 18018 20596
rect 18049 20587 18107 20593
rect 18049 20584 18061 20587
rect 18012 20556 18061 20584
rect 18012 20544 18018 20556
rect 18049 20553 18061 20556
rect 18095 20553 18107 20587
rect 18049 20547 18107 20553
rect 18230 20544 18236 20596
rect 18288 20584 18294 20596
rect 18693 20587 18751 20593
rect 18693 20584 18705 20587
rect 18288 20556 18705 20584
rect 18288 20544 18294 20556
rect 18693 20553 18705 20556
rect 18739 20553 18751 20587
rect 18693 20547 18751 20553
rect 2041 20519 2099 20525
rect 2041 20485 2053 20519
rect 2087 20485 2099 20519
rect 6914 20516 6920 20528
rect 2041 20479 2099 20485
rect 2700 20488 6920 20516
rect 1762 20408 1768 20460
rect 1820 20408 1826 20460
rect 2700 20457 2728 20488
rect 6914 20476 6920 20488
rect 6972 20476 6978 20528
rect 9950 20525 9956 20528
rect 9944 20516 9956 20525
rect 9911 20488 9956 20516
rect 9944 20479 9956 20488
rect 9950 20476 9956 20479
rect 10008 20476 10014 20528
rect 12704 20519 12762 20525
rect 12704 20485 12716 20519
rect 12750 20516 12762 20519
rect 15749 20519 15807 20525
rect 15749 20516 15761 20519
rect 12750 20488 15761 20516
rect 12750 20485 12762 20488
rect 12704 20479 12762 20485
rect 15749 20485 15761 20488
rect 15795 20485 15807 20519
rect 20438 20516 20444 20528
rect 15749 20479 15807 20485
rect 18892 20488 20444 20516
rect 2685 20451 2743 20457
rect 2685 20417 2697 20451
rect 2731 20417 2743 20451
rect 2685 20411 2743 20417
rect 3050 20408 3056 20460
rect 3108 20448 3114 20460
rect 5454 20451 5512 20457
rect 5454 20448 5466 20451
rect 3108 20420 5466 20448
rect 3108 20408 3114 20420
rect 5454 20417 5466 20420
rect 5500 20417 5512 20451
rect 5454 20411 5512 20417
rect 7006 20408 7012 20460
rect 7064 20408 7070 20460
rect 7265 20451 7323 20457
rect 7265 20448 7277 20451
rect 7116 20420 7277 20448
rect 2501 20383 2559 20389
rect 2501 20349 2513 20383
rect 2547 20380 2559 20383
rect 5721 20383 5779 20389
rect 2547 20352 2728 20380
rect 2547 20349 2559 20352
rect 2501 20343 2559 20349
rect 2700 20324 2728 20352
rect 5721 20349 5733 20383
rect 5767 20380 5779 20383
rect 5994 20380 6000 20392
rect 5767 20352 6000 20380
rect 5767 20349 5779 20352
rect 5721 20343 5779 20349
rect 5994 20340 6000 20352
rect 6052 20340 6058 20392
rect 7116 20380 7144 20420
rect 7265 20417 7277 20420
rect 7311 20417 7323 20451
rect 7265 20411 7323 20417
rect 9306 20408 9312 20460
rect 9364 20448 9370 20460
rect 14366 20448 14372 20460
rect 9364 20420 14372 20448
rect 9364 20408 9370 20420
rect 14366 20408 14372 20420
rect 14424 20448 14430 20460
rect 14461 20451 14519 20457
rect 14461 20448 14473 20451
rect 14424 20420 14473 20448
rect 14424 20408 14430 20420
rect 14461 20417 14473 20420
rect 14507 20417 14519 20451
rect 14461 20411 14519 20417
rect 15289 20451 15347 20457
rect 15289 20417 15301 20451
rect 15335 20448 15347 20451
rect 15378 20448 15384 20460
rect 15335 20420 15384 20448
rect 15335 20417 15347 20420
rect 15289 20411 15347 20417
rect 15378 20408 15384 20420
rect 15436 20408 15442 20460
rect 15930 20408 15936 20460
rect 15988 20408 15994 20460
rect 16209 20451 16267 20457
rect 16209 20417 16221 20451
rect 16255 20448 16267 20451
rect 16482 20448 16488 20460
rect 16255 20420 16488 20448
rect 16255 20417 16267 20420
rect 16209 20411 16267 20417
rect 16482 20408 16488 20420
rect 16540 20408 16546 20460
rect 17034 20408 17040 20460
rect 17092 20408 17098 20460
rect 17218 20408 17224 20460
rect 17276 20408 17282 20460
rect 18892 20457 18920 20488
rect 20438 20476 20444 20488
rect 20496 20476 20502 20528
rect 18877 20451 18935 20457
rect 18877 20417 18889 20451
rect 18923 20417 18935 20451
rect 18877 20411 18935 20417
rect 19153 20451 19211 20457
rect 19153 20417 19165 20451
rect 19199 20448 19211 20451
rect 19426 20448 19432 20460
rect 19199 20420 19432 20448
rect 19199 20417 19211 20420
rect 19153 20411 19211 20417
rect 19426 20408 19432 20420
rect 19484 20408 19490 20460
rect 6104 20352 7144 20380
rect 2682 20272 2688 20324
rect 2740 20272 2746 20324
rect 2041 20247 2099 20253
rect 2041 20213 2053 20247
rect 2087 20244 2099 20247
rect 2222 20244 2228 20256
rect 2087 20216 2228 20244
rect 2087 20213 2099 20216
rect 2041 20207 2099 20213
rect 2222 20204 2228 20216
rect 2280 20204 2286 20256
rect 2866 20204 2872 20256
rect 2924 20204 2930 20256
rect 3970 20204 3976 20256
rect 4028 20244 4034 20256
rect 6104 20244 6132 20352
rect 9490 20340 9496 20392
rect 9548 20380 9554 20392
rect 9677 20383 9735 20389
rect 9677 20380 9689 20383
rect 9548 20352 9689 20380
rect 9548 20340 9554 20352
rect 9677 20349 9689 20352
rect 9723 20349 9735 20383
rect 9677 20343 9735 20349
rect 12158 20340 12164 20392
rect 12216 20380 12222 20392
rect 12437 20383 12495 20389
rect 12437 20380 12449 20383
rect 12216 20352 12449 20380
rect 12216 20340 12222 20352
rect 12437 20349 12449 20352
rect 12483 20349 12495 20383
rect 12437 20343 12495 20349
rect 18966 20340 18972 20392
rect 19024 20340 19030 20392
rect 19061 20383 19119 20389
rect 19061 20349 19073 20383
rect 19107 20349 19119 20383
rect 19061 20343 19119 20349
rect 15194 20312 15200 20324
rect 13740 20284 15200 20312
rect 4028 20216 6132 20244
rect 11057 20247 11115 20253
rect 4028 20204 4034 20216
rect 11057 20213 11069 20247
rect 11103 20244 11115 20247
rect 13740 20244 13768 20284
rect 15194 20272 15200 20284
rect 15252 20272 15258 20324
rect 18690 20272 18696 20324
rect 18748 20312 18754 20324
rect 19076 20312 19104 20343
rect 18748 20284 19104 20312
rect 18748 20272 18754 20284
rect 11103 20216 13768 20244
rect 11103 20213 11115 20216
rect 11057 20207 11115 20213
rect 16114 20204 16120 20256
rect 16172 20204 16178 20256
rect 1104 20154 22816 20176
rect 1104 20102 3664 20154
rect 3716 20102 3728 20154
rect 3780 20102 3792 20154
rect 3844 20102 3856 20154
rect 3908 20102 3920 20154
rect 3972 20102 9092 20154
rect 9144 20102 9156 20154
rect 9208 20102 9220 20154
rect 9272 20102 9284 20154
rect 9336 20102 9348 20154
rect 9400 20102 14520 20154
rect 14572 20102 14584 20154
rect 14636 20102 14648 20154
rect 14700 20102 14712 20154
rect 14764 20102 14776 20154
rect 14828 20102 19948 20154
rect 20000 20102 20012 20154
rect 20064 20102 20076 20154
rect 20128 20102 20140 20154
rect 20192 20102 20204 20154
rect 20256 20102 22816 20154
rect 1104 20080 22816 20102
rect 3050 20000 3056 20052
rect 3108 20000 3114 20052
rect 16022 20000 16028 20052
rect 16080 20000 16086 20052
rect 1762 19932 1768 19984
rect 1820 19972 1826 19984
rect 2041 19975 2099 19981
rect 2041 19972 2053 19975
rect 1820 19944 2053 19972
rect 1820 19932 1826 19944
rect 2041 19941 2053 19944
rect 2087 19972 2099 19975
rect 4433 19975 4491 19981
rect 4433 19972 4445 19975
rect 2087 19944 4445 19972
rect 2087 19941 2099 19944
rect 2041 19935 2099 19941
rect 4433 19941 4445 19944
rect 4479 19941 4491 19975
rect 4433 19935 4491 19941
rect 13541 19975 13599 19981
rect 13541 19941 13553 19975
rect 13587 19972 13599 19975
rect 17034 19972 17040 19984
rect 13587 19944 17040 19972
rect 13587 19941 13599 19944
rect 13541 19935 13599 19941
rect 17034 19932 17040 19944
rect 17092 19932 17098 19984
rect 1854 19864 1860 19916
rect 1912 19904 1918 19916
rect 1949 19907 2007 19913
rect 1949 19904 1961 19907
rect 1912 19876 1961 19904
rect 1912 19864 1918 19876
rect 1949 19873 1961 19876
rect 1995 19873 2007 19907
rect 1949 19867 2007 19873
rect 14645 19907 14703 19913
rect 14645 19873 14657 19907
rect 14691 19904 14703 19907
rect 16390 19904 16396 19916
rect 14691 19876 15700 19904
rect 14691 19873 14703 19876
rect 14645 19867 14703 19873
rect 2222 19796 2228 19848
rect 2280 19796 2286 19848
rect 2866 19796 2872 19848
rect 2924 19836 2930 19848
rect 5546 19839 5604 19845
rect 5546 19836 5558 19839
rect 2924 19808 5558 19836
rect 2924 19796 2930 19808
rect 5546 19805 5558 19808
rect 5592 19805 5604 19839
rect 5546 19799 5604 19805
rect 5813 19839 5871 19845
rect 5813 19805 5825 19839
rect 5859 19836 5871 19839
rect 5994 19836 6000 19848
rect 5859 19808 6000 19836
rect 5859 19805 5871 19808
rect 5813 19799 5871 19805
rect 5994 19796 6000 19808
rect 6052 19796 6058 19848
rect 11698 19796 11704 19848
rect 11756 19836 11762 19848
rect 12158 19836 12164 19848
rect 11756 19808 12164 19836
rect 11756 19796 11762 19808
rect 12158 19796 12164 19808
rect 12216 19796 12222 19848
rect 13354 19796 13360 19848
rect 13412 19836 13418 19848
rect 15565 19839 15623 19845
rect 15565 19836 15577 19839
rect 13412 19808 15577 19836
rect 13412 19796 13418 19808
rect 15565 19805 15577 19808
rect 15611 19805 15623 19839
rect 15565 19799 15623 19805
rect 2498 19728 2504 19780
rect 2556 19768 2562 19780
rect 2958 19768 2964 19780
rect 2556 19740 2964 19768
rect 2556 19728 2562 19740
rect 2958 19728 2964 19740
rect 3016 19768 3022 19780
rect 3237 19771 3295 19777
rect 3237 19768 3249 19771
rect 3016 19740 3249 19768
rect 3016 19728 3022 19740
rect 3237 19737 3249 19740
rect 3283 19737 3295 19771
rect 3237 19731 3295 19737
rect 3421 19771 3479 19777
rect 3421 19737 3433 19771
rect 3467 19768 3479 19771
rect 4522 19768 4528 19780
rect 3467 19740 4528 19768
rect 3467 19737 3479 19740
rect 3421 19731 3479 19737
rect 4522 19728 4528 19740
rect 4580 19728 4586 19780
rect 12428 19771 12486 19777
rect 12428 19737 12440 19771
rect 12474 19768 12486 19771
rect 14274 19768 14280 19780
rect 12474 19740 14280 19768
rect 12474 19737 12486 19740
rect 12428 19731 12486 19737
rect 14274 19728 14280 19740
rect 14332 19728 14338 19780
rect 14366 19728 14372 19780
rect 14424 19728 14430 19780
rect 15194 19728 15200 19780
rect 15252 19728 15258 19780
rect 15381 19771 15439 19777
rect 15381 19737 15393 19771
rect 15427 19768 15439 19771
rect 15672 19768 15700 19876
rect 16132 19876 16396 19904
rect 16132 19768 16160 19876
rect 16390 19864 16396 19876
rect 16448 19864 16454 19916
rect 17218 19836 17224 19848
rect 16224 19808 17224 19836
rect 16224 19777 16252 19808
rect 17218 19796 17224 19808
rect 17276 19796 17282 19848
rect 15427 19740 16160 19768
rect 16209 19771 16267 19777
rect 15427 19737 15439 19740
rect 15381 19731 15439 19737
rect 16209 19737 16221 19771
rect 16255 19737 16267 19771
rect 16209 19731 16267 19737
rect 2406 19660 2412 19712
rect 2464 19660 2470 19712
rect 4062 19660 4068 19712
rect 4120 19700 4126 19712
rect 8294 19700 8300 19712
rect 4120 19672 8300 19700
rect 4120 19660 4126 19672
rect 8294 19660 8300 19672
rect 8352 19660 8358 19712
rect 15102 19660 15108 19712
rect 15160 19700 15166 19712
rect 16224 19700 16252 19731
rect 16390 19728 16396 19780
rect 16448 19728 16454 19780
rect 15160 19672 16252 19700
rect 15160 19660 15166 19672
rect 1104 19610 22976 19632
rect 1104 19558 6378 19610
rect 6430 19558 6442 19610
rect 6494 19558 6506 19610
rect 6558 19558 6570 19610
rect 6622 19558 6634 19610
rect 6686 19558 11806 19610
rect 11858 19558 11870 19610
rect 11922 19558 11934 19610
rect 11986 19558 11998 19610
rect 12050 19558 12062 19610
rect 12114 19558 17234 19610
rect 17286 19558 17298 19610
rect 17350 19558 17362 19610
rect 17414 19558 17426 19610
rect 17478 19558 17490 19610
rect 17542 19558 22662 19610
rect 22714 19558 22726 19610
rect 22778 19558 22790 19610
rect 22842 19558 22854 19610
rect 22906 19558 22918 19610
rect 22970 19558 22976 19610
rect 1104 19536 22976 19558
rect 2501 19499 2559 19505
rect 2501 19465 2513 19499
rect 2547 19496 2559 19499
rect 10873 19499 10931 19505
rect 2547 19468 7144 19496
rect 2547 19465 2559 19468
rect 2501 19459 2559 19465
rect 2406 19388 2412 19440
rect 2464 19428 2470 19440
rect 2464 19400 4016 19428
rect 2464 19388 2470 19400
rect 1854 19320 1860 19372
rect 1912 19360 1918 19372
rect 2133 19363 2191 19369
rect 2133 19360 2145 19363
rect 1912 19332 2145 19360
rect 1912 19320 1918 19332
rect 2133 19329 2145 19332
rect 2179 19329 2191 19363
rect 2133 19323 2191 19329
rect 2317 19363 2375 19369
rect 2317 19329 2329 19363
rect 2363 19360 2375 19363
rect 2682 19360 2688 19372
rect 2363 19332 2688 19360
rect 2363 19329 2375 19332
rect 2317 19323 2375 19329
rect 2682 19320 2688 19332
rect 2740 19320 2746 19372
rect 3988 19360 4016 19400
rect 5730 19363 5788 19369
rect 5730 19360 5742 19363
rect 3988 19332 5742 19360
rect 5730 19329 5742 19332
rect 5776 19329 5788 19363
rect 5730 19323 5788 19329
rect 5994 19320 6000 19372
rect 6052 19360 6058 19372
rect 6917 19363 6975 19369
rect 6917 19360 6929 19363
rect 6052 19332 6929 19360
rect 6052 19320 6058 19332
rect 6917 19329 6929 19332
rect 6963 19360 6975 19363
rect 7006 19360 7012 19372
rect 6963 19332 7012 19360
rect 6963 19329 6975 19332
rect 6917 19323 6975 19329
rect 7006 19320 7012 19332
rect 7064 19320 7070 19372
rect 7116 19360 7144 19468
rect 10873 19465 10885 19499
rect 10919 19496 10931 19499
rect 16114 19496 16120 19508
rect 10919 19468 16120 19496
rect 10919 19465 10931 19468
rect 10873 19459 10931 19465
rect 16114 19456 16120 19468
rect 16172 19456 16178 19508
rect 16853 19499 16911 19505
rect 16853 19465 16865 19499
rect 16899 19465 16911 19499
rect 16853 19459 16911 19465
rect 12336 19431 12394 19437
rect 12336 19397 12348 19431
rect 12382 19428 12394 19431
rect 13354 19428 13360 19440
rect 12382 19400 13360 19428
rect 12382 19397 12394 19400
rect 12336 19391 12394 19397
rect 13354 19388 13360 19400
rect 13412 19388 13418 19440
rect 13538 19388 13544 19440
rect 13596 19428 13602 19440
rect 14645 19431 14703 19437
rect 14645 19428 14657 19431
rect 13596 19400 14657 19428
rect 13596 19388 13602 19400
rect 14645 19397 14657 19400
rect 14691 19397 14703 19431
rect 16868 19428 16896 19459
rect 14645 19391 14703 19397
rect 16132 19400 16896 19428
rect 9766 19369 9772 19372
rect 7173 19363 7231 19369
rect 7173 19360 7185 19363
rect 7116 19332 7185 19360
rect 7173 19329 7185 19332
rect 7219 19329 7231 19363
rect 7173 19323 7231 19329
rect 9760 19323 9772 19369
rect 9766 19320 9772 19323
rect 9824 19320 9830 19372
rect 16132 19369 16160 19400
rect 17034 19388 17040 19440
rect 17092 19428 17098 19440
rect 17092 19400 17264 19428
rect 17092 19388 17098 19400
rect 14829 19363 14887 19369
rect 14829 19360 14841 19363
rect 13464 19332 14841 19360
rect 9490 19252 9496 19304
rect 9548 19252 9554 19304
rect 11698 19252 11704 19304
rect 11756 19292 11762 19304
rect 12069 19295 12127 19301
rect 12069 19292 12081 19295
rect 11756 19264 12081 19292
rect 11756 19252 11762 19264
rect 12069 19261 12081 19264
rect 12115 19261 12127 19295
rect 12069 19255 12127 19261
rect 13464 19233 13492 19332
rect 14829 19329 14841 19332
rect 14875 19329 14887 19363
rect 14829 19323 14887 19329
rect 16117 19363 16175 19369
rect 16117 19329 16129 19363
rect 16163 19329 16175 19363
rect 16117 19323 16175 19329
rect 16301 19363 16359 19369
rect 16301 19329 16313 19363
rect 16347 19360 16359 19363
rect 16574 19360 16580 19372
rect 16347 19332 16580 19360
rect 16347 19329 16359 19332
rect 16301 19323 16359 19329
rect 16574 19320 16580 19332
rect 16632 19320 16638 19372
rect 17236 19369 17264 19400
rect 18690 19388 18696 19440
rect 18748 19428 18754 19440
rect 18877 19431 18935 19437
rect 18877 19428 18889 19431
rect 18748 19400 18889 19428
rect 18748 19388 18754 19400
rect 18877 19397 18889 19400
rect 18923 19428 18935 19431
rect 18923 19400 19748 19428
rect 18923 19397 18935 19400
rect 18877 19391 18935 19397
rect 17221 19363 17279 19369
rect 17221 19329 17233 19363
rect 17267 19329 17279 19363
rect 17221 19323 17279 19329
rect 18598 19320 18604 19372
rect 18656 19360 18662 19372
rect 18966 19360 18972 19372
rect 18656 19332 18972 19360
rect 18656 19320 18662 19332
rect 18966 19320 18972 19332
rect 19024 19360 19030 19372
rect 19720 19369 19748 19400
rect 19061 19363 19119 19369
rect 19061 19360 19073 19363
rect 19024 19332 19073 19360
rect 19024 19320 19030 19332
rect 19061 19329 19073 19332
rect 19107 19360 19119 19363
rect 19521 19363 19579 19369
rect 19521 19360 19533 19363
rect 19107 19332 19533 19360
rect 19107 19329 19119 19332
rect 19061 19323 19119 19329
rect 19521 19329 19533 19332
rect 19567 19329 19579 19363
rect 19521 19323 19579 19329
rect 19705 19363 19763 19369
rect 19705 19329 19717 19363
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19292 15071 19295
rect 15470 19292 15476 19304
rect 15059 19264 15476 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 15470 19252 15476 19264
rect 15528 19292 15534 19304
rect 16022 19292 16028 19304
rect 15528 19264 16028 19292
rect 15528 19252 15534 19264
rect 16022 19252 16028 19264
rect 16080 19252 16086 19304
rect 16482 19252 16488 19304
rect 16540 19292 16546 19304
rect 17037 19295 17095 19301
rect 17037 19292 17049 19295
rect 16540 19264 17049 19292
rect 16540 19252 16546 19264
rect 17037 19261 17049 19264
rect 17083 19261 17095 19295
rect 17037 19255 17095 19261
rect 17126 19252 17132 19304
rect 17184 19252 17190 19304
rect 17313 19295 17371 19301
rect 17313 19261 17325 19295
rect 17359 19292 17371 19295
rect 19334 19292 19340 19304
rect 17359 19264 19340 19292
rect 17359 19261 17371 19264
rect 17313 19255 17371 19261
rect 13449 19227 13507 19233
rect 13449 19193 13461 19227
rect 13495 19193 13507 19227
rect 13449 19187 13507 19193
rect 14274 19184 14280 19236
rect 14332 19224 14338 19236
rect 16117 19227 16175 19233
rect 16117 19224 16129 19227
rect 14332 19196 16129 19224
rect 14332 19184 14338 19196
rect 16117 19193 16129 19196
rect 16163 19193 16175 19227
rect 16117 19187 16175 19193
rect 4614 19116 4620 19168
rect 4672 19116 4678 19168
rect 8297 19159 8355 19165
rect 8297 19125 8309 19159
rect 8343 19156 8355 19159
rect 8386 19156 8392 19168
rect 8343 19128 8392 19156
rect 8343 19125 8355 19128
rect 8297 19119 8355 19125
rect 8386 19116 8392 19128
rect 8444 19116 8450 19168
rect 16390 19116 16396 19168
rect 16448 19156 16454 19168
rect 17328 19156 17356 19255
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 16448 19128 17356 19156
rect 16448 19116 16454 19128
rect 18690 19116 18696 19168
rect 18748 19116 18754 19168
rect 19610 19116 19616 19168
rect 19668 19116 19674 19168
rect 1104 19066 22816 19088
rect 1104 19014 3664 19066
rect 3716 19014 3728 19066
rect 3780 19014 3792 19066
rect 3844 19014 3856 19066
rect 3908 19014 3920 19066
rect 3972 19014 9092 19066
rect 9144 19014 9156 19066
rect 9208 19014 9220 19066
rect 9272 19014 9284 19066
rect 9336 19014 9348 19066
rect 9400 19014 14520 19066
rect 14572 19014 14584 19066
rect 14636 19014 14648 19066
rect 14700 19014 14712 19066
rect 14764 19014 14776 19066
rect 14828 19014 19948 19066
rect 20000 19014 20012 19066
rect 20064 19014 20076 19066
rect 20128 19014 20140 19066
rect 20192 19014 20204 19066
rect 20256 19014 22816 19066
rect 1104 18992 22816 19014
rect 4522 18912 4528 18964
rect 4580 18912 4586 18964
rect 8389 18955 8447 18961
rect 8389 18921 8401 18955
rect 8435 18952 8447 18955
rect 9674 18952 9680 18964
rect 8435 18924 9680 18952
rect 8435 18921 8447 18924
rect 8389 18915 8447 18921
rect 9674 18912 9680 18924
rect 9732 18912 9738 18964
rect 10689 18955 10747 18961
rect 10689 18921 10701 18955
rect 10735 18952 10747 18955
rect 15102 18952 15108 18964
rect 10735 18924 15108 18952
rect 10735 18921 10747 18924
rect 10689 18915 10747 18921
rect 15102 18912 15108 18924
rect 15160 18912 15166 18964
rect 16574 18912 16580 18964
rect 16632 18912 16638 18964
rect 5905 18819 5963 18825
rect 5905 18785 5917 18819
rect 5951 18816 5963 18819
rect 5994 18816 6000 18828
rect 5951 18788 6000 18816
rect 5951 18785 5963 18788
rect 5905 18779 5963 18785
rect 5994 18776 6000 18788
rect 6052 18776 6058 18828
rect 13538 18816 13544 18828
rect 10980 18788 13544 18816
rect 2682 18708 2688 18760
rect 2740 18748 2746 18760
rect 3053 18751 3111 18757
rect 3053 18748 3065 18751
rect 2740 18720 3065 18748
rect 2740 18708 2746 18720
rect 3053 18717 3065 18720
rect 3099 18717 3111 18751
rect 3053 18711 3111 18717
rect 3237 18751 3295 18757
rect 3237 18717 3249 18751
rect 3283 18748 3295 18751
rect 4614 18748 4620 18760
rect 3283 18720 4620 18748
rect 3283 18717 3295 18720
rect 3237 18711 3295 18717
rect 4614 18708 4620 18720
rect 4672 18708 4678 18760
rect 8110 18708 8116 18760
rect 8168 18708 8174 18760
rect 8205 18751 8263 18757
rect 8205 18717 8217 18751
rect 8251 18748 8263 18751
rect 8386 18748 8392 18760
rect 8251 18720 8392 18748
rect 8251 18717 8263 18720
rect 8205 18711 8263 18717
rect 8386 18708 8392 18720
rect 8444 18708 8450 18760
rect 9309 18751 9367 18757
rect 9309 18717 9321 18751
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 9576 18751 9634 18757
rect 9576 18717 9588 18751
rect 9622 18748 9634 18751
rect 10980 18748 11008 18788
rect 13538 18776 13544 18788
rect 13596 18776 13602 18828
rect 20349 18819 20407 18825
rect 18708 18788 19472 18816
rect 18708 18760 18736 18788
rect 9622 18720 11008 18748
rect 9622 18717 9634 18720
rect 9576 18711 9634 18717
rect 4062 18640 4068 18692
rect 4120 18680 4126 18692
rect 5638 18683 5696 18689
rect 5638 18680 5650 18683
rect 4120 18652 5650 18680
rect 4120 18640 4126 18652
rect 5638 18649 5650 18652
rect 5684 18649 5696 18683
rect 9324 18680 9352 18711
rect 11698 18708 11704 18760
rect 11756 18748 11762 18760
rect 12069 18751 12127 18757
rect 12069 18748 12081 18751
rect 11756 18720 12081 18748
rect 11756 18708 11762 18720
rect 12069 18717 12081 18720
rect 12115 18717 12127 18751
rect 12069 18711 12127 18717
rect 12345 18751 12403 18757
rect 12345 18717 12357 18751
rect 12391 18748 12403 18751
rect 15286 18748 15292 18760
rect 12391 18720 15292 18748
rect 12391 18717 12403 18720
rect 12345 18711 12403 18717
rect 15286 18708 15292 18720
rect 15344 18708 15350 18760
rect 15654 18708 15660 18760
rect 15712 18748 15718 18760
rect 16482 18748 16488 18760
rect 15712 18720 16488 18748
rect 15712 18708 15718 18720
rect 16482 18708 16488 18720
rect 16540 18748 16546 18760
rect 16853 18751 16911 18757
rect 16853 18748 16865 18751
rect 16540 18720 16865 18748
rect 16540 18708 16546 18720
rect 16853 18717 16865 18720
rect 16899 18748 16911 18751
rect 18598 18748 18604 18760
rect 16899 18720 18604 18748
rect 16899 18717 16911 18720
rect 16853 18711 16911 18717
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 18690 18708 18696 18760
rect 18748 18708 18754 18760
rect 19444 18757 19472 18788
rect 20349 18785 20361 18819
rect 20395 18816 20407 18819
rect 20438 18816 20444 18828
rect 20395 18788 20444 18816
rect 20395 18785 20407 18788
rect 20349 18779 20407 18785
rect 20438 18776 20444 18788
rect 20496 18776 20502 18828
rect 18877 18751 18935 18757
rect 18877 18717 18889 18751
rect 18923 18717 18935 18751
rect 18877 18711 18935 18717
rect 19429 18751 19487 18757
rect 19429 18717 19441 18751
rect 19475 18717 19487 18751
rect 19429 18711 19487 18717
rect 16577 18683 16635 18689
rect 9324 18652 9628 18680
rect 5638 18643 5696 18649
rect 9600 18624 9628 18652
rect 16577 18649 16589 18683
rect 16623 18680 16635 18683
rect 17034 18680 17040 18692
rect 16623 18652 17040 18680
rect 16623 18649 16635 18652
rect 16577 18643 16635 18649
rect 17034 18640 17040 18652
rect 17092 18640 17098 18692
rect 18892 18680 18920 18711
rect 19610 18708 19616 18760
rect 19668 18708 19674 18760
rect 19628 18680 19656 18708
rect 20272 18680 20300 18734
rect 18892 18652 20300 18680
rect 20901 18683 20959 18689
rect 20901 18649 20913 18683
rect 20947 18680 20959 18683
rect 20990 18680 20996 18692
rect 20947 18652 20996 18680
rect 20947 18649 20959 18652
rect 20901 18643 20959 18649
rect 20990 18640 20996 18652
rect 21048 18640 21054 18692
rect 3418 18572 3424 18624
rect 3476 18572 3482 18624
rect 9582 18572 9588 18624
rect 9640 18572 9646 18624
rect 13633 18615 13691 18621
rect 13633 18581 13645 18615
rect 13679 18612 13691 18615
rect 15746 18612 15752 18624
rect 13679 18584 15752 18612
rect 13679 18581 13691 18584
rect 13633 18575 13691 18581
rect 15746 18572 15752 18584
rect 15804 18612 15810 18624
rect 16761 18615 16819 18621
rect 16761 18612 16773 18615
rect 15804 18584 16773 18612
rect 15804 18572 15810 18584
rect 16761 18581 16773 18584
rect 16807 18612 16819 18615
rect 17126 18612 17132 18624
rect 16807 18584 17132 18612
rect 16807 18581 16819 18584
rect 16761 18575 16819 18581
rect 17126 18572 17132 18584
rect 17184 18572 17190 18624
rect 18506 18572 18512 18624
rect 18564 18572 18570 18624
rect 19610 18572 19616 18624
rect 19668 18572 19674 18624
rect 1104 18522 22976 18544
rect 1104 18470 6378 18522
rect 6430 18470 6442 18522
rect 6494 18470 6506 18522
rect 6558 18470 6570 18522
rect 6622 18470 6634 18522
rect 6686 18470 11806 18522
rect 11858 18470 11870 18522
rect 11922 18470 11934 18522
rect 11986 18470 11998 18522
rect 12050 18470 12062 18522
rect 12114 18470 17234 18522
rect 17286 18470 17298 18522
rect 17350 18470 17362 18522
rect 17414 18470 17426 18522
rect 17478 18470 17490 18522
rect 17542 18470 22662 18522
rect 22714 18470 22726 18522
rect 22778 18470 22790 18522
rect 22842 18470 22854 18522
rect 22906 18470 22918 18522
rect 22970 18470 22976 18522
rect 1104 18448 22976 18470
rect 4062 18368 4068 18420
rect 4120 18368 4126 18420
rect 15286 18368 15292 18420
rect 15344 18368 15350 18420
rect 2682 18340 2688 18352
rect 1964 18312 2688 18340
rect 1964 18281 1992 18312
rect 2682 18300 2688 18312
rect 2740 18340 2746 18352
rect 2740 18300 2774 18340
rect 3418 18300 3424 18352
rect 3476 18340 3482 18352
rect 5638 18343 5696 18349
rect 5638 18340 5650 18343
rect 3476 18312 5650 18340
rect 3476 18300 3482 18312
rect 5638 18309 5650 18312
rect 5684 18309 5696 18343
rect 7622 18343 7680 18349
rect 7622 18340 7634 18343
rect 5638 18303 5696 18309
rect 5736 18312 7634 18340
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18241 1823 18275
rect 1765 18235 1823 18241
rect 1949 18275 2007 18281
rect 1949 18241 1961 18275
rect 1995 18241 2007 18275
rect 1949 18235 2007 18241
rect 2409 18275 2467 18281
rect 2409 18241 2421 18275
rect 2455 18241 2467 18275
rect 2746 18272 2774 18300
rect 3697 18275 3755 18281
rect 3697 18272 3709 18275
rect 2746 18244 3709 18272
rect 2409 18235 2467 18241
rect 3697 18241 3709 18244
rect 3743 18241 3755 18275
rect 3697 18235 3755 18241
rect 3881 18275 3939 18281
rect 3881 18241 3893 18275
rect 3927 18272 3939 18275
rect 3927 18244 4568 18272
rect 3927 18241 3939 18244
rect 3881 18235 3939 18241
rect 1780 18136 1808 18235
rect 1854 18164 1860 18216
rect 1912 18204 1918 18216
rect 2424 18204 2452 18235
rect 1912 18176 2452 18204
rect 1912 18164 1918 18176
rect 2590 18136 2596 18148
rect 1780 18108 2596 18136
rect 2590 18096 2596 18108
rect 2648 18096 2654 18148
rect 4540 18145 4568 18244
rect 4614 18232 4620 18284
rect 4672 18272 4678 18284
rect 5736 18272 5764 18312
rect 7622 18309 7634 18312
rect 7668 18309 7680 18343
rect 7622 18303 7680 18309
rect 18506 18300 18512 18352
rect 18564 18300 18570 18352
rect 18693 18343 18751 18349
rect 18693 18309 18705 18343
rect 18739 18340 18751 18343
rect 19426 18340 19432 18352
rect 18739 18312 19432 18340
rect 18739 18309 18751 18312
rect 18693 18303 18751 18309
rect 19426 18300 19432 18312
rect 19484 18300 19490 18352
rect 4672 18244 5764 18272
rect 5905 18275 5963 18281
rect 4672 18232 4678 18244
rect 5905 18241 5917 18275
rect 5951 18272 5963 18275
rect 5994 18272 6000 18284
rect 5951 18244 6000 18272
rect 5951 18241 5963 18244
rect 5905 18235 5963 18241
rect 5994 18232 6000 18244
rect 6052 18272 6058 18284
rect 7377 18275 7435 18281
rect 7377 18272 7389 18275
rect 6052 18244 7389 18272
rect 6052 18232 6058 18244
rect 7377 18241 7389 18244
rect 7423 18241 7435 18275
rect 7377 18235 7435 18241
rect 8110 18232 8116 18284
rect 8168 18272 8174 18284
rect 8168 18244 12296 18272
rect 8168 18232 8174 18244
rect 12268 18216 12296 18244
rect 15470 18232 15476 18284
rect 15528 18232 15534 18284
rect 15746 18232 15752 18284
rect 15804 18232 15810 18284
rect 18524 18272 18552 18300
rect 19337 18275 19395 18281
rect 19337 18272 19349 18275
rect 18524 18244 19349 18272
rect 19337 18241 19349 18244
rect 19383 18241 19395 18275
rect 19337 18235 19395 18241
rect 19521 18275 19579 18281
rect 19521 18241 19533 18275
rect 19567 18272 19579 18275
rect 20438 18272 20444 18284
rect 19567 18244 20444 18272
rect 19567 18241 19579 18244
rect 19521 18235 19579 18241
rect 20438 18232 20444 18244
rect 20496 18232 20502 18284
rect 12250 18164 12256 18216
rect 12308 18204 12314 18216
rect 16022 18204 16028 18216
rect 12308 18176 16028 18204
rect 12308 18164 12314 18176
rect 16022 18164 16028 18176
rect 16080 18164 16086 18216
rect 18782 18164 18788 18216
rect 18840 18164 18846 18216
rect 4525 18139 4583 18145
rect 4525 18105 4537 18139
rect 4571 18105 4583 18139
rect 4525 18099 4583 18105
rect 8757 18139 8815 18145
rect 8757 18105 8769 18139
rect 8803 18136 8815 18139
rect 16206 18136 16212 18148
rect 8803 18108 16212 18136
rect 8803 18105 8815 18108
rect 8757 18099 8815 18105
rect 16206 18096 16212 18108
rect 16264 18096 16270 18148
rect 2501 18071 2559 18077
rect 2501 18037 2513 18071
rect 2547 18068 2559 18071
rect 3234 18068 3240 18080
rect 2547 18040 3240 18068
rect 2547 18037 2559 18040
rect 2501 18031 2559 18037
rect 3234 18028 3240 18040
rect 3292 18028 3298 18080
rect 15654 18028 15660 18080
rect 15712 18028 15718 18080
rect 18230 18028 18236 18080
rect 18288 18028 18294 18080
rect 1104 17978 22816 18000
rect 1104 17926 3664 17978
rect 3716 17926 3728 17978
rect 3780 17926 3792 17978
rect 3844 17926 3856 17978
rect 3908 17926 3920 17978
rect 3972 17926 9092 17978
rect 9144 17926 9156 17978
rect 9208 17926 9220 17978
rect 9272 17926 9284 17978
rect 9336 17926 9348 17978
rect 9400 17926 14520 17978
rect 14572 17926 14584 17978
rect 14636 17926 14648 17978
rect 14700 17926 14712 17978
rect 14764 17926 14776 17978
rect 14828 17926 19948 17978
rect 20000 17926 20012 17978
rect 20064 17926 20076 17978
rect 20128 17926 20140 17978
rect 20192 17926 20204 17978
rect 20256 17926 22816 17978
rect 1104 17904 22816 17926
rect 2961 17867 3019 17873
rect 2961 17864 2973 17867
rect 2746 17836 2973 17864
rect 1854 17620 1860 17672
rect 1912 17660 1918 17672
rect 1949 17663 2007 17669
rect 1949 17660 1961 17663
rect 1912 17632 1961 17660
rect 1912 17620 1918 17632
rect 1949 17629 1961 17632
rect 1995 17629 2007 17663
rect 1949 17623 2007 17629
rect 2225 17663 2283 17669
rect 2225 17629 2237 17663
rect 2271 17660 2283 17663
rect 2314 17660 2320 17672
rect 2271 17632 2320 17660
rect 2271 17629 2283 17632
rect 2225 17623 2283 17629
rect 2314 17620 2320 17632
rect 2372 17660 2378 17672
rect 2746 17660 2774 17836
rect 2961 17833 2973 17836
rect 3007 17864 3019 17867
rect 4614 17864 4620 17876
rect 3007 17836 4620 17864
rect 3007 17833 3019 17836
rect 2961 17827 3019 17833
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 5721 17867 5779 17873
rect 5721 17833 5733 17867
rect 5767 17864 5779 17867
rect 5994 17864 6000 17876
rect 5767 17836 6000 17864
rect 5767 17833 5779 17836
rect 5721 17827 5779 17833
rect 5994 17824 6000 17836
rect 6052 17824 6058 17876
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 11698 17864 11704 17876
rect 9732 17836 11704 17864
rect 9732 17824 9738 17836
rect 11698 17824 11704 17836
rect 11756 17824 11762 17876
rect 15470 17824 15476 17876
rect 15528 17824 15534 17876
rect 2372 17632 2774 17660
rect 2372 17620 2378 17632
rect 3050 17620 3056 17672
rect 3108 17620 3114 17672
rect 14829 17663 14887 17669
rect 14829 17629 14841 17663
rect 14875 17629 14887 17663
rect 14829 17623 14887 17629
rect 15013 17663 15071 17669
rect 15013 17629 15025 17663
rect 15059 17660 15071 17663
rect 15194 17660 15200 17672
rect 15059 17632 15200 17660
rect 15059 17629 15071 17632
rect 15013 17623 15071 17629
rect 2041 17595 2099 17601
rect 2041 17561 2053 17595
rect 2087 17592 2099 17595
rect 2498 17592 2504 17604
rect 2087 17564 2504 17592
rect 2087 17561 2099 17564
rect 2041 17555 2099 17561
rect 2498 17552 2504 17564
rect 2556 17552 2562 17604
rect 7009 17595 7067 17601
rect 7009 17561 7021 17595
rect 7055 17592 7067 17595
rect 10413 17595 10471 17601
rect 10413 17592 10425 17595
rect 7055 17564 10425 17592
rect 7055 17561 7067 17564
rect 7009 17555 7067 17561
rect 10413 17561 10425 17564
rect 10459 17592 10471 17595
rect 10594 17592 10600 17604
rect 10459 17564 10600 17592
rect 10459 17561 10471 17564
rect 10413 17555 10471 17561
rect 10594 17552 10600 17564
rect 10652 17552 10658 17604
rect 14844 17592 14872 17623
rect 15194 17620 15200 17632
rect 15252 17660 15258 17672
rect 15654 17660 15660 17672
rect 15252 17632 15660 17660
rect 15252 17620 15258 17632
rect 15654 17620 15660 17632
rect 15712 17660 15718 17672
rect 15749 17663 15807 17669
rect 15749 17660 15761 17663
rect 15712 17632 15761 17660
rect 15712 17620 15718 17632
rect 15749 17629 15761 17632
rect 15795 17629 15807 17663
rect 15749 17623 15807 17629
rect 16206 17620 16212 17672
rect 16264 17620 16270 17672
rect 19426 17620 19432 17672
rect 19484 17620 19490 17672
rect 15473 17595 15531 17601
rect 15473 17592 15485 17595
rect 14844 17564 15485 17592
rect 15473 17561 15485 17564
rect 15519 17592 15531 17595
rect 16390 17592 16396 17604
rect 15519 17564 16396 17592
rect 15519 17561 15531 17564
rect 15473 17555 15531 17561
rect 16390 17552 16396 17564
rect 16448 17552 16454 17604
rect 18782 17552 18788 17604
rect 18840 17592 18846 17604
rect 19242 17592 19248 17604
rect 18840 17564 19248 17592
rect 18840 17552 18846 17564
rect 19242 17552 19248 17564
rect 19300 17592 19306 17604
rect 19613 17595 19671 17601
rect 19613 17592 19625 17595
rect 19300 17564 19625 17592
rect 19300 17552 19306 17564
rect 19613 17561 19625 17564
rect 19659 17561 19671 17595
rect 19613 17555 19671 17561
rect 19794 17552 19800 17604
rect 19852 17552 19858 17604
rect 1946 17484 1952 17536
rect 2004 17524 2010 17536
rect 2409 17527 2467 17533
rect 2409 17524 2421 17527
rect 2004 17496 2421 17524
rect 2004 17484 2010 17496
rect 2409 17493 2421 17496
rect 2455 17493 2467 17527
rect 2409 17487 2467 17493
rect 2590 17484 2596 17536
rect 2648 17524 2654 17536
rect 2866 17524 2872 17536
rect 2648 17496 2872 17524
rect 2648 17484 2654 17496
rect 2866 17484 2872 17496
rect 2924 17484 2930 17536
rect 12894 17484 12900 17536
rect 12952 17524 12958 17536
rect 14921 17527 14979 17533
rect 14921 17524 14933 17527
rect 12952 17496 14933 17524
rect 12952 17484 12958 17496
rect 14921 17493 14933 17496
rect 14967 17493 14979 17527
rect 14921 17487 14979 17493
rect 15657 17527 15715 17533
rect 15657 17493 15669 17527
rect 15703 17524 15715 17527
rect 15746 17524 15752 17536
rect 15703 17496 15752 17524
rect 15703 17493 15715 17496
rect 15657 17487 15715 17493
rect 15746 17484 15752 17496
rect 15804 17484 15810 17536
rect 16301 17527 16359 17533
rect 16301 17493 16313 17527
rect 16347 17524 16359 17527
rect 16942 17524 16948 17536
rect 16347 17496 16948 17524
rect 16347 17493 16359 17496
rect 16301 17487 16359 17493
rect 16942 17484 16948 17496
rect 17000 17484 17006 17536
rect 1104 17434 22976 17456
rect 1104 17382 6378 17434
rect 6430 17382 6442 17434
rect 6494 17382 6506 17434
rect 6558 17382 6570 17434
rect 6622 17382 6634 17434
rect 6686 17382 11806 17434
rect 11858 17382 11870 17434
rect 11922 17382 11934 17434
rect 11986 17382 11998 17434
rect 12050 17382 12062 17434
rect 12114 17382 17234 17434
rect 17286 17382 17298 17434
rect 17350 17382 17362 17434
rect 17414 17382 17426 17434
rect 17478 17382 17490 17434
rect 17542 17382 22662 17434
rect 22714 17382 22726 17434
rect 22778 17382 22790 17434
rect 22842 17382 22854 17434
rect 22906 17382 22918 17434
rect 22970 17382 22976 17434
rect 1104 17360 22976 17382
rect 1946 17280 1952 17332
rect 2004 17280 2010 17332
rect 2866 17280 2872 17332
rect 2924 17320 2930 17332
rect 2924 17292 18552 17320
rect 2924 17280 2930 17292
rect 9922 17255 9980 17261
rect 9922 17252 9934 17255
rect 4172 17224 9934 17252
rect 2314 17144 2320 17196
rect 2372 17144 2378 17196
rect 3050 17144 3056 17196
rect 3108 17144 3114 17196
rect 3234 17144 3240 17196
rect 3292 17184 3298 17196
rect 4172 17184 4200 17224
rect 9922 17221 9934 17224
rect 9968 17221 9980 17255
rect 9922 17215 9980 17221
rect 14277 17255 14335 17261
rect 14277 17221 14289 17255
rect 14323 17252 14335 17255
rect 15194 17252 15200 17264
rect 14323 17224 15200 17252
rect 14323 17221 14335 17224
rect 14277 17215 14335 17221
rect 15194 17212 15200 17224
rect 15252 17212 15258 17264
rect 18524 17261 18552 17292
rect 19242 17280 19248 17332
rect 19300 17320 19306 17332
rect 19300 17292 20852 17320
rect 19300 17280 19306 17292
rect 18509 17255 18567 17261
rect 18509 17221 18521 17255
rect 18555 17221 18567 17255
rect 18509 17215 18567 17221
rect 19334 17212 19340 17264
rect 19392 17252 19398 17264
rect 19794 17252 19800 17264
rect 19392 17224 19800 17252
rect 19392 17212 19398 17224
rect 19794 17212 19800 17224
rect 19852 17212 19858 17264
rect 5730 17187 5788 17193
rect 5730 17184 5742 17187
rect 3292 17156 4200 17184
rect 4264 17156 5742 17184
rect 3292 17144 3298 17156
rect 2409 17119 2467 17125
rect 2409 17085 2421 17119
rect 2455 17116 2467 17119
rect 2498 17116 2504 17128
rect 2455 17088 2504 17116
rect 2455 17085 2467 17088
rect 2409 17079 2467 17085
rect 2498 17076 2504 17088
rect 2556 17076 2562 17128
rect 2593 17119 2651 17125
rect 2593 17085 2605 17119
rect 2639 17116 2651 17119
rect 4264 17116 4292 17156
rect 5730 17153 5742 17156
rect 5776 17153 5788 17187
rect 5730 17147 5788 17153
rect 5994 17144 6000 17196
rect 6052 17184 6058 17196
rect 7006 17184 7012 17196
rect 6052 17156 7012 17184
rect 6052 17144 6058 17156
rect 7006 17144 7012 17156
rect 7064 17184 7070 17196
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 7064 17156 7389 17184
rect 7064 17144 7070 17156
rect 7377 17153 7389 17156
rect 7423 17153 7435 17187
rect 7377 17147 7435 17153
rect 7466 17144 7472 17196
rect 7524 17184 7530 17196
rect 7633 17187 7691 17193
rect 7633 17184 7645 17187
rect 7524 17156 7645 17184
rect 7524 17144 7530 17156
rect 7633 17153 7645 17156
rect 7679 17153 7691 17187
rect 7633 17147 7691 17153
rect 11698 17144 11704 17196
rect 11756 17184 11762 17196
rect 12621 17187 12679 17193
rect 12621 17184 12633 17187
rect 11756 17156 12633 17184
rect 11756 17144 11762 17156
rect 12621 17153 12633 17156
rect 12667 17153 12679 17187
rect 12621 17147 12679 17153
rect 12894 17144 12900 17196
rect 12952 17144 12958 17196
rect 16482 17144 16488 17196
rect 16540 17184 16546 17196
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 16540 17156 16865 17184
rect 16540 17144 16546 17156
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 16853 17147 16911 17153
rect 17589 17187 17647 17193
rect 17589 17153 17601 17187
rect 17635 17184 17647 17187
rect 18230 17184 18236 17196
rect 17635 17156 18236 17184
rect 17635 17153 17647 17156
rect 17589 17147 17647 17153
rect 18230 17144 18236 17156
rect 18288 17144 18294 17196
rect 18690 17144 18696 17196
rect 18748 17184 18754 17196
rect 18969 17187 19027 17193
rect 18969 17184 18981 17187
rect 18748 17156 18981 17184
rect 18748 17144 18754 17156
rect 18969 17153 18981 17156
rect 19015 17153 19027 17187
rect 18969 17147 19027 17153
rect 19429 17187 19487 17193
rect 19429 17153 19441 17187
rect 19475 17184 19487 17187
rect 19518 17184 19524 17196
rect 19475 17156 19524 17184
rect 19475 17153 19487 17156
rect 19429 17147 19487 17153
rect 19518 17144 19524 17156
rect 19576 17144 19582 17196
rect 19610 17144 19616 17196
rect 19668 17184 19674 17196
rect 20824 17193 20852 17292
rect 20165 17187 20223 17193
rect 20165 17184 20177 17187
rect 19668 17156 20177 17184
rect 19668 17144 19674 17156
rect 20165 17153 20177 17156
rect 20211 17153 20223 17187
rect 20165 17147 20223 17153
rect 20349 17187 20407 17193
rect 20349 17153 20361 17187
rect 20395 17153 20407 17187
rect 20349 17147 20407 17153
rect 20809 17187 20867 17193
rect 20809 17153 20821 17187
rect 20855 17153 20867 17187
rect 20809 17147 20867 17153
rect 2639 17088 4292 17116
rect 2639 17085 2651 17088
rect 2593 17079 2651 17085
rect 9674 17076 9680 17128
rect 9732 17076 9738 17128
rect 12406 17088 17080 17116
rect 11057 17051 11115 17057
rect 11057 17017 11069 17051
rect 11103 17048 11115 17051
rect 12406 17048 12434 17088
rect 11103 17020 12434 17048
rect 11103 17017 11115 17020
rect 11057 17011 11115 17017
rect 14918 17008 14924 17060
rect 14976 17048 14982 17060
rect 16945 17051 17003 17057
rect 16945 17048 16957 17051
rect 14976 17020 16957 17048
rect 14976 17008 14982 17020
rect 16945 17017 16957 17020
rect 16991 17017 17003 17051
rect 17052 17048 17080 17088
rect 17678 17076 17684 17128
rect 17736 17076 17742 17128
rect 19705 17119 19763 17125
rect 19705 17085 19717 17119
rect 19751 17116 19763 17119
rect 20257 17119 20315 17125
rect 20257 17116 20269 17119
rect 19751 17088 20269 17116
rect 19751 17085 19763 17088
rect 19705 17079 19763 17085
rect 20257 17085 20269 17088
rect 20303 17085 20315 17119
rect 20257 17079 20315 17085
rect 20364 17116 20392 17147
rect 20990 17144 20996 17196
rect 21048 17144 21054 17196
rect 21008 17116 21036 17144
rect 20364 17088 21036 17116
rect 18230 17048 18236 17060
rect 17052 17020 18236 17048
rect 16945 17011 17003 17017
rect 18230 17008 18236 17020
rect 18288 17008 18294 17060
rect 3142 16940 3148 16992
rect 3200 16940 3206 16992
rect 4617 16983 4675 16989
rect 4617 16949 4629 16983
rect 4663 16980 4675 16983
rect 4982 16980 4988 16992
rect 4663 16952 4988 16980
rect 4663 16949 4675 16952
rect 4617 16943 4675 16949
rect 4982 16940 4988 16952
rect 5040 16940 5046 16992
rect 8754 16940 8760 16992
rect 8812 16940 8818 16992
rect 19702 16940 19708 16992
rect 19760 16980 19766 16992
rect 20364 16980 20392 17088
rect 19760 16952 20392 16980
rect 19760 16940 19766 16952
rect 20898 16940 20904 16992
rect 20956 16940 20962 16992
rect 1104 16890 22816 16912
rect 1104 16838 3664 16890
rect 3716 16838 3728 16890
rect 3780 16838 3792 16890
rect 3844 16838 3856 16890
rect 3908 16838 3920 16890
rect 3972 16838 9092 16890
rect 9144 16838 9156 16890
rect 9208 16838 9220 16890
rect 9272 16838 9284 16890
rect 9336 16838 9348 16890
rect 9400 16838 14520 16890
rect 14572 16838 14584 16890
rect 14636 16838 14648 16890
rect 14700 16838 14712 16890
rect 14764 16838 14776 16890
rect 14828 16838 19948 16890
rect 20000 16838 20012 16890
rect 20064 16838 20076 16890
rect 20128 16838 20140 16890
rect 20192 16838 20204 16890
rect 20256 16838 22816 16890
rect 1104 16816 22816 16838
rect 5994 16776 6000 16788
rect 4540 16748 6000 16776
rect 1946 16600 1952 16652
rect 2004 16640 2010 16652
rect 4540 16649 4568 16748
rect 5994 16736 6000 16748
rect 6052 16736 6058 16788
rect 16482 16736 16488 16788
rect 16540 16736 16546 16788
rect 18690 16736 18696 16788
rect 18748 16736 18754 16788
rect 11149 16711 11207 16717
rect 11149 16677 11161 16711
rect 11195 16677 11207 16711
rect 19981 16711 20039 16717
rect 19981 16708 19993 16711
rect 11149 16671 11207 16677
rect 17512 16680 19993 16708
rect 3421 16643 3479 16649
rect 2004 16612 2452 16640
rect 2004 16600 2010 16612
rect 2424 16581 2452 16612
rect 3421 16609 3433 16643
rect 3467 16640 3479 16643
rect 4525 16643 4583 16649
rect 3467 16612 4476 16640
rect 3467 16609 3479 16612
rect 3421 16603 3479 16609
rect 2225 16575 2283 16581
rect 2225 16541 2237 16575
rect 2271 16541 2283 16575
rect 2225 16535 2283 16541
rect 2409 16575 2467 16581
rect 2409 16541 2421 16575
rect 2455 16574 2467 16575
rect 3053 16575 3111 16581
rect 2455 16546 2489 16574
rect 2455 16541 2467 16546
rect 2409 16535 2467 16541
rect 3053 16541 3065 16575
rect 3099 16572 3111 16575
rect 3142 16572 3148 16584
rect 3099 16544 3148 16572
rect 3099 16541 3111 16544
rect 3053 16535 3111 16541
rect 1762 16464 1768 16516
rect 1820 16504 1826 16516
rect 2240 16504 2268 16535
rect 3142 16532 3148 16544
rect 3200 16532 3206 16584
rect 3234 16532 3240 16584
rect 3292 16572 3298 16584
rect 3878 16572 3884 16584
rect 3292 16544 3884 16572
rect 3292 16532 3298 16544
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 4448 16572 4476 16612
rect 4525 16609 4537 16643
rect 4571 16609 4583 16643
rect 4525 16603 4583 16609
rect 7006 16600 7012 16652
rect 7064 16600 7070 16652
rect 9674 16600 9680 16652
rect 9732 16640 9738 16652
rect 9769 16643 9827 16649
rect 9769 16640 9781 16643
rect 9732 16612 9781 16640
rect 9732 16600 9738 16612
rect 9769 16609 9781 16612
rect 9815 16609 9827 16643
rect 9769 16603 9827 16609
rect 7265 16575 7323 16581
rect 7265 16572 7277 16575
rect 4448 16544 7277 16572
rect 7265 16541 7277 16544
rect 7311 16541 7323 16575
rect 11164 16572 11192 16671
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 12069 16643 12127 16649
rect 12069 16640 12081 16643
rect 11756 16612 12081 16640
rect 11756 16600 11762 16612
rect 12069 16609 12081 16612
rect 12115 16609 12127 16643
rect 12069 16603 12127 16609
rect 16114 16600 16120 16652
rect 16172 16600 16178 16652
rect 17512 16649 17540 16680
rect 19981 16677 19993 16680
rect 20027 16677 20039 16711
rect 19981 16671 20039 16677
rect 16209 16643 16267 16649
rect 16209 16609 16221 16643
rect 16255 16640 16267 16643
rect 17497 16643 17555 16649
rect 16255 16612 17264 16640
rect 16255 16609 16267 16612
rect 16209 16603 16267 16609
rect 17236 16584 17264 16612
rect 17497 16609 17509 16643
rect 17543 16609 17555 16643
rect 17497 16603 17555 16609
rect 17678 16600 17684 16652
rect 17736 16600 17742 16652
rect 18417 16643 18475 16649
rect 18417 16640 18429 16643
rect 17880 16612 18429 16640
rect 15197 16575 15255 16581
rect 15197 16572 15209 16575
rect 11164 16544 15209 16572
rect 7265 16535 7323 16541
rect 15197 16541 15209 16544
rect 15243 16541 15255 16575
rect 15197 16535 15255 16541
rect 15289 16575 15347 16581
rect 15289 16541 15301 16575
rect 15335 16572 15347 16575
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 15335 16544 15853 16572
rect 15335 16541 15347 16544
rect 15289 16535 15347 16541
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 16022 16532 16028 16584
rect 16080 16532 16086 16584
rect 16301 16575 16359 16581
rect 16301 16541 16313 16575
rect 16347 16572 16359 16575
rect 17129 16575 17187 16581
rect 17129 16572 17141 16575
rect 16347 16544 17141 16572
rect 16347 16541 16359 16544
rect 16301 16535 16359 16541
rect 17129 16541 17141 16544
rect 17175 16541 17187 16575
rect 17129 16535 17187 16541
rect 4770 16507 4828 16513
rect 4770 16504 4782 16507
rect 1820 16476 2544 16504
rect 1820 16464 1826 16476
rect 2406 16396 2412 16448
rect 2464 16396 2470 16448
rect 2516 16436 2544 16476
rect 3804 16476 4782 16504
rect 3804 16436 3832 16476
rect 4770 16473 4782 16476
rect 4816 16473 4828 16507
rect 10036 16507 10094 16513
rect 10036 16504 10048 16507
rect 4770 16467 4828 16473
rect 4908 16476 10048 16504
rect 2516 16408 3832 16436
rect 3878 16396 3884 16448
rect 3936 16436 3942 16448
rect 4908 16436 4936 16476
rect 10036 16473 10048 16476
rect 10082 16473 10094 16507
rect 10036 16467 10094 16473
rect 3936 16408 4936 16436
rect 3936 16396 3942 16408
rect 5810 16396 5816 16448
rect 5868 16436 5874 16448
rect 5905 16439 5963 16445
rect 5905 16436 5917 16439
rect 5868 16408 5917 16436
rect 5868 16396 5874 16408
rect 5905 16405 5917 16408
rect 5951 16405 5963 16439
rect 5905 16399 5963 16405
rect 8386 16396 8392 16448
rect 8444 16396 8450 16448
rect 10060 16436 10088 16467
rect 12158 16464 12164 16516
rect 12216 16504 12222 16516
rect 12314 16507 12372 16513
rect 12314 16504 12326 16507
rect 12216 16476 12326 16504
rect 12216 16464 12222 16476
rect 12314 16473 12326 16476
rect 12360 16473 12372 16507
rect 14918 16504 14924 16516
rect 12314 16467 12372 16473
rect 12406 16476 14924 16504
rect 12406 16436 12434 16476
rect 14918 16464 14924 16476
rect 14976 16464 14982 16516
rect 17144 16504 17172 16535
rect 17218 16532 17224 16584
rect 17276 16572 17282 16584
rect 17405 16575 17463 16581
rect 17405 16572 17417 16575
rect 17276 16544 17417 16572
rect 17276 16532 17282 16544
rect 17405 16541 17417 16544
rect 17451 16572 17463 16575
rect 17880 16572 17908 16612
rect 18417 16609 18429 16612
rect 18463 16640 18475 16643
rect 19242 16640 19248 16652
rect 18463 16612 19248 16640
rect 18463 16609 18475 16612
rect 18417 16603 18475 16609
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 19610 16600 19616 16652
rect 19668 16640 19674 16652
rect 19668 16612 19840 16640
rect 19668 16600 19674 16612
rect 17451 16544 17908 16572
rect 17451 16541 17463 16544
rect 17405 16535 17463 16541
rect 18230 16532 18236 16584
rect 18288 16532 18294 16584
rect 18322 16532 18328 16584
rect 18380 16532 18386 16584
rect 18506 16532 18512 16584
rect 18564 16532 18570 16584
rect 19426 16532 19432 16584
rect 19484 16532 19490 16584
rect 19521 16575 19579 16581
rect 19521 16541 19533 16575
rect 19567 16572 19579 16575
rect 19567 16544 19656 16572
rect 19567 16541 19579 16544
rect 19521 16535 19579 16541
rect 18524 16504 18552 16532
rect 19628 16516 19656 16544
rect 19702 16532 19708 16584
rect 19760 16532 19766 16584
rect 19812 16581 19840 16612
rect 19797 16575 19855 16581
rect 19797 16541 19809 16575
rect 19843 16541 19855 16575
rect 19797 16535 19855 16541
rect 17144 16476 18552 16504
rect 19610 16464 19616 16516
rect 19668 16464 19674 16516
rect 10060 16408 12434 16436
rect 13449 16439 13507 16445
rect 13449 16405 13461 16439
rect 13495 16436 13507 16439
rect 15010 16436 15016 16448
rect 13495 16408 15016 16436
rect 13495 16405 13507 16408
rect 13449 16399 13507 16405
rect 15010 16396 15016 16408
rect 15068 16396 15074 16448
rect 1104 16346 22976 16368
rect 1104 16294 6378 16346
rect 6430 16294 6442 16346
rect 6494 16294 6506 16346
rect 6558 16294 6570 16346
rect 6622 16294 6634 16346
rect 6686 16294 11806 16346
rect 11858 16294 11870 16346
rect 11922 16294 11934 16346
rect 11986 16294 11998 16346
rect 12050 16294 12062 16346
rect 12114 16294 17234 16346
rect 17286 16294 17298 16346
rect 17350 16294 17362 16346
rect 17414 16294 17426 16346
rect 17478 16294 17490 16346
rect 17542 16294 22662 16346
rect 22714 16294 22726 16346
rect 22778 16294 22790 16346
rect 22842 16294 22854 16346
rect 22906 16294 22918 16346
rect 22970 16294 22976 16346
rect 1104 16272 22976 16294
rect 1762 16192 1768 16244
rect 1820 16192 1826 16244
rect 2406 16192 2412 16244
rect 2464 16232 2470 16244
rect 2958 16232 2964 16244
rect 2464 16204 2964 16232
rect 2464 16192 2470 16204
rect 2958 16192 2964 16204
rect 3016 16192 3022 16244
rect 3234 16232 3240 16244
rect 3068 16204 3240 16232
rect 2314 16164 2320 16176
rect 1872 16136 2320 16164
rect 1872 16105 1900 16136
rect 2314 16124 2320 16136
rect 2372 16164 2378 16176
rect 2590 16164 2596 16176
rect 2372 16136 2596 16164
rect 2372 16124 2378 16136
rect 2590 16124 2596 16136
rect 2648 16124 2654 16176
rect 3068 16164 3096 16204
rect 3234 16192 3240 16204
rect 3292 16192 3298 16244
rect 4062 16192 4068 16244
rect 4120 16232 4126 16244
rect 4120 16204 19104 16232
rect 4120 16192 4126 16204
rect 2700 16136 3096 16164
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16065 1915 16099
rect 1857 16059 1915 16065
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16096 2099 16099
rect 2498 16096 2504 16108
rect 2087 16068 2504 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 2498 16056 2504 16068
rect 2556 16096 2562 16108
rect 2700 16096 2728 16136
rect 3142 16124 3148 16176
rect 3200 16164 3206 16176
rect 3200 16136 3648 16164
rect 3200 16124 3206 16136
rect 2556 16068 2728 16096
rect 2556 16056 2562 16068
rect 2866 16056 2872 16108
rect 2924 16056 2930 16108
rect 3620 16105 3648 16136
rect 8294 16124 8300 16176
rect 8352 16164 8358 16176
rect 9309 16167 9367 16173
rect 9309 16164 9321 16167
rect 8352 16136 9321 16164
rect 8352 16124 8358 16136
rect 9309 16133 9321 16136
rect 9355 16133 9367 16167
rect 18506 16164 18512 16176
rect 9309 16127 9367 16133
rect 17236 16136 18512 16164
rect 3421 16099 3479 16105
rect 3421 16065 3433 16099
rect 3467 16065 3479 16099
rect 3421 16059 3479 16065
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16065 3663 16099
rect 3605 16059 3663 16065
rect 1581 16031 1639 16037
rect 1581 15997 1593 16031
rect 1627 16028 1639 16031
rect 2130 16028 2136 16040
rect 1627 16000 2136 16028
rect 1627 15997 1639 16000
rect 1581 15991 1639 15997
rect 2130 15988 2136 16000
rect 2188 16028 2194 16040
rect 3436 16028 3464 16059
rect 16942 16056 16948 16108
rect 17000 16056 17006 16108
rect 17126 16056 17132 16108
rect 17184 16056 17190 16108
rect 17236 16105 17264 16136
rect 18506 16124 18512 16136
rect 18564 16124 18570 16176
rect 19076 16173 19104 16204
rect 19061 16167 19119 16173
rect 19061 16133 19073 16167
rect 19107 16133 19119 16167
rect 19061 16127 19119 16133
rect 17221 16099 17279 16105
rect 17221 16065 17233 16099
rect 17267 16065 17279 16099
rect 17221 16059 17279 16065
rect 17405 16099 17463 16105
rect 17405 16065 17417 16099
rect 17451 16096 17463 16099
rect 18693 16099 18751 16105
rect 18693 16096 18705 16099
rect 17451 16068 18705 16096
rect 17451 16065 17463 16068
rect 17405 16059 17463 16065
rect 18693 16065 18705 16068
rect 18739 16065 18751 16099
rect 18693 16059 18751 16065
rect 19334 16056 19340 16108
rect 19392 16096 19398 16108
rect 19429 16099 19487 16105
rect 19429 16096 19441 16099
rect 19392 16068 19441 16096
rect 19392 16056 19398 16068
rect 19429 16065 19441 16068
rect 19475 16065 19487 16099
rect 19429 16059 19487 16065
rect 19518 16056 19524 16108
rect 19576 16056 19582 16108
rect 19889 16099 19947 16105
rect 19889 16065 19901 16099
rect 19935 16096 19947 16099
rect 20898 16096 20904 16108
rect 19935 16068 20904 16096
rect 19935 16065 19947 16068
rect 19889 16059 19947 16065
rect 20898 16056 20904 16068
rect 20956 16056 20962 16108
rect 2188 16000 3464 16028
rect 2188 15988 2194 16000
rect 12342 15988 12348 16040
rect 12400 16028 12406 16040
rect 12621 16031 12679 16037
rect 12621 16028 12633 16031
rect 12400 16000 12633 16028
rect 12400 15988 12406 16000
rect 12621 15997 12633 16000
rect 12667 15997 12679 16031
rect 12621 15991 12679 15997
rect 12897 16031 12955 16037
rect 12897 15997 12909 16031
rect 12943 16028 12955 16031
rect 16758 16028 16764 16040
rect 12943 16000 16764 16028
rect 12943 15997 12955 16000
rect 12897 15991 12955 15997
rect 16758 15988 16764 16000
rect 16816 15988 16822 16040
rect 18509 16031 18567 16037
rect 18509 15997 18521 16031
rect 18555 16028 18567 16031
rect 18598 16028 18604 16040
rect 18555 16000 18604 16028
rect 18555 15997 18567 16000
rect 18509 15991 18567 15997
rect 18598 15988 18604 16000
rect 18656 15988 18662 16040
rect 2682 15920 2688 15972
rect 2740 15920 2746 15972
rect 2958 15920 2964 15972
rect 3016 15960 3022 15972
rect 7466 15960 7472 15972
rect 3016 15932 7472 15960
rect 3016 15920 3022 15932
rect 7466 15920 7472 15932
rect 7524 15920 7530 15972
rect 16114 15920 16120 15972
rect 16172 15960 16178 15972
rect 17037 15963 17095 15969
rect 17037 15960 17049 15963
rect 16172 15932 17049 15960
rect 16172 15920 16178 15932
rect 17037 15929 17049 15932
rect 17083 15960 17095 15963
rect 18322 15960 18328 15972
rect 17083 15932 18328 15960
rect 17083 15929 17095 15932
rect 17037 15923 17095 15929
rect 18322 15920 18328 15932
rect 18380 15920 18386 15972
rect 3513 15895 3571 15901
rect 3513 15861 3525 15895
rect 3559 15892 3571 15895
rect 9674 15892 9680 15904
rect 3559 15864 9680 15892
rect 3559 15861 3571 15864
rect 3513 15855 3571 15861
rect 9674 15852 9680 15864
rect 9732 15852 9738 15904
rect 10594 15852 10600 15904
rect 10652 15852 10658 15904
rect 14185 15895 14243 15901
rect 14185 15861 14197 15895
rect 14231 15892 14243 15895
rect 16850 15892 16856 15904
rect 14231 15864 16856 15892
rect 14231 15861 14243 15864
rect 14185 15855 14243 15861
rect 16850 15852 16856 15864
rect 16908 15852 16914 15904
rect 1104 15802 22816 15824
rect 1104 15750 3664 15802
rect 3716 15750 3728 15802
rect 3780 15750 3792 15802
rect 3844 15750 3856 15802
rect 3908 15750 3920 15802
rect 3972 15750 9092 15802
rect 9144 15750 9156 15802
rect 9208 15750 9220 15802
rect 9272 15750 9284 15802
rect 9336 15750 9348 15802
rect 9400 15750 14520 15802
rect 14572 15750 14584 15802
rect 14636 15750 14648 15802
rect 14700 15750 14712 15802
rect 14764 15750 14776 15802
rect 14828 15750 19948 15802
rect 20000 15750 20012 15802
rect 20064 15750 20076 15802
rect 20128 15750 20140 15802
rect 20192 15750 20204 15802
rect 20256 15750 22816 15802
rect 1104 15728 22816 15750
rect 2130 15648 2136 15700
rect 2188 15648 2194 15700
rect 16758 15648 16764 15700
rect 16816 15688 16822 15700
rect 17037 15691 17095 15697
rect 17037 15688 17049 15691
rect 16816 15660 17049 15688
rect 16816 15648 16822 15660
rect 17037 15657 17049 15660
rect 17083 15657 17095 15691
rect 17037 15651 17095 15657
rect 17126 15648 17132 15700
rect 17184 15688 17190 15700
rect 17221 15691 17279 15697
rect 17221 15688 17233 15691
rect 17184 15660 17233 15688
rect 17184 15648 17190 15660
rect 17221 15657 17233 15660
rect 17267 15657 17279 15691
rect 17221 15651 17279 15657
rect 2498 15580 2504 15632
rect 2556 15580 2562 15632
rect 19705 15623 19763 15629
rect 19705 15589 19717 15623
rect 19751 15620 19763 15623
rect 20070 15620 20076 15632
rect 19751 15592 20076 15620
rect 19751 15589 19763 15592
rect 19705 15583 19763 15589
rect 20070 15580 20076 15592
rect 20128 15580 20134 15632
rect 2314 15512 2320 15564
rect 2372 15512 2378 15564
rect 2409 15555 2467 15561
rect 2409 15521 2421 15555
rect 2455 15552 2467 15555
rect 2516 15552 2544 15580
rect 2455 15524 2544 15552
rect 2455 15521 2467 15524
rect 2409 15515 2467 15521
rect 2590 15512 2596 15564
rect 2648 15552 2654 15564
rect 3050 15552 3056 15564
rect 2648 15524 3056 15552
rect 2648 15512 2654 15524
rect 3050 15512 3056 15524
rect 3108 15552 3114 15564
rect 4062 15552 4068 15564
rect 3108 15524 4068 15552
rect 3108 15512 3114 15524
rect 4062 15512 4068 15524
rect 4120 15512 4126 15564
rect 1946 15444 1952 15496
rect 2004 15484 2010 15496
rect 2501 15487 2559 15493
rect 2501 15484 2513 15487
rect 2004 15456 2513 15484
rect 2004 15444 2010 15456
rect 2501 15453 2513 15456
rect 2547 15484 2559 15487
rect 2682 15484 2688 15496
rect 2547 15456 2688 15484
rect 2547 15453 2559 15456
rect 2501 15447 2559 15453
rect 2682 15444 2688 15456
rect 2740 15444 2746 15496
rect 9582 15444 9588 15496
rect 9640 15444 9646 15496
rect 9674 15444 9680 15496
rect 9732 15484 9738 15496
rect 9841 15487 9899 15493
rect 9841 15484 9853 15487
rect 9732 15456 9853 15484
rect 9732 15444 9738 15456
rect 9841 15453 9853 15456
rect 9887 15453 9899 15487
rect 9841 15447 9899 15453
rect 12342 15444 12348 15496
rect 12400 15444 12406 15496
rect 15378 15444 15384 15496
rect 15436 15484 15442 15496
rect 15933 15487 15991 15493
rect 15933 15484 15945 15487
rect 15436 15456 15945 15484
rect 15436 15444 15442 15456
rect 15933 15453 15945 15456
rect 15979 15453 15991 15487
rect 15933 15447 15991 15453
rect 16022 15444 16028 15496
rect 16080 15484 16086 15496
rect 16080 15456 17448 15484
rect 16080 15444 16086 15456
rect 12612 15419 12670 15425
rect 12612 15385 12624 15419
rect 12658 15416 12670 15419
rect 15102 15416 15108 15428
rect 12658 15388 15108 15416
rect 12658 15385 12670 15388
rect 12612 15379 12670 15385
rect 15102 15376 15108 15388
rect 15160 15376 15166 15428
rect 16482 15376 16488 15428
rect 16540 15376 16546 15428
rect 17420 15425 17448 15456
rect 18322 15444 18328 15496
rect 18380 15484 18386 15496
rect 19334 15484 19340 15496
rect 18380 15456 19340 15484
rect 18380 15444 18386 15456
rect 19334 15444 19340 15456
rect 19392 15484 19398 15496
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 19392 15456 19441 15484
rect 19392 15444 19398 15456
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 17405 15419 17463 15425
rect 17405 15385 17417 15419
rect 17451 15385 17463 15419
rect 17405 15379 17463 15385
rect 19702 15376 19708 15428
rect 19760 15376 19766 15428
rect 10870 15308 10876 15360
rect 10928 15348 10934 15360
rect 10965 15351 11023 15357
rect 10965 15348 10977 15351
rect 10928 15320 10977 15348
rect 10928 15308 10934 15320
rect 10965 15317 10977 15320
rect 11011 15317 11023 15351
rect 10965 15311 11023 15317
rect 13725 15351 13783 15357
rect 13725 15317 13737 15351
rect 13771 15348 13783 15351
rect 15562 15348 15568 15360
rect 13771 15320 15568 15348
rect 13771 15317 13783 15320
rect 13725 15311 13783 15317
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 17205 15351 17263 15357
rect 17205 15317 17217 15351
rect 17251 15348 17263 15351
rect 17586 15348 17592 15360
rect 17251 15320 17592 15348
rect 17251 15317 17263 15320
rect 17205 15311 17263 15317
rect 17586 15308 17592 15320
rect 17644 15308 17650 15360
rect 18782 15308 18788 15360
rect 18840 15348 18846 15360
rect 19521 15351 19579 15357
rect 19521 15348 19533 15351
rect 18840 15320 19533 15348
rect 18840 15308 18846 15320
rect 19521 15317 19533 15320
rect 19567 15317 19579 15351
rect 19521 15311 19579 15317
rect 1104 15258 22976 15280
rect 1104 15206 6378 15258
rect 6430 15206 6442 15258
rect 6494 15206 6506 15258
rect 6558 15206 6570 15258
rect 6622 15206 6634 15258
rect 6686 15206 11806 15258
rect 11858 15206 11870 15258
rect 11922 15206 11934 15258
rect 11986 15206 11998 15258
rect 12050 15206 12062 15258
rect 12114 15206 17234 15258
rect 17286 15206 17298 15258
rect 17350 15206 17362 15258
rect 17414 15206 17426 15258
rect 17478 15206 17490 15258
rect 17542 15206 22662 15258
rect 22714 15206 22726 15258
rect 22778 15206 22790 15258
rect 22842 15206 22854 15258
rect 22906 15206 22918 15258
rect 22970 15206 22976 15258
rect 1104 15184 22976 15206
rect 2498 15104 2504 15156
rect 2556 15144 2562 15156
rect 2556 15116 2820 15144
rect 2556 15104 2562 15116
rect 2590 15076 2596 15088
rect 2332 15048 2596 15076
rect 2332 15017 2360 15048
rect 2590 15036 2596 15048
rect 2648 15036 2654 15088
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 14977 2375 15011
rect 2317 14971 2375 14977
rect 2406 14968 2412 15020
rect 2464 15008 2470 15020
rect 2792 15017 2820 15116
rect 2866 15104 2872 15156
rect 2924 15144 2930 15156
rect 3789 15147 3847 15153
rect 3789 15144 3801 15147
rect 2924 15116 3801 15144
rect 2924 15104 2930 15116
rect 3789 15113 3801 15116
rect 3835 15144 3847 15147
rect 8110 15144 8116 15156
rect 3835 15116 8116 15144
rect 3835 15113 3847 15116
rect 3789 15107 3847 15113
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 15102 15104 15108 15156
rect 15160 15144 15166 15156
rect 15289 15147 15347 15153
rect 15289 15144 15301 15147
rect 15160 15116 15301 15144
rect 15160 15104 15166 15116
rect 15289 15113 15301 15116
rect 15335 15113 15347 15147
rect 15289 15107 15347 15113
rect 17126 15104 17132 15156
rect 17184 15144 17190 15156
rect 17221 15147 17279 15153
rect 17221 15144 17233 15147
rect 17184 15116 17233 15144
rect 17184 15104 17190 15116
rect 17221 15113 17233 15116
rect 17267 15113 17279 15147
rect 17221 15107 17279 15113
rect 18785 15147 18843 15153
rect 18785 15113 18797 15147
rect 18831 15144 18843 15147
rect 18874 15144 18880 15156
rect 18831 15116 18880 15144
rect 18831 15113 18843 15116
rect 18785 15107 18843 15113
rect 18874 15104 18880 15116
rect 18932 15144 18938 15156
rect 19518 15144 19524 15156
rect 18932 15116 19524 15144
rect 18932 15104 18938 15116
rect 19518 15104 19524 15116
rect 19576 15104 19582 15156
rect 20073 15147 20131 15153
rect 20073 15113 20085 15147
rect 20119 15113 20131 15147
rect 20073 15107 20131 15113
rect 2961 15079 3019 15085
rect 2961 15045 2973 15079
rect 3007 15076 3019 15079
rect 7898 15079 7956 15085
rect 7898 15076 7910 15079
rect 3007 15048 7910 15076
rect 3007 15045 3019 15048
rect 2961 15039 3019 15045
rect 7898 15045 7910 15048
rect 7944 15045 7956 15079
rect 7898 15039 7956 15045
rect 12158 15036 12164 15088
rect 12216 15076 12222 15088
rect 20088 15076 20116 15107
rect 12216 15048 20116 15076
rect 12216 15036 12222 15048
rect 2501 15011 2559 15017
rect 2501 15008 2513 15011
rect 2464 14980 2513 15008
rect 2464 14968 2470 14980
rect 2501 14977 2513 14980
rect 2547 14977 2559 15011
rect 2501 14971 2559 14977
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 14977 2835 15011
rect 2777 14971 2835 14977
rect 3510 14968 3516 15020
rect 3568 14968 3574 15020
rect 4062 14968 4068 15020
rect 4120 15008 4126 15020
rect 4689 15011 4747 15017
rect 4689 15008 4701 15011
rect 4120 14980 4701 15008
rect 4120 14968 4126 14980
rect 4689 14977 4701 14980
rect 4735 14977 4747 15011
rect 4689 14971 4747 14977
rect 12612 15011 12670 15017
rect 12612 14977 12624 15011
rect 12658 15008 12670 15011
rect 13722 15008 13728 15020
rect 12658 14980 13728 15008
rect 12658 14977 12670 14980
rect 12612 14971 12670 14977
rect 13722 14968 13728 14980
rect 13780 14968 13786 15020
rect 15473 15011 15531 15017
rect 15473 14977 15485 15011
rect 15519 14977 15531 15011
rect 15473 14971 15531 14977
rect 4433 14943 4491 14949
rect 4433 14909 4445 14943
rect 4479 14909 4491 14943
rect 4433 14903 4491 14909
rect 4448 14804 4476 14903
rect 7650 14900 7656 14952
rect 7708 14900 7714 14952
rect 12342 14900 12348 14952
rect 12400 14900 12406 14952
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 15488 14940 15516 14971
rect 15562 14968 15568 15020
rect 15620 14968 15626 15020
rect 15749 15011 15807 15017
rect 15749 14977 15761 15011
rect 15795 14977 15807 15011
rect 15749 14971 15807 14977
rect 15841 15011 15899 15017
rect 15841 14977 15853 15011
rect 15887 15008 15899 15011
rect 16114 15008 16120 15020
rect 15887 14980 16120 15008
rect 15887 14977 15899 14980
rect 15841 14971 15899 14977
rect 13688 14912 15516 14940
rect 15764 14940 15792 14971
rect 16114 14968 16120 14980
rect 16172 14968 16178 15020
rect 16758 14968 16764 15020
rect 16816 15008 16822 15020
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 16816 14980 16865 15008
rect 16816 14968 16822 14980
rect 16853 14977 16865 14980
rect 16899 15008 16911 15011
rect 17954 15008 17960 15020
rect 16899 14980 17960 15008
rect 16899 14977 16911 14980
rect 16853 14971 16911 14977
rect 17954 14968 17960 14980
rect 18012 14968 18018 15020
rect 18046 14968 18052 15020
rect 18104 15008 18110 15020
rect 18506 15008 18512 15020
rect 18104 14980 18512 15008
rect 18104 14968 18110 14980
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 19334 14968 19340 15020
rect 19392 14968 19398 15020
rect 20070 14968 20076 15020
rect 20128 14968 20134 15020
rect 16482 14940 16488 14952
rect 15764 14912 16488 14940
rect 13688 14900 13694 14912
rect 15378 14832 15384 14884
rect 15436 14872 15442 14884
rect 15764 14872 15792 14912
rect 16482 14900 16488 14912
rect 16540 14900 16546 14952
rect 16945 14943 17003 14949
rect 16945 14909 16957 14943
rect 16991 14940 17003 14943
rect 16991 14912 19196 14940
rect 16991 14909 17003 14912
rect 16945 14903 17003 14909
rect 18782 14872 18788 14884
rect 15436 14844 15792 14872
rect 16776 14844 18788 14872
rect 15436 14832 15442 14844
rect 5626 14804 5632 14816
rect 4448 14776 5632 14804
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 5813 14807 5871 14813
rect 5813 14773 5825 14807
rect 5859 14804 5871 14807
rect 5994 14804 6000 14816
rect 5859 14776 6000 14804
rect 5859 14773 5871 14776
rect 5813 14767 5871 14773
rect 5994 14764 6000 14776
rect 6052 14764 6058 14816
rect 8846 14764 8852 14816
rect 8904 14804 8910 14816
rect 9033 14807 9091 14813
rect 9033 14804 9045 14807
rect 8904 14776 9045 14804
rect 8904 14764 8910 14776
rect 9033 14773 9045 14776
rect 9079 14773 9091 14807
rect 9033 14767 9091 14773
rect 13725 14807 13783 14813
rect 13725 14773 13737 14807
rect 13771 14804 13783 14807
rect 16776 14804 16804 14844
rect 18782 14832 18788 14844
rect 18840 14832 18846 14884
rect 19168 14872 19196 14912
rect 19242 14900 19248 14952
rect 19300 14900 19306 14952
rect 19518 14900 19524 14952
rect 19576 14940 19582 14952
rect 20349 14943 20407 14949
rect 20349 14940 20361 14943
rect 19576 14912 20361 14940
rect 19576 14900 19582 14912
rect 20349 14909 20361 14912
rect 20395 14909 20407 14943
rect 20349 14903 20407 14909
rect 19426 14872 19432 14884
rect 19168 14844 19432 14872
rect 19426 14832 19432 14844
rect 19484 14832 19490 14884
rect 19794 14832 19800 14884
rect 19852 14872 19858 14884
rect 20165 14875 20223 14881
rect 20165 14872 20177 14875
rect 19852 14844 20177 14872
rect 19852 14832 19858 14844
rect 20165 14841 20177 14844
rect 20211 14841 20223 14875
rect 20165 14835 20223 14841
rect 13771 14776 16804 14804
rect 13771 14773 13783 14776
rect 13725 14767 13783 14773
rect 16850 14764 16856 14816
rect 16908 14764 16914 14816
rect 1104 14714 22816 14736
rect 1104 14662 3664 14714
rect 3716 14662 3728 14714
rect 3780 14662 3792 14714
rect 3844 14662 3856 14714
rect 3908 14662 3920 14714
rect 3972 14662 9092 14714
rect 9144 14662 9156 14714
rect 9208 14662 9220 14714
rect 9272 14662 9284 14714
rect 9336 14662 9348 14714
rect 9400 14662 14520 14714
rect 14572 14662 14584 14714
rect 14636 14662 14648 14714
rect 14700 14662 14712 14714
rect 14764 14662 14776 14714
rect 14828 14662 19948 14714
rect 20000 14662 20012 14714
rect 20064 14662 20076 14714
rect 20128 14662 20140 14714
rect 20192 14662 20204 14714
rect 20256 14662 22816 14714
rect 1104 14640 22816 14662
rect 2222 14560 2228 14612
rect 2280 14560 2286 14612
rect 2317 14603 2375 14609
rect 2317 14569 2329 14603
rect 2363 14600 2375 14603
rect 4062 14600 4068 14612
rect 2363 14572 4068 14600
rect 2363 14569 2375 14572
rect 2317 14563 2375 14569
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 12250 14560 12256 14612
rect 12308 14600 12314 14612
rect 13354 14600 13360 14612
rect 12308 14572 13360 14600
rect 12308 14560 12314 14572
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 16482 14560 16488 14612
rect 16540 14600 16546 14612
rect 17034 14600 17040 14612
rect 16540 14572 17040 14600
rect 16540 14560 16546 14572
rect 17034 14560 17040 14572
rect 17092 14600 17098 14612
rect 18598 14600 18604 14612
rect 17092 14572 18604 14600
rect 17092 14560 17098 14572
rect 18598 14560 18604 14572
rect 18656 14560 18662 14612
rect 19610 14560 19616 14612
rect 19668 14560 19674 14612
rect 19794 14560 19800 14612
rect 19852 14560 19858 14612
rect 2130 14492 2136 14544
rect 2188 14492 2194 14544
rect 15841 14535 15899 14541
rect 15841 14501 15853 14535
rect 15887 14501 15899 14535
rect 17586 14532 17592 14544
rect 15841 14495 15899 14501
rect 16132 14504 17592 14532
rect 2148 14464 2176 14492
rect 2409 14467 2467 14473
rect 2409 14464 2421 14467
rect 2148 14436 2421 14464
rect 2409 14433 2421 14436
rect 2455 14433 2467 14467
rect 2409 14427 2467 14433
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 2498 14396 2504 14408
rect 2179 14368 2504 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 5626 14356 5632 14408
rect 5684 14356 5690 14408
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14396 8171 14399
rect 8202 14396 8208 14408
rect 8159 14368 8208 14396
rect 8159 14365 8171 14368
rect 8113 14359 8171 14365
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 9493 14399 9551 14405
rect 9493 14365 9505 14399
rect 9539 14396 9551 14399
rect 9582 14396 9588 14408
rect 9539 14368 9588 14396
rect 9539 14365 9551 14368
rect 9493 14359 9551 14365
rect 9582 14356 9588 14368
rect 9640 14356 9646 14408
rect 9769 14399 9827 14405
rect 9769 14365 9781 14399
rect 9815 14396 9827 14399
rect 11054 14396 11060 14408
rect 9815 14368 11060 14396
rect 9815 14365 9827 14368
rect 9769 14359 9827 14365
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 12342 14356 12348 14408
rect 12400 14356 12406 14408
rect 12612 14399 12670 14405
rect 12612 14365 12624 14399
rect 12658 14396 12670 14399
rect 15856 14396 15884 14495
rect 16132 14405 16160 14504
rect 17586 14492 17592 14504
rect 17644 14492 17650 14544
rect 18782 14492 18788 14544
rect 18840 14492 18846 14544
rect 19628 14532 19656 14560
rect 20254 14532 20260 14544
rect 19628 14504 20260 14532
rect 20254 14492 20260 14504
rect 20312 14492 20318 14544
rect 16666 14424 16672 14476
rect 16724 14464 16730 14476
rect 16853 14467 16911 14473
rect 16853 14464 16865 14467
rect 16724 14436 16865 14464
rect 16724 14424 16730 14436
rect 16853 14433 16865 14436
rect 16899 14433 16911 14467
rect 18800 14464 18828 14492
rect 18800 14436 19656 14464
rect 16853 14427 16911 14433
rect 12658 14368 15884 14396
rect 16117 14399 16175 14405
rect 12658 14365 12670 14368
rect 12612 14359 12670 14365
rect 16117 14365 16129 14399
rect 16163 14365 16175 14399
rect 16117 14359 16175 14365
rect 16758 14356 16764 14408
rect 16816 14356 16822 14408
rect 16945 14399 17003 14405
rect 16945 14365 16957 14399
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 4614 14288 4620 14340
rect 4672 14328 4678 14340
rect 5362 14331 5420 14337
rect 5362 14328 5374 14331
rect 4672 14300 5374 14328
rect 4672 14288 4678 14300
rect 5362 14297 5374 14300
rect 5408 14297 5420 14331
rect 5362 14291 5420 14297
rect 7558 14288 7564 14340
rect 7616 14328 7622 14340
rect 7846 14331 7904 14337
rect 7846 14328 7858 14331
rect 7616 14300 7858 14328
rect 7616 14288 7622 14300
rect 7846 14297 7858 14300
rect 7892 14297 7904 14331
rect 7846 14291 7904 14297
rect 4154 14220 4160 14272
rect 4212 14260 4218 14272
rect 4249 14263 4307 14269
rect 4249 14260 4261 14263
rect 4212 14232 4261 14260
rect 4212 14220 4218 14232
rect 4249 14229 4261 14232
rect 4295 14229 4307 14263
rect 4249 14223 4307 14229
rect 5902 14220 5908 14272
rect 5960 14260 5966 14272
rect 6733 14263 6791 14269
rect 6733 14260 6745 14263
rect 5960 14232 6745 14260
rect 5960 14220 5966 14232
rect 6733 14229 6745 14232
rect 6779 14229 6791 14263
rect 9600 14260 9628 14356
rect 14642 14328 14648 14340
rect 12406 14300 14648 14328
rect 9766 14260 9772 14272
rect 9600 14232 9772 14260
rect 6733 14223 6791 14229
rect 9766 14220 9772 14232
rect 9824 14220 9830 14272
rect 10686 14220 10692 14272
rect 10744 14260 10750 14272
rect 11057 14263 11115 14269
rect 11057 14260 11069 14263
rect 10744 14232 11069 14260
rect 10744 14220 10750 14232
rect 11057 14229 11069 14232
rect 11103 14260 11115 14263
rect 12406 14260 12434 14300
rect 14642 14288 14648 14300
rect 14700 14328 14706 14340
rect 15746 14328 15752 14340
rect 14700 14300 15752 14328
rect 14700 14288 14706 14300
rect 15746 14288 15752 14300
rect 15804 14288 15810 14340
rect 15841 14331 15899 14337
rect 15841 14297 15853 14331
rect 15887 14328 15899 14331
rect 15887 14300 16620 14328
rect 15887 14297 15899 14300
rect 15841 14291 15899 14297
rect 11103 14232 12434 14260
rect 13725 14263 13783 14269
rect 11103 14229 11115 14232
rect 11057 14223 11115 14229
rect 13725 14229 13737 14263
rect 13771 14260 13783 14263
rect 15654 14260 15660 14272
rect 13771 14232 15660 14260
rect 13771 14229 13783 14232
rect 13725 14223 13783 14229
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 16022 14220 16028 14272
rect 16080 14220 16086 14272
rect 16592 14269 16620 14300
rect 16850 14288 16856 14340
rect 16908 14328 16914 14340
rect 16960 14328 16988 14359
rect 17034 14356 17040 14408
rect 17092 14356 17098 14408
rect 17589 14399 17647 14405
rect 17589 14365 17601 14399
rect 17635 14365 17647 14399
rect 17589 14359 17647 14365
rect 17773 14399 17831 14405
rect 17773 14365 17785 14399
rect 17819 14396 17831 14399
rect 17954 14396 17960 14408
rect 17819 14368 17960 14396
rect 17819 14365 17831 14368
rect 17773 14359 17831 14365
rect 17604 14328 17632 14359
rect 17954 14356 17960 14368
rect 18012 14396 18018 14408
rect 18417 14399 18475 14405
rect 18417 14396 18429 14399
rect 18012 14368 18429 14396
rect 18012 14356 18018 14368
rect 18417 14365 18429 14368
rect 18463 14365 18475 14399
rect 18417 14359 18475 14365
rect 18598 14356 18604 14408
rect 18656 14396 18662 14408
rect 18782 14396 18788 14408
rect 18656 14368 18788 14396
rect 18656 14356 18662 14368
rect 18782 14356 18788 14368
rect 18840 14396 18846 14408
rect 19518 14396 19524 14408
rect 18840 14368 19524 14396
rect 18840 14356 18846 14368
rect 19518 14356 19524 14368
rect 19576 14356 19582 14408
rect 16908 14300 17632 14328
rect 19429 14331 19487 14337
rect 16908 14288 16914 14300
rect 19429 14297 19441 14331
rect 19475 14328 19487 14331
rect 19628 14328 19656 14436
rect 20438 14328 20444 14340
rect 19475 14300 20444 14328
rect 19475 14297 19487 14300
rect 19429 14291 19487 14297
rect 20438 14288 20444 14300
rect 20496 14288 20502 14340
rect 16577 14263 16635 14269
rect 16577 14229 16589 14263
rect 16623 14229 16635 14263
rect 16577 14223 16635 14229
rect 17586 14220 17592 14272
rect 17644 14220 17650 14272
rect 18509 14263 18567 14269
rect 18509 14229 18521 14263
rect 18555 14260 18567 14263
rect 18690 14260 18696 14272
rect 18555 14232 18696 14260
rect 18555 14229 18567 14232
rect 18509 14223 18567 14229
rect 18690 14220 18696 14232
rect 18748 14220 18754 14272
rect 19639 14263 19697 14269
rect 19639 14229 19651 14263
rect 19685 14260 19697 14263
rect 19794 14260 19800 14272
rect 19685 14232 19800 14260
rect 19685 14229 19697 14232
rect 19639 14223 19697 14229
rect 19794 14220 19800 14232
rect 19852 14220 19858 14272
rect 1104 14170 22976 14192
rect 1104 14118 6378 14170
rect 6430 14118 6442 14170
rect 6494 14118 6506 14170
rect 6558 14118 6570 14170
rect 6622 14118 6634 14170
rect 6686 14118 11806 14170
rect 11858 14118 11870 14170
rect 11922 14118 11934 14170
rect 11986 14118 11998 14170
rect 12050 14118 12062 14170
rect 12114 14118 17234 14170
rect 17286 14118 17298 14170
rect 17350 14118 17362 14170
rect 17414 14118 17426 14170
rect 17478 14118 17490 14170
rect 17542 14118 22662 14170
rect 22714 14118 22726 14170
rect 22778 14118 22790 14170
rect 22842 14118 22854 14170
rect 22906 14118 22918 14170
rect 22970 14118 22976 14170
rect 1104 14096 22976 14118
rect 2409 14059 2467 14065
rect 2409 14025 2421 14059
rect 2455 14056 2467 14059
rect 3510 14056 3516 14068
rect 2455 14028 3516 14056
rect 2455 14025 2467 14028
rect 2409 14019 2467 14025
rect 3510 14016 3516 14028
rect 3568 14016 3574 14068
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 15473 14059 15531 14065
rect 15473 14056 15485 14059
rect 11112 14028 15485 14056
rect 11112 14016 11118 14028
rect 15473 14025 15485 14028
rect 15519 14025 15531 14059
rect 15473 14019 15531 14025
rect 15562 14016 15568 14068
rect 15620 14056 15626 14068
rect 20990 14056 20996 14068
rect 15620 14028 20996 14056
rect 15620 14016 15626 14028
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 5626 13988 5632 14000
rect 4264 13960 5632 13988
rect 2038 13880 2044 13932
rect 2096 13920 2102 13932
rect 4264 13929 4292 13960
rect 5626 13948 5632 13960
rect 5684 13948 5690 14000
rect 7650 13988 7656 14000
rect 7300 13960 7656 13988
rect 7300 13932 7328 13960
rect 7650 13948 7656 13960
rect 7708 13988 7714 14000
rect 8202 13988 8208 14000
rect 7708 13960 8208 13988
rect 7708 13948 7714 13960
rect 8202 13948 8208 13960
rect 8260 13948 8266 14000
rect 13906 13948 13912 14000
rect 13964 13988 13970 14000
rect 15746 13988 15752 14000
rect 13964 13960 15752 13988
rect 13964 13948 13970 13960
rect 15746 13948 15752 13960
rect 15804 13948 15810 14000
rect 4522 13929 4528 13932
rect 2317 13923 2375 13929
rect 2317 13920 2329 13923
rect 2096 13892 2329 13920
rect 2096 13880 2102 13892
rect 2317 13889 2329 13892
rect 2363 13889 2375 13923
rect 2317 13883 2375 13889
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 4516 13883 4528 13929
rect 4522 13880 4528 13883
rect 4580 13880 4586 13932
rect 7282 13880 7288 13932
rect 7340 13880 7346 13932
rect 10042 13929 10048 13932
rect 7541 13923 7599 13929
rect 7541 13920 7553 13923
rect 7392 13892 7553 13920
rect 6822 13812 6828 13864
rect 6880 13852 6886 13864
rect 7392 13852 7420 13892
rect 7541 13889 7553 13892
rect 7587 13889 7599 13923
rect 7541 13883 7599 13889
rect 10036 13883 10048 13929
rect 10042 13880 10048 13883
rect 10100 13880 10106 13932
rect 12796 13923 12854 13929
rect 12796 13889 12808 13923
rect 12842 13920 12854 13923
rect 12842 13892 13584 13920
rect 12842 13889 12854 13892
rect 12796 13883 12854 13889
rect 6880 13824 7420 13852
rect 6880 13812 6886 13824
rect 9766 13812 9772 13864
rect 9824 13812 9830 13864
rect 12342 13812 12348 13864
rect 12400 13852 12406 13864
rect 12529 13855 12587 13861
rect 12529 13852 12541 13855
rect 12400 13824 12541 13852
rect 12400 13812 12406 13824
rect 12529 13821 12541 13824
rect 12575 13821 12587 13855
rect 12529 13815 12587 13821
rect 13556 13784 13584 13892
rect 13630 13880 13636 13932
rect 13688 13920 13694 13932
rect 13688 13918 14044 13920
rect 13688 13892 14136 13918
rect 13688 13880 13694 13892
rect 14016 13890 14136 13892
rect 14108 13852 14136 13890
rect 14642 13880 14648 13932
rect 14700 13880 14706 13932
rect 14737 13923 14795 13929
rect 14737 13889 14749 13923
rect 14783 13889 14795 13923
rect 14737 13883 14795 13889
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13920 14979 13923
rect 15194 13920 15200 13932
rect 14967 13892 15200 13920
rect 14967 13889 14979 13892
rect 14921 13883 14979 13889
rect 14752 13852 14780 13883
rect 15194 13880 15200 13892
rect 15252 13880 15258 13932
rect 15565 13923 15623 13929
rect 15565 13920 15577 13923
rect 15304 13892 15577 13920
rect 15304 13852 15332 13892
rect 15565 13889 15577 13892
rect 15611 13889 15623 13923
rect 15565 13883 15623 13889
rect 15838 13880 15844 13932
rect 15896 13880 15902 13932
rect 16022 13880 16028 13932
rect 16080 13920 16086 13932
rect 16482 13920 16488 13932
rect 16080 13892 16488 13920
rect 16080 13880 16086 13892
rect 16482 13880 16488 13892
rect 16540 13920 16546 13932
rect 17037 13923 17095 13929
rect 17037 13920 17049 13923
rect 16540 13892 17049 13920
rect 16540 13880 16546 13892
rect 17037 13889 17049 13892
rect 17083 13889 17095 13923
rect 17037 13883 17095 13889
rect 18690 13880 18696 13932
rect 18748 13880 18754 13932
rect 19889 13923 19947 13929
rect 19889 13889 19901 13923
rect 19935 13920 19947 13923
rect 20346 13920 20352 13932
rect 19935 13892 20352 13920
rect 19935 13889 19947 13892
rect 19889 13883 19947 13889
rect 20346 13880 20352 13892
rect 20404 13880 20410 13932
rect 14108 13824 14780 13852
rect 14936 13824 15332 13852
rect 13556 13756 13860 13784
rect 5629 13719 5687 13725
rect 5629 13685 5641 13719
rect 5675 13716 5687 13719
rect 5718 13716 5724 13728
rect 5675 13688 5724 13716
rect 5675 13685 5687 13688
rect 5629 13679 5687 13685
rect 5718 13676 5724 13688
rect 5776 13676 5782 13728
rect 8662 13676 8668 13728
rect 8720 13676 8726 13728
rect 11146 13676 11152 13728
rect 11204 13676 11210 13728
rect 13832 13716 13860 13756
rect 13906 13744 13912 13796
rect 13964 13744 13970 13796
rect 14936 13793 14964 13824
rect 15378 13812 15384 13864
rect 15436 13812 15442 13864
rect 16206 13812 16212 13864
rect 16264 13812 16270 13864
rect 16666 13812 16672 13864
rect 16724 13852 16730 13864
rect 16942 13852 16948 13864
rect 16724 13824 16948 13852
rect 16724 13812 16730 13824
rect 16942 13812 16948 13824
rect 17000 13812 17006 13864
rect 18874 13812 18880 13864
rect 18932 13812 18938 13864
rect 18966 13812 18972 13864
rect 19024 13812 19030 13864
rect 19518 13812 19524 13864
rect 19576 13852 19582 13864
rect 19613 13855 19671 13861
rect 19613 13852 19625 13855
rect 19576 13824 19625 13852
rect 19576 13812 19582 13824
rect 19613 13821 19625 13824
rect 19659 13821 19671 13855
rect 19613 13815 19671 13821
rect 14921 13787 14979 13793
rect 14921 13753 14933 13787
rect 14967 13753 14979 13787
rect 14921 13747 14979 13753
rect 18509 13719 18567 13725
rect 18509 13716 18521 13719
rect 13832 13688 18521 13716
rect 18509 13685 18521 13688
rect 18555 13685 18567 13719
rect 18509 13679 18567 13685
rect 1104 13626 22816 13648
rect 1104 13574 3664 13626
rect 3716 13574 3728 13626
rect 3780 13574 3792 13626
rect 3844 13574 3856 13626
rect 3908 13574 3920 13626
rect 3972 13574 9092 13626
rect 9144 13574 9156 13626
rect 9208 13574 9220 13626
rect 9272 13574 9284 13626
rect 9336 13574 9348 13626
rect 9400 13574 14520 13626
rect 14572 13574 14584 13626
rect 14636 13574 14648 13626
rect 14700 13574 14712 13626
rect 14764 13574 14776 13626
rect 14828 13574 19948 13626
rect 20000 13574 20012 13626
rect 20064 13574 20076 13626
rect 20128 13574 20140 13626
rect 20192 13574 20204 13626
rect 20256 13574 22816 13626
rect 1104 13552 22816 13574
rect 5626 13472 5632 13524
rect 5684 13512 5690 13524
rect 5721 13515 5779 13521
rect 5721 13512 5733 13515
rect 5684 13484 5733 13512
rect 5684 13472 5690 13484
rect 5721 13481 5733 13484
rect 5767 13512 5779 13515
rect 7282 13512 7288 13524
rect 5767 13484 7288 13512
rect 5767 13481 5779 13484
rect 5721 13475 5779 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 19702 13404 19708 13456
rect 19760 13404 19766 13456
rect 16758 13376 16764 13388
rect 16408 13348 16764 13376
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13308 7067 13311
rect 10413 13311 10471 13317
rect 10413 13308 10425 13311
rect 7055 13280 10425 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 10413 13277 10425 13280
rect 10459 13308 10471 13311
rect 10594 13308 10600 13320
rect 10459 13280 10600 13308
rect 10459 13277 10471 13280
rect 10413 13271 10471 13277
rect 10594 13268 10600 13280
rect 10652 13268 10658 13320
rect 16408 13317 16436 13348
rect 16758 13336 16764 13348
rect 16816 13376 16822 13388
rect 18233 13379 18291 13385
rect 18233 13376 18245 13379
rect 16816 13348 18245 13376
rect 16816 13336 16822 13348
rect 18233 13345 18245 13348
rect 18279 13345 18291 13379
rect 18233 13339 18291 13345
rect 19426 13336 19432 13388
rect 19484 13376 19490 13388
rect 19886 13376 19892 13388
rect 19484 13348 19892 13376
rect 19484 13336 19490 13348
rect 19886 13336 19892 13348
rect 19944 13376 19950 13388
rect 19981 13379 20039 13385
rect 19981 13376 19993 13379
rect 19944 13348 19993 13376
rect 19944 13336 19950 13348
rect 19981 13345 19993 13348
rect 20027 13345 20039 13379
rect 19981 13339 20039 13345
rect 16393 13311 16451 13317
rect 16393 13277 16405 13311
rect 16439 13277 16451 13311
rect 16393 13271 16451 13277
rect 16485 13311 16543 13317
rect 16485 13277 16497 13311
rect 16531 13308 16543 13311
rect 16942 13308 16948 13320
rect 16531 13280 16948 13308
rect 16531 13277 16543 13280
rect 16485 13271 16543 13277
rect 16942 13268 16948 13280
rect 17000 13268 17006 13320
rect 18046 13268 18052 13320
rect 18104 13268 18110 13320
rect 18601 13311 18659 13317
rect 18601 13277 18613 13311
rect 18647 13308 18659 13311
rect 18966 13308 18972 13320
rect 18647 13280 18972 13308
rect 18647 13277 18659 13280
rect 18601 13271 18659 13277
rect 18966 13268 18972 13280
rect 19024 13268 19030 13320
rect 12161 13243 12219 13249
rect 12161 13209 12173 13243
rect 12207 13240 12219 13243
rect 12342 13240 12348 13252
rect 12207 13212 12348 13240
rect 12207 13209 12219 13212
rect 12161 13203 12219 13209
rect 12342 13200 12348 13212
rect 12400 13200 12406 13252
rect 16761 13243 16819 13249
rect 16761 13209 16773 13243
rect 16807 13240 16819 13243
rect 16850 13240 16856 13252
rect 16807 13212 16856 13240
rect 16807 13209 16819 13212
rect 16761 13203 16819 13209
rect 16850 13200 16856 13212
rect 16908 13200 16914 13252
rect 18785 13243 18843 13249
rect 18785 13209 18797 13243
rect 18831 13240 18843 13243
rect 19242 13240 19248 13252
rect 18831 13212 19248 13240
rect 18831 13209 18843 13212
rect 18785 13203 18843 13209
rect 19242 13200 19248 13212
rect 19300 13200 19306 13252
rect 16206 13132 16212 13184
rect 16264 13132 16270 13184
rect 16574 13132 16580 13184
rect 16632 13132 16638 13184
rect 18690 13132 18696 13184
rect 18748 13132 18754 13184
rect 18966 13132 18972 13184
rect 19024 13172 19030 13184
rect 19521 13175 19579 13181
rect 19521 13172 19533 13175
rect 19024 13144 19533 13172
rect 19024 13132 19030 13144
rect 19521 13141 19533 13144
rect 19567 13141 19579 13175
rect 19521 13135 19579 13141
rect 1104 13082 22976 13104
rect 1104 13030 6378 13082
rect 6430 13030 6442 13082
rect 6494 13030 6506 13082
rect 6558 13030 6570 13082
rect 6622 13030 6634 13082
rect 6686 13030 11806 13082
rect 11858 13030 11870 13082
rect 11922 13030 11934 13082
rect 11986 13030 11998 13082
rect 12050 13030 12062 13082
rect 12114 13030 17234 13082
rect 17286 13030 17298 13082
rect 17350 13030 17362 13082
rect 17414 13030 17426 13082
rect 17478 13030 17490 13082
rect 17542 13030 22662 13082
rect 22714 13030 22726 13082
rect 22778 13030 22790 13082
rect 22842 13030 22854 13082
rect 22906 13030 22918 13082
rect 22970 13030 22976 13082
rect 1104 13008 22976 13030
rect 16025 12971 16083 12977
rect 16025 12937 16037 12971
rect 16071 12937 16083 12971
rect 16025 12931 16083 12937
rect 8196 12903 8254 12909
rect 8196 12869 8208 12903
rect 8242 12900 8254 12903
rect 8294 12900 8300 12912
rect 8242 12872 8300 12900
rect 8242 12869 8254 12872
rect 8196 12863 8254 12869
rect 8294 12860 8300 12872
rect 8352 12860 8358 12912
rect 12888 12903 12946 12909
rect 12888 12869 12900 12903
rect 12934 12900 12946 12903
rect 16040 12900 16068 12931
rect 19886 12928 19892 12980
rect 19944 12928 19950 12980
rect 12934 12872 16068 12900
rect 12934 12869 12946 12872
rect 12888 12863 12946 12869
rect 19058 12860 19064 12912
rect 19116 12900 19122 12912
rect 19518 12900 19524 12912
rect 19116 12872 19524 12900
rect 19116 12860 19122 12872
rect 19518 12860 19524 12872
rect 19576 12900 19582 12912
rect 19797 12903 19855 12909
rect 19797 12900 19809 12903
rect 19576 12872 19809 12900
rect 19576 12860 19582 12872
rect 19797 12869 19809 12872
rect 19843 12869 19855 12903
rect 19797 12863 19855 12869
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 5270 12835 5328 12841
rect 5270 12832 5282 12835
rect 4304 12804 5282 12832
rect 4304 12792 4310 12804
rect 5270 12801 5282 12804
rect 5316 12801 5328 12835
rect 5270 12795 5328 12801
rect 5537 12835 5595 12841
rect 5537 12801 5549 12835
rect 5583 12832 5595 12835
rect 5626 12832 5632 12844
rect 5583 12804 5632 12832
rect 5583 12801 5595 12804
rect 5537 12795 5595 12801
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 10036 12835 10094 12841
rect 10036 12801 10048 12835
rect 10082 12832 10094 12835
rect 11606 12832 11612 12844
rect 10082 12804 11612 12832
rect 10082 12801 10094 12804
rect 10036 12795 10094 12801
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 15194 12792 15200 12844
rect 15252 12832 15258 12844
rect 16025 12835 16083 12841
rect 16025 12832 16037 12835
rect 15252 12804 16037 12832
rect 15252 12792 15258 12804
rect 16025 12801 16037 12804
rect 16071 12832 16083 12835
rect 16206 12832 16212 12844
rect 16071 12804 16212 12832
rect 16071 12801 16083 12804
rect 16025 12795 16083 12801
rect 16206 12792 16212 12804
rect 16264 12792 16270 12844
rect 19245 12835 19303 12841
rect 19245 12801 19257 12835
rect 19291 12832 19303 12835
rect 19610 12832 19616 12844
rect 19291 12804 19616 12832
rect 19291 12801 19303 12804
rect 19245 12795 19303 12801
rect 19610 12792 19616 12804
rect 19668 12792 19674 12844
rect 7929 12767 7987 12773
rect 7929 12733 7941 12767
rect 7975 12733 7987 12767
rect 7929 12727 7987 12733
rect 4157 12631 4215 12637
rect 4157 12597 4169 12631
rect 4203 12628 4215 12631
rect 4430 12628 4436 12640
rect 4203 12600 4436 12628
rect 4203 12597 4215 12600
rect 4157 12591 4215 12597
rect 4430 12588 4436 12600
rect 4488 12588 4494 12640
rect 7944 12628 7972 12727
rect 9766 12724 9772 12776
rect 9824 12724 9830 12776
rect 12342 12724 12348 12776
rect 12400 12764 12406 12776
rect 12621 12767 12679 12773
rect 12621 12764 12633 12767
rect 12400 12736 12633 12764
rect 12400 12724 12406 12736
rect 12621 12733 12633 12736
rect 12667 12733 12679 12767
rect 12621 12727 12679 12733
rect 15378 12724 15384 12776
rect 15436 12764 15442 12776
rect 15749 12767 15807 12773
rect 15749 12764 15761 12767
rect 15436 12736 15761 12764
rect 15436 12724 15442 12736
rect 15749 12733 15761 12736
rect 15795 12733 15807 12767
rect 15749 12727 15807 12733
rect 18598 12724 18604 12776
rect 18656 12764 18662 12776
rect 18877 12767 18935 12773
rect 18877 12764 18889 12767
rect 18656 12736 18889 12764
rect 18656 12724 18662 12736
rect 18877 12733 18889 12736
rect 18923 12733 18935 12767
rect 18877 12727 18935 12733
rect 8202 12628 8208 12640
rect 7944 12600 8208 12628
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 9309 12631 9367 12637
rect 9309 12597 9321 12631
rect 9355 12628 9367 12631
rect 9582 12628 9588 12640
rect 9355 12600 9588 12628
rect 9355 12597 9367 12600
rect 9309 12591 9367 12597
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 9784 12628 9812 12724
rect 15933 12699 15991 12705
rect 15933 12665 15945 12699
rect 15979 12696 15991 12699
rect 16850 12696 16856 12708
rect 15979 12668 16856 12696
rect 15979 12665 15991 12668
rect 15933 12659 15991 12665
rect 16850 12656 16856 12668
rect 16908 12656 16914 12708
rect 18506 12656 18512 12708
rect 18564 12696 18570 12708
rect 19080 12699 19138 12705
rect 19080 12696 19092 12699
rect 18564 12668 19092 12696
rect 18564 12656 18570 12668
rect 19080 12665 19092 12668
rect 19126 12665 19138 12699
rect 19080 12659 19138 12665
rect 11054 12628 11060 12640
rect 9784 12600 11060 12628
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 11149 12631 11207 12637
rect 11149 12597 11161 12631
rect 11195 12628 11207 12631
rect 13262 12628 13268 12640
rect 11195 12600 13268 12628
rect 11195 12597 11207 12600
rect 11149 12591 11207 12597
rect 13262 12588 13268 12600
rect 13320 12588 13326 12640
rect 14001 12631 14059 12637
rect 14001 12597 14013 12631
rect 14047 12628 14059 12631
rect 16574 12628 16580 12640
rect 14047 12600 16580 12628
rect 14047 12597 14059 12600
rect 14001 12591 14059 12597
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 18138 12588 18144 12640
rect 18196 12628 18202 12640
rect 18601 12631 18659 12637
rect 18601 12628 18613 12631
rect 18196 12600 18613 12628
rect 18196 12588 18202 12600
rect 18601 12597 18613 12600
rect 18647 12628 18659 12631
rect 18690 12628 18696 12640
rect 18647 12600 18696 12628
rect 18647 12597 18659 12600
rect 18601 12591 18659 12597
rect 18690 12588 18696 12600
rect 18748 12588 18754 12640
rect 18966 12588 18972 12640
rect 19024 12588 19030 12640
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 19886 12628 19892 12640
rect 19392 12600 19892 12628
rect 19392 12588 19398 12600
rect 19886 12588 19892 12600
rect 19944 12588 19950 12640
rect 1104 12538 22816 12560
rect 1104 12486 3664 12538
rect 3716 12486 3728 12538
rect 3780 12486 3792 12538
rect 3844 12486 3856 12538
rect 3908 12486 3920 12538
rect 3972 12486 9092 12538
rect 9144 12486 9156 12538
rect 9208 12486 9220 12538
rect 9272 12486 9284 12538
rect 9336 12486 9348 12538
rect 9400 12486 14520 12538
rect 14572 12486 14584 12538
rect 14636 12486 14648 12538
rect 14700 12486 14712 12538
rect 14764 12486 14776 12538
rect 14828 12486 19948 12538
rect 20000 12486 20012 12538
rect 20064 12486 20076 12538
rect 20128 12486 20140 12538
rect 20192 12486 20204 12538
rect 20256 12486 22816 12538
rect 1104 12464 22816 12486
rect 5718 12384 5724 12436
rect 5776 12424 5782 12436
rect 6178 12424 6184 12436
rect 5776 12396 6184 12424
rect 5776 12384 5782 12396
rect 6178 12384 6184 12396
rect 6236 12384 6242 12436
rect 15286 12384 15292 12436
rect 15344 12424 15350 12436
rect 15657 12427 15715 12433
rect 15657 12424 15669 12427
rect 15344 12396 15669 12424
rect 15344 12384 15350 12396
rect 15657 12393 15669 12396
rect 15703 12424 15715 12427
rect 15703 12396 19472 12424
rect 15703 12393 15715 12396
rect 15657 12387 15715 12393
rect 15838 12316 15844 12368
rect 15896 12356 15902 12368
rect 16209 12359 16267 12365
rect 16209 12356 16221 12359
rect 15896 12328 16221 12356
rect 15896 12316 15902 12328
rect 16209 12325 16221 12328
rect 16255 12325 16267 12359
rect 16209 12319 16267 12325
rect 16942 12316 16948 12368
rect 17000 12356 17006 12368
rect 17000 12328 19334 12356
rect 17000 12316 17006 12328
rect 3142 12288 3148 12300
rect 2516 12260 3148 12288
rect 1946 12180 1952 12232
rect 2004 12220 2010 12232
rect 2222 12220 2228 12232
rect 2004 12192 2228 12220
rect 2004 12180 2010 12192
rect 2222 12180 2228 12192
rect 2280 12180 2286 12232
rect 2516 12229 2544 12260
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 11054 12248 11060 12300
rect 11112 12288 11118 12300
rect 11333 12291 11391 12297
rect 11333 12288 11345 12291
rect 11112 12260 11345 12288
rect 11112 12248 11118 12260
rect 11333 12257 11345 12260
rect 11379 12257 11391 12291
rect 11333 12251 11391 12257
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12189 2467 12223
rect 2409 12183 2467 12189
rect 2501 12223 2559 12229
rect 2501 12189 2513 12223
rect 2547 12189 2559 12223
rect 2501 12183 2559 12189
rect 2424 12152 2452 12183
rect 2590 12180 2596 12232
rect 2648 12180 2654 12232
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 6365 12223 6423 12229
rect 6365 12220 6377 12223
rect 5684 12192 6377 12220
rect 5684 12180 5690 12192
rect 6365 12189 6377 12192
rect 6411 12189 6423 12223
rect 6365 12183 6423 12189
rect 8202 12180 8208 12232
rect 8260 12220 8266 12232
rect 9217 12223 9275 12229
rect 9217 12220 9229 12223
rect 8260 12192 9229 12220
rect 8260 12180 8266 12192
rect 9217 12189 9229 12192
rect 9263 12189 9275 12223
rect 9217 12183 9275 12189
rect 9493 12223 9551 12229
rect 9493 12189 9505 12223
rect 9539 12220 9551 12223
rect 10318 12220 10324 12232
rect 9539 12192 10324 12220
rect 9539 12189 9551 12192
rect 9493 12183 9551 12189
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 11348 12220 11376 12251
rect 15654 12248 15660 12300
rect 15712 12288 15718 12300
rect 15712 12260 16436 12288
rect 15712 12248 15718 12260
rect 12342 12220 12348 12232
rect 11348 12192 12348 12220
rect 12342 12180 12348 12192
rect 12400 12220 12406 12232
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 12400 12192 14289 12220
rect 12400 12180 12406 12192
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 16114 12180 16120 12232
rect 16172 12180 16178 12232
rect 16408 12229 16436 12260
rect 16574 12248 16580 12300
rect 16632 12288 16638 12300
rect 17862 12288 17868 12300
rect 16632 12260 17868 12288
rect 16632 12248 16638 12260
rect 17862 12248 17868 12260
rect 17920 12288 17926 12300
rect 17920 12260 18276 12288
rect 17920 12248 17926 12260
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12189 16451 12223
rect 18141 12223 18199 12229
rect 18141 12220 18153 12223
rect 16393 12183 16451 12189
rect 16500 12192 18153 12220
rect 2774 12152 2780 12164
rect 2424 12124 2780 12152
rect 2774 12112 2780 12124
rect 2832 12112 2838 12164
rect 2869 12155 2927 12161
rect 2869 12121 2881 12155
rect 2915 12152 2927 12155
rect 5362 12155 5420 12161
rect 5362 12152 5374 12155
rect 2915 12124 5374 12152
rect 2915 12121 2927 12124
rect 2869 12115 2927 12121
rect 5362 12121 5374 12124
rect 5408 12121 5420 12155
rect 5362 12115 5420 12121
rect 6632 12155 6690 12161
rect 6632 12121 6644 12155
rect 6678 12152 6690 12155
rect 6730 12152 6736 12164
rect 6678 12124 6736 12152
rect 6678 12121 6690 12124
rect 6632 12115 6690 12121
rect 6730 12112 6736 12124
rect 6788 12112 6794 12164
rect 11238 12112 11244 12164
rect 11296 12152 11302 12164
rect 11578 12155 11636 12161
rect 11578 12152 11590 12155
rect 11296 12124 11590 12152
rect 11296 12112 11302 12124
rect 11578 12121 11590 12124
rect 11624 12121 11636 12155
rect 11578 12115 11636 12121
rect 13906 12112 13912 12164
rect 13964 12152 13970 12164
rect 14522 12155 14580 12161
rect 14522 12152 14534 12155
rect 13964 12124 14534 12152
rect 13964 12112 13970 12124
rect 14522 12121 14534 12124
rect 14568 12121 14580 12155
rect 14522 12115 14580 12121
rect 4154 12044 4160 12096
rect 4212 12084 4218 12096
rect 4249 12087 4307 12093
rect 4249 12084 4261 12087
rect 4212 12056 4261 12084
rect 4212 12044 4218 12056
rect 4249 12053 4261 12056
rect 4295 12053 4307 12087
rect 4249 12047 4307 12053
rect 7374 12044 7380 12096
rect 7432 12084 7438 12096
rect 7745 12087 7803 12093
rect 7745 12084 7757 12087
rect 7432 12056 7757 12084
rect 7432 12044 7438 12056
rect 7745 12053 7757 12056
rect 7791 12053 7803 12087
rect 7745 12047 7803 12053
rect 10502 12044 10508 12096
rect 10560 12084 10566 12096
rect 10597 12087 10655 12093
rect 10597 12084 10609 12087
rect 10560 12056 10609 12084
rect 10560 12044 10566 12056
rect 10597 12053 10609 12056
rect 10643 12053 10655 12087
rect 10597 12047 10655 12053
rect 12713 12087 12771 12093
rect 12713 12053 12725 12087
rect 12759 12084 12771 12087
rect 13630 12084 13636 12096
rect 12759 12056 13636 12084
rect 12759 12053 12771 12056
rect 12713 12047 12771 12053
rect 13630 12044 13636 12056
rect 13688 12084 13694 12096
rect 16500 12084 16528 12192
rect 18141 12189 18153 12192
rect 18187 12189 18199 12223
rect 18248 12220 18276 12260
rect 18322 12248 18328 12300
rect 18380 12288 18386 12300
rect 18601 12291 18659 12297
rect 18601 12288 18613 12291
rect 18380 12260 18613 12288
rect 18380 12248 18386 12260
rect 18601 12257 18613 12260
rect 18647 12257 18659 12291
rect 18601 12251 18659 12257
rect 18693 12223 18751 12229
rect 18693 12220 18705 12223
rect 18248 12192 18705 12220
rect 18141 12183 18199 12189
rect 18693 12189 18705 12192
rect 18739 12189 18751 12223
rect 19306 12220 19334 12328
rect 19444 12297 19472 12396
rect 19429 12291 19487 12297
rect 19429 12257 19441 12291
rect 19475 12257 19487 12291
rect 19429 12251 19487 12257
rect 19610 12248 19616 12300
rect 19668 12248 19674 12300
rect 19886 12248 19892 12300
rect 19944 12248 19950 12300
rect 19981 12223 20039 12229
rect 19981 12220 19993 12223
rect 19306 12192 19993 12220
rect 18693 12183 18751 12189
rect 19444 12164 19472 12192
rect 19981 12189 19993 12192
rect 20027 12189 20039 12223
rect 19981 12183 20039 12189
rect 16853 12155 16911 12161
rect 16853 12121 16865 12155
rect 16899 12152 16911 12155
rect 18230 12152 18236 12164
rect 16899 12124 18236 12152
rect 16899 12121 16911 12124
rect 16853 12115 16911 12121
rect 18230 12112 18236 12124
rect 18288 12152 18294 12164
rect 18598 12152 18604 12164
rect 18288 12124 18604 12152
rect 18288 12112 18294 12124
rect 18598 12112 18604 12124
rect 18656 12112 18662 12164
rect 19426 12112 19432 12164
rect 19484 12112 19490 12164
rect 13688 12056 16528 12084
rect 18325 12087 18383 12093
rect 13688 12044 13694 12056
rect 18325 12053 18337 12087
rect 18371 12084 18383 12087
rect 18506 12084 18512 12096
rect 18371 12056 18512 12084
rect 18371 12053 18383 12056
rect 18325 12047 18383 12053
rect 18506 12044 18512 12056
rect 18564 12084 18570 12096
rect 19150 12084 19156 12096
rect 18564 12056 19156 12084
rect 18564 12044 18570 12056
rect 19150 12044 19156 12056
rect 19208 12044 19214 12096
rect 19334 12044 19340 12096
rect 19392 12084 19398 12096
rect 19886 12084 19892 12096
rect 19392 12056 19892 12084
rect 19392 12044 19398 12056
rect 19886 12044 19892 12056
rect 19944 12044 19950 12096
rect 1104 11994 22976 12016
rect 1104 11942 6378 11994
rect 6430 11942 6442 11994
rect 6494 11942 6506 11994
rect 6558 11942 6570 11994
rect 6622 11942 6634 11994
rect 6686 11942 11806 11994
rect 11858 11942 11870 11994
rect 11922 11942 11934 11994
rect 11986 11942 11998 11994
rect 12050 11942 12062 11994
rect 12114 11942 17234 11994
rect 17286 11942 17298 11994
rect 17350 11942 17362 11994
rect 17414 11942 17426 11994
rect 17478 11942 17490 11994
rect 17542 11942 22662 11994
rect 22714 11942 22726 11994
rect 22778 11942 22790 11994
rect 22842 11942 22854 11994
rect 22906 11942 22918 11994
rect 22970 11942 22976 11994
rect 1104 11920 22976 11942
rect 2501 11883 2559 11889
rect 2501 11849 2513 11883
rect 2547 11880 2559 11883
rect 2590 11880 2596 11892
rect 2547 11852 2596 11880
rect 2547 11849 2559 11852
rect 2501 11843 2559 11849
rect 2590 11840 2596 11852
rect 2648 11840 2654 11892
rect 2774 11840 2780 11892
rect 2832 11880 2838 11892
rect 2961 11883 3019 11889
rect 2961 11880 2973 11883
rect 2832 11852 2973 11880
rect 2832 11840 2838 11852
rect 2961 11849 2973 11852
rect 3007 11849 3019 11883
rect 2961 11843 3019 11849
rect 16850 11840 16856 11892
rect 16908 11840 16914 11892
rect 18322 11840 18328 11892
rect 18380 11880 18386 11892
rect 19334 11880 19340 11892
rect 18380 11852 19340 11880
rect 18380 11840 18386 11852
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 19518 11840 19524 11892
rect 19576 11840 19582 11892
rect 4154 11812 4160 11824
rect 2976 11784 4160 11812
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11744 2375 11747
rect 2682 11744 2688 11756
rect 2363 11716 2688 11744
rect 2363 11713 2375 11716
rect 2317 11707 2375 11713
rect 2682 11704 2688 11716
rect 2740 11744 2746 11756
rect 2976 11753 3004 11784
rect 4154 11772 4160 11784
rect 4212 11772 4218 11824
rect 5626 11812 5632 11824
rect 4264 11784 5632 11812
rect 2961 11747 3019 11753
rect 2961 11744 2973 11747
rect 2740 11716 2973 11744
rect 2740 11704 2746 11716
rect 2961 11713 2973 11716
rect 3007 11713 3019 11747
rect 2961 11707 3019 11713
rect 3142 11704 3148 11756
rect 3200 11704 3206 11756
rect 4264 11753 4292 11784
rect 5626 11772 5632 11784
rect 5684 11772 5690 11824
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11713 4307 11747
rect 4505 11747 4563 11753
rect 4505 11744 4517 11747
rect 4249 11707 4307 11713
rect 4356 11716 4517 11744
rect 2133 11679 2191 11685
rect 2133 11645 2145 11679
rect 2179 11676 2191 11679
rect 2590 11676 2596 11688
rect 2179 11648 2596 11676
rect 2179 11645 2191 11648
rect 2133 11639 2191 11645
rect 2590 11636 2596 11648
rect 2648 11636 2654 11688
rect 4154 11636 4160 11688
rect 4212 11676 4218 11688
rect 4356 11676 4384 11716
rect 4505 11713 4517 11716
rect 4551 11713 4563 11747
rect 4505 11707 4563 11713
rect 8202 11704 8208 11756
rect 8260 11744 8266 11756
rect 8570 11753 8576 11756
rect 8297 11747 8355 11753
rect 8297 11744 8309 11747
rect 8260 11716 8309 11744
rect 8260 11704 8266 11716
rect 8297 11713 8309 11716
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 8564 11707 8576 11753
rect 8570 11704 8576 11707
rect 8628 11704 8634 11756
rect 12342 11704 12348 11756
rect 12400 11744 12406 11756
rect 12621 11747 12679 11753
rect 12621 11744 12633 11747
rect 12400 11716 12633 11744
rect 12400 11704 12406 11716
rect 12621 11713 12633 11716
rect 12667 11713 12679 11747
rect 12621 11707 12679 11713
rect 12888 11747 12946 11753
rect 12888 11713 12900 11747
rect 12934 11744 12946 11747
rect 13170 11744 13176 11756
rect 12934 11716 13176 11744
rect 12934 11713 12946 11716
rect 12888 11707 12946 11713
rect 13170 11704 13176 11716
rect 13228 11704 13234 11756
rect 15654 11704 15660 11756
rect 15712 11704 15718 11756
rect 16117 11747 16175 11753
rect 16117 11713 16129 11747
rect 16163 11713 16175 11747
rect 16117 11707 16175 11713
rect 4212 11648 4384 11676
rect 4212 11636 4218 11648
rect 15194 11636 15200 11688
rect 15252 11676 15258 11688
rect 16132 11676 16160 11707
rect 17034 11704 17040 11756
rect 17092 11704 17098 11756
rect 17221 11747 17279 11753
rect 17221 11713 17233 11747
rect 17267 11744 17279 11747
rect 17586 11744 17592 11756
rect 17267 11716 17592 11744
rect 17267 11713 17279 11716
rect 17221 11707 17279 11713
rect 17586 11704 17592 11716
rect 17644 11704 17650 11756
rect 18230 11704 18236 11756
rect 18288 11744 18294 11756
rect 18325 11747 18383 11753
rect 18325 11744 18337 11747
rect 18288 11716 18337 11744
rect 18288 11704 18294 11716
rect 18325 11713 18337 11716
rect 18371 11713 18383 11747
rect 18325 11707 18383 11713
rect 18966 11704 18972 11756
rect 19024 11704 19030 11756
rect 19150 11704 19156 11756
rect 19208 11704 19214 11756
rect 19610 11704 19616 11756
rect 19668 11704 19674 11756
rect 15252 11648 16160 11676
rect 17313 11679 17371 11685
rect 15252 11636 15258 11648
rect 17313 11645 17325 11679
rect 17359 11645 17371 11679
rect 17313 11639 17371 11645
rect 15470 11568 15476 11620
rect 15528 11608 15534 11620
rect 15749 11611 15807 11617
rect 15749 11608 15761 11611
rect 15528 11580 15761 11608
rect 15528 11568 15534 11580
rect 15749 11577 15761 11580
rect 15795 11608 15807 11611
rect 16482 11608 16488 11620
rect 15795 11580 16488 11608
rect 15795 11577 15807 11580
rect 15749 11571 15807 11577
rect 16482 11568 16488 11580
rect 16540 11608 16546 11620
rect 17328 11608 17356 11639
rect 16540 11580 17356 11608
rect 16540 11568 16546 11580
rect 5629 11543 5687 11549
rect 5629 11509 5641 11543
rect 5675 11540 5687 11543
rect 5994 11540 6000 11552
rect 5675 11512 6000 11540
rect 5675 11509 5687 11512
rect 5629 11503 5687 11509
rect 5994 11500 6000 11512
rect 6052 11500 6058 11552
rect 9674 11500 9680 11552
rect 9732 11500 9738 11552
rect 14001 11543 14059 11549
rect 14001 11509 14013 11543
rect 14047 11540 14059 11543
rect 15562 11540 15568 11552
rect 14047 11512 15568 11540
rect 14047 11509 14059 11512
rect 14001 11503 14059 11509
rect 15562 11500 15568 11512
rect 15620 11500 15626 11552
rect 1104 11450 22816 11472
rect 1104 11398 3664 11450
rect 3716 11398 3728 11450
rect 3780 11398 3792 11450
rect 3844 11398 3856 11450
rect 3908 11398 3920 11450
rect 3972 11398 9092 11450
rect 9144 11398 9156 11450
rect 9208 11398 9220 11450
rect 9272 11398 9284 11450
rect 9336 11398 9348 11450
rect 9400 11398 14520 11450
rect 14572 11398 14584 11450
rect 14636 11398 14648 11450
rect 14700 11398 14712 11450
rect 14764 11398 14776 11450
rect 14828 11398 19948 11450
rect 20000 11398 20012 11450
rect 20064 11398 20076 11450
rect 20128 11398 20140 11450
rect 20192 11398 20204 11450
rect 20256 11398 22816 11450
rect 1104 11376 22816 11398
rect 7466 11228 7472 11280
rect 7524 11268 7530 11280
rect 7653 11271 7711 11277
rect 7653 11268 7665 11271
rect 7524 11240 7665 11268
rect 7524 11228 7530 11240
rect 7653 11237 7665 11240
rect 7699 11237 7711 11271
rect 7653 11231 7711 11237
rect 15562 11228 15568 11280
rect 15620 11268 15626 11280
rect 16025 11271 16083 11277
rect 16025 11268 16037 11271
rect 15620 11240 16037 11268
rect 15620 11228 15626 11240
rect 16025 11237 16037 11240
rect 16071 11268 16083 11271
rect 16298 11268 16304 11280
rect 16071 11240 16304 11268
rect 16071 11237 16083 11240
rect 16025 11231 16083 11237
rect 16298 11228 16304 11240
rect 16356 11228 16362 11280
rect 5626 11160 5632 11212
rect 5684 11200 5690 11212
rect 6273 11203 6331 11209
rect 6273 11200 6285 11203
rect 5684 11172 6285 11200
rect 5684 11160 5690 11172
rect 6273 11169 6285 11172
rect 6319 11169 6331 11203
rect 6273 11163 6331 11169
rect 15654 11160 15660 11212
rect 15712 11200 15718 11212
rect 15749 11203 15807 11209
rect 15749 11200 15761 11203
rect 15712 11172 15761 11200
rect 15712 11160 15718 11172
rect 15749 11169 15761 11172
rect 15795 11169 15807 11203
rect 15749 11163 15807 11169
rect 16209 11203 16267 11209
rect 16209 11169 16221 11203
rect 16255 11200 16267 11203
rect 18598 11200 18604 11212
rect 16255 11172 18604 11200
rect 16255 11169 16267 11172
rect 16209 11163 16267 11169
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 17862 11092 17868 11144
rect 17920 11132 17926 11144
rect 18171 11135 18229 11141
rect 18171 11132 18183 11135
rect 17920 11104 18183 11132
rect 17920 11092 17926 11104
rect 18171 11101 18183 11104
rect 18217 11101 18229 11135
rect 18171 11095 18229 11101
rect 18322 11092 18328 11144
rect 18380 11092 18386 11144
rect 5902 11024 5908 11076
rect 5960 11064 5966 11076
rect 6518 11067 6576 11073
rect 6518 11064 6530 11067
rect 5960 11036 6530 11064
rect 5960 11024 5966 11036
rect 6518 11033 6530 11036
rect 6564 11033 6576 11067
rect 6518 11027 6576 11033
rect 17034 11024 17040 11076
rect 17092 11064 17098 11076
rect 17957 11067 18015 11073
rect 17957 11064 17969 11067
rect 17092 11036 17969 11064
rect 17092 11024 17098 11036
rect 17957 11033 17969 11036
rect 18003 11033 18015 11067
rect 17957 11027 18015 11033
rect 1104 10906 22976 10928
rect 1104 10854 6378 10906
rect 6430 10854 6442 10906
rect 6494 10854 6506 10906
rect 6558 10854 6570 10906
rect 6622 10854 6634 10906
rect 6686 10854 11806 10906
rect 11858 10854 11870 10906
rect 11922 10854 11934 10906
rect 11986 10854 11998 10906
rect 12050 10854 12062 10906
rect 12114 10854 17234 10906
rect 17286 10854 17298 10906
rect 17350 10854 17362 10906
rect 17414 10854 17426 10906
rect 17478 10854 17490 10906
rect 17542 10854 22662 10906
rect 22714 10854 22726 10906
rect 22778 10854 22790 10906
rect 22842 10854 22854 10906
rect 22906 10854 22918 10906
rect 22970 10854 22976 10906
rect 1104 10832 22976 10854
rect 2133 10795 2191 10801
rect 2133 10761 2145 10795
rect 2179 10761 2191 10795
rect 2133 10755 2191 10761
rect 1857 10727 1915 10733
rect 1857 10693 1869 10727
rect 1903 10724 1915 10727
rect 2038 10724 2044 10736
rect 1903 10696 2044 10724
rect 1903 10693 1915 10696
rect 1857 10687 1915 10693
rect 2038 10684 2044 10696
rect 2096 10684 2102 10736
rect 2148 10724 2176 10755
rect 2590 10752 2596 10804
rect 2648 10792 2654 10804
rect 2961 10795 3019 10801
rect 2961 10792 2973 10795
rect 2648 10764 2973 10792
rect 2648 10752 2654 10764
rect 2961 10761 2973 10764
rect 3007 10761 3019 10795
rect 2961 10755 3019 10761
rect 3513 10795 3571 10801
rect 3513 10761 3525 10795
rect 3559 10792 3571 10795
rect 4338 10792 4344 10804
rect 3559 10764 4344 10792
rect 3559 10761 3571 10764
rect 3513 10755 3571 10761
rect 4338 10752 4344 10764
rect 4396 10752 4402 10804
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 6638 10792 6644 10804
rect 5684 10764 6644 10792
rect 5684 10752 5690 10764
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 8389 10795 8447 10801
rect 8389 10792 8401 10795
rect 8352 10764 8401 10792
rect 8352 10752 8358 10764
rect 8389 10761 8401 10764
rect 8435 10761 8447 10795
rect 8389 10755 8447 10761
rect 13357 10795 13415 10801
rect 13357 10761 13369 10795
rect 13403 10792 13415 10795
rect 13906 10792 13912 10804
rect 13403 10764 13912 10792
rect 13403 10761 13415 10764
rect 13357 10755 13415 10761
rect 13906 10752 13912 10764
rect 13964 10752 13970 10804
rect 4154 10724 4160 10736
rect 2148 10696 4160 10724
rect 4154 10684 4160 10696
rect 4212 10684 4218 10736
rect 7285 10727 7343 10733
rect 7285 10724 7297 10727
rect 5736 10696 6500 10724
rect 2056 10588 2084 10684
rect 2133 10659 2191 10665
rect 2133 10625 2145 10659
rect 2179 10656 2191 10659
rect 2314 10656 2320 10668
rect 2179 10628 2320 10656
rect 2179 10625 2191 10628
rect 2133 10619 2191 10625
rect 2314 10616 2320 10628
rect 2372 10656 2378 10668
rect 2777 10659 2835 10665
rect 2777 10656 2789 10659
rect 2372 10628 2789 10656
rect 2372 10616 2378 10628
rect 2777 10625 2789 10628
rect 2823 10625 2835 10659
rect 2777 10619 2835 10625
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10625 3111 10659
rect 3053 10619 3111 10625
rect 3068 10588 3096 10619
rect 3510 10616 3516 10668
rect 3568 10616 3574 10668
rect 4430 10656 4436 10668
rect 3620 10628 4436 10656
rect 3620 10588 3648 10628
rect 4430 10616 4436 10628
rect 4488 10616 4494 10668
rect 5736 10665 5764 10696
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 5828 10628 6408 10656
rect 3789 10591 3847 10597
rect 3789 10588 3801 10591
rect 2056 10560 2728 10588
rect 3068 10560 3648 10588
rect 3712 10560 3801 10588
rect 2038 10480 2044 10532
rect 2096 10480 2102 10532
rect 2700 10452 2728 10560
rect 2777 10523 2835 10529
rect 2777 10489 2789 10523
rect 2823 10520 2835 10523
rect 3605 10523 3663 10529
rect 3605 10520 3617 10523
rect 2823 10492 3617 10520
rect 2823 10489 2835 10492
rect 2777 10483 2835 10489
rect 3605 10489 3617 10492
rect 3651 10489 3663 10523
rect 3605 10483 3663 10489
rect 3712 10452 3740 10560
rect 3789 10557 3801 10560
rect 3835 10588 3847 10591
rect 5828 10588 5856 10628
rect 3835 10560 5856 10588
rect 5997 10591 6055 10597
rect 3835 10557 3847 10560
rect 3789 10551 3847 10557
rect 5997 10557 6009 10591
rect 6043 10588 6055 10591
rect 6043 10560 6316 10588
rect 6043 10557 6055 10560
rect 5997 10551 6055 10557
rect 5813 10523 5871 10529
rect 5813 10489 5825 10523
rect 5859 10520 5871 10523
rect 6178 10520 6184 10532
rect 5859 10492 6184 10520
rect 5859 10489 5871 10492
rect 5813 10483 5871 10489
rect 6178 10480 6184 10492
rect 6236 10480 6242 10532
rect 2700 10424 3740 10452
rect 5902 10412 5908 10464
rect 5960 10412 5966 10464
rect 6288 10452 6316 10560
rect 6380 10520 6408 10628
rect 6472 10588 6500 10696
rect 6564 10696 7297 10724
rect 6564 10665 6592 10696
rect 7285 10693 7297 10696
rect 7331 10724 7343 10727
rect 7742 10724 7748 10736
rect 7331 10696 7748 10724
rect 7331 10693 7343 10696
rect 7285 10687 7343 10693
rect 7742 10684 7748 10696
rect 7800 10684 7806 10736
rect 9674 10724 9680 10736
rect 8220 10696 9680 10724
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 6638 10616 6644 10668
rect 6696 10656 6702 10668
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 6696 10628 6745 10656
rect 6696 10616 6702 10628
rect 6733 10625 6745 10628
rect 6779 10656 6791 10659
rect 7193 10659 7251 10665
rect 7193 10656 7205 10659
rect 6779 10628 7205 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 7193 10625 7205 10628
rect 7239 10625 7251 10659
rect 7193 10619 7251 10625
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10656 7619 10659
rect 7650 10656 7656 10668
rect 7607 10628 7656 10656
rect 7607 10625 7619 10628
rect 7561 10619 7619 10625
rect 7650 10616 7656 10628
rect 7708 10656 7714 10668
rect 8220 10656 8248 10696
rect 9674 10684 9680 10696
rect 9732 10684 9738 10736
rect 12406 10696 18460 10724
rect 7708 10628 8248 10656
rect 8297 10659 8355 10665
rect 7708 10616 7714 10628
rect 8297 10625 8309 10659
rect 8343 10625 8355 10659
rect 8297 10619 8355 10625
rect 7282 10588 7288 10600
rect 6472 10560 7288 10588
rect 7282 10548 7288 10560
rect 7340 10548 7346 10600
rect 7374 10548 7380 10600
rect 7432 10548 7438 10600
rect 8312 10532 8340 10619
rect 8478 10616 8484 10668
rect 8536 10616 8542 10668
rect 9582 10616 9588 10668
rect 9640 10656 9646 10668
rect 12406 10656 12434 10696
rect 9640 10628 12434 10656
rect 9640 10616 9646 10628
rect 13078 10616 13084 10668
rect 13136 10616 13142 10668
rect 13446 10616 13452 10668
rect 13504 10656 13510 10668
rect 14001 10659 14059 10665
rect 14001 10656 14013 10659
rect 13504 10628 14013 10656
rect 13504 10616 13510 10628
rect 14001 10625 14013 10628
rect 14047 10656 14059 10659
rect 15286 10656 15292 10668
rect 14047 10628 15292 10656
rect 14047 10625 14059 10628
rect 14001 10619 14059 10625
rect 15286 10616 15292 10628
rect 15344 10616 15350 10668
rect 15746 10616 15752 10668
rect 15804 10656 15810 10668
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 15804 10628 15853 10656
rect 15804 10616 15810 10628
rect 15841 10625 15853 10628
rect 15887 10656 15899 10659
rect 16117 10659 16175 10665
rect 15887 10628 16068 10656
rect 15887 10625 15899 10628
rect 15841 10619 15899 10625
rect 13354 10548 13360 10600
rect 13412 10548 13418 10600
rect 8294 10520 8300 10532
rect 6380 10492 8300 10520
rect 8294 10480 8300 10492
rect 8352 10480 8358 10532
rect 9490 10480 9496 10532
rect 9548 10520 9554 10532
rect 13909 10523 13967 10529
rect 13909 10520 13921 10523
rect 9548 10492 13921 10520
rect 9548 10480 9554 10492
rect 13909 10489 13921 10492
rect 13955 10520 13967 10523
rect 14918 10520 14924 10532
rect 13955 10492 14924 10520
rect 13955 10489 13967 10492
rect 13909 10483 13967 10489
rect 14918 10480 14924 10492
rect 14976 10480 14982 10532
rect 15304 10520 15332 10616
rect 15654 10548 15660 10600
rect 15712 10588 15718 10600
rect 15933 10591 15991 10597
rect 15933 10588 15945 10591
rect 15712 10560 15945 10588
rect 15712 10548 15718 10560
rect 15933 10557 15945 10560
rect 15979 10557 15991 10591
rect 16040 10588 16068 10628
rect 16117 10625 16129 10659
rect 16163 10656 16175 10659
rect 16574 10656 16580 10668
rect 16163 10628 16580 10656
rect 16163 10625 16175 10628
rect 16117 10619 16175 10625
rect 16574 10616 16580 10628
rect 16632 10616 16638 10668
rect 18230 10616 18236 10668
rect 18288 10616 18294 10668
rect 18432 10665 18460 10696
rect 18417 10659 18475 10665
rect 18417 10625 18429 10659
rect 18463 10625 18475 10659
rect 18417 10619 18475 10625
rect 18598 10616 18604 10668
rect 18656 10616 18662 10668
rect 18690 10616 18696 10668
rect 18748 10616 18754 10668
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 19797 10659 19855 10665
rect 19797 10656 19809 10659
rect 19392 10628 19809 10656
rect 19392 10616 19398 10628
rect 19797 10625 19809 10628
rect 19843 10656 19855 10659
rect 20438 10656 20444 10668
rect 19843 10628 20444 10656
rect 19843 10625 19855 10628
rect 19797 10619 19855 10625
rect 20438 10616 20444 10628
rect 20496 10616 20502 10668
rect 19702 10588 19708 10600
rect 16040 10560 19708 10588
rect 15933 10551 15991 10557
rect 19702 10548 19708 10560
rect 19760 10548 19766 10600
rect 16206 10520 16212 10532
rect 15304 10492 16212 10520
rect 16206 10480 16212 10492
rect 16264 10480 16270 10532
rect 18509 10523 18567 10529
rect 18509 10489 18521 10523
rect 18555 10520 18567 10523
rect 19429 10523 19487 10529
rect 19429 10520 19441 10523
rect 18555 10492 19441 10520
rect 18555 10489 18567 10492
rect 18509 10483 18567 10489
rect 19429 10489 19441 10492
rect 19475 10489 19487 10523
rect 19429 10483 19487 10489
rect 6638 10452 6644 10464
rect 6288 10424 6644 10452
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 7561 10455 7619 10461
rect 7561 10421 7573 10455
rect 7607 10452 7619 10455
rect 8110 10452 8116 10464
rect 7607 10424 8116 10452
rect 7607 10421 7619 10424
rect 7561 10415 7619 10421
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 13173 10455 13231 10461
rect 13173 10421 13185 10455
rect 13219 10452 13231 10455
rect 13814 10452 13820 10464
rect 13219 10424 13820 10452
rect 13219 10421 13231 10424
rect 13173 10415 13231 10421
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 15654 10412 15660 10464
rect 15712 10412 15718 10464
rect 16117 10455 16175 10461
rect 16117 10421 16129 10455
rect 16163 10452 16175 10455
rect 16942 10452 16948 10464
rect 16163 10424 16948 10452
rect 16163 10421 16175 10424
rect 16117 10415 16175 10421
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 18966 10412 18972 10464
rect 19024 10412 19030 10464
rect 1104 10362 22816 10384
rect 1104 10310 3664 10362
rect 3716 10310 3728 10362
rect 3780 10310 3792 10362
rect 3844 10310 3856 10362
rect 3908 10310 3920 10362
rect 3972 10310 9092 10362
rect 9144 10310 9156 10362
rect 9208 10310 9220 10362
rect 9272 10310 9284 10362
rect 9336 10310 9348 10362
rect 9400 10310 14520 10362
rect 14572 10310 14584 10362
rect 14636 10310 14648 10362
rect 14700 10310 14712 10362
rect 14764 10310 14776 10362
rect 14828 10310 19948 10362
rect 20000 10310 20012 10362
rect 20064 10310 20076 10362
rect 20128 10310 20140 10362
rect 20192 10310 20204 10362
rect 20256 10310 22816 10362
rect 1104 10288 22816 10310
rect 2133 10251 2191 10257
rect 2133 10217 2145 10251
rect 2179 10248 2191 10251
rect 2179 10220 2268 10248
rect 2179 10217 2191 10220
rect 2133 10211 2191 10217
rect 2240 10180 2268 10220
rect 2314 10208 2320 10260
rect 2372 10208 2378 10260
rect 2682 10208 2688 10260
rect 2740 10248 2746 10260
rect 4157 10251 4215 10257
rect 4157 10248 4169 10251
rect 2740 10220 4169 10248
rect 2740 10208 2746 10220
rect 4157 10217 4169 10220
rect 4203 10217 4215 10251
rect 5626 10248 5632 10260
rect 4157 10211 4215 10217
rect 4264 10220 5632 10248
rect 2406 10180 2412 10192
rect 2240 10152 2412 10180
rect 2406 10140 2412 10152
rect 2464 10180 2470 10192
rect 3329 10183 3387 10189
rect 2464 10152 2912 10180
rect 2464 10140 2470 10152
rect 2682 10072 2688 10124
rect 2740 10112 2746 10124
rect 2777 10115 2835 10121
rect 2777 10112 2789 10115
rect 2740 10084 2789 10112
rect 2740 10072 2746 10084
rect 2777 10081 2789 10084
rect 2823 10081 2835 10115
rect 2777 10075 2835 10081
rect 1854 9936 1860 9988
rect 1912 9976 1918 9988
rect 1949 9979 2007 9985
rect 1949 9976 1961 9979
rect 1912 9948 1961 9976
rect 1912 9936 1918 9948
rect 1949 9945 1961 9948
rect 1995 9976 2007 9979
rect 2700 9976 2728 10072
rect 2884 10044 2912 10152
rect 3329 10149 3341 10183
rect 3375 10180 3387 10183
rect 3510 10180 3516 10192
rect 3375 10152 3516 10180
rect 3375 10149 3387 10152
rect 3329 10143 3387 10149
rect 3510 10140 3516 10152
rect 3568 10180 3574 10192
rect 4264 10180 4292 10220
rect 5626 10208 5632 10220
rect 5684 10208 5690 10260
rect 6365 10251 6423 10257
rect 6365 10217 6377 10251
rect 6411 10248 6423 10251
rect 6730 10248 6736 10260
rect 6411 10220 6736 10248
rect 6411 10217 6423 10220
rect 6365 10211 6423 10217
rect 6730 10208 6736 10220
rect 6788 10208 6794 10260
rect 8478 10208 8484 10260
rect 8536 10248 8542 10260
rect 9125 10251 9183 10257
rect 9125 10248 9137 10251
rect 8536 10220 9137 10248
rect 8536 10208 8542 10220
rect 9125 10217 9137 10220
rect 9171 10217 9183 10251
rect 9125 10211 9183 10217
rect 10318 10208 10324 10260
rect 10376 10208 10382 10260
rect 11238 10208 11244 10260
rect 11296 10208 11302 10260
rect 11609 10251 11667 10257
rect 11609 10217 11621 10251
rect 11655 10248 11667 10251
rect 12069 10251 12127 10257
rect 12069 10248 12081 10251
rect 11655 10220 12081 10248
rect 11655 10217 11667 10220
rect 11609 10211 11667 10217
rect 12069 10217 12081 10220
rect 12115 10217 12127 10251
rect 12069 10211 12127 10217
rect 12250 10208 12256 10260
rect 12308 10208 12314 10260
rect 12342 10208 12348 10260
rect 12400 10248 12406 10260
rect 13078 10248 13084 10260
rect 12400 10220 13084 10248
rect 12400 10208 12406 10220
rect 13078 10208 13084 10220
rect 13136 10248 13142 10260
rect 13173 10251 13231 10257
rect 13173 10248 13185 10251
rect 13136 10220 13185 10248
rect 13136 10208 13142 10220
rect 13173 10217 13185 10220
rect 13219 10217 13231 10251
rect 13173 10211 13231 10217
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 14277 10251 14335 10257
rect 14277 10248 14289 10251
rect 13872 10220 14289 10248
rect 13872 10208 13878 10220
rect 14277 10217 14289 10220
rect 14323 10217 14335 10251
rect 14277 10211 14335 10217
rect 18325 10251 18383 10257
rect 18325 10217 18337 10251
rect 18371 10248 18383 10251
rect 18966 10248 18972 10260
rect 18371 10220 18972 10248
rect 18371 10217 18383 10220
rect 18325 10211 18383 10217
rect 18966 10208 18972 10220
rect 19024 10208 19030 10260
rect 19794 10208 19800 10260
rect 19852 10248 19858 10260
rect 20073 10251 20131 10257
rect 20073 10248 20085 10251
rect 19852 10220 20085 10248
rect 19852 10208 19858 10220
rect 20073 10217 20085 10220
rect 20119 10217 20131 10251
rect 20073 10211 20131 10217
rect 3568 10152 4292 10180
rect 4341 10183 4399 10189
rect 3568 10140 3574 10152
rect 4341 10149 4353 10183
rect 4387 10180 4399 10183
rect 15378 10180 15384 10192
rect 4387 10152 6960 10180
rect 4387 10149 4399 10152
rect 4341 10143 4399 10149
rect 4154 10112 4160 10124
rect 4080 10084 4160 10112
rect 4080 10053 4108 10084
rect 4154 10072 4160 10084
rect 4212 10072 4218 10124
rect 6638 10112 6644 10124
rect 6012 10084 6644 10112
rect 3053 10047 3111 10053
rect 3053 10044 3065 10047
rect 2884 10016 3065 10044
rect 3053 10013 3065 10016
rect 3099 10013 3111 10047
rect 3053 10007 3111 10013
rect 4065 10047 4123 10053
rect 4065 10013 4077 10047
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 1995 9948 2728 9976
rect 2961 9979 3019 9985
rect 1995 9945 2007 9948
rect 1949 9939 2007 9945
rect 2961 9945 2973 9979
rect 3007 9976 3019 9979
rect 4264 9976 4292 10007
rect 4338 10004 4344 10056
rect 4396 10044 4402 10056
rect 4433 10047 4491 10053
rect 4433 10044 4445 10047
rect 4396 10016 4445 10044
rect 4396 10004 4402 10016
rect 4433 10013 4445 10016
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 5718 10004 5724 10056
rect 5776 10004 5782 10056
rect 5902 10004 5908 10056
rect 5960 10004 5966 10056
rect 6012 10053 6040 10084
rect 6638 10072 6644 10084
rect 6696 10072 6702 10124
rect 6932 10112 6960 10152
rect 11532 10152 15384 10180
rect 7374 10112 7380 10124
rect 6932 10084 7380 10112
rect 5997 10047 6055 10053
rect 5997 10013 6009 10047
rect 6043 10013 6055 10047
rect 5997 10007 6055 10013
rect 6089 10047 6147 10053
rect 6089 10013 6101 10047
rect 6135 10044 6147 10047
rect 6178 10044 6184 10056
rect 6135 10016 6184 10044
rect 6135 10013 6147 10016
rect 6089 10007 6147 10013
rect 6178 10004 6184 10016
rect 6236 10044 6242 10056
rect 7024 10053 7052 10084
rect 7374 10072 7380 10084
rect 7432 10112 7438 10124
rect 7469 10115 7527 10121
rect 7469 10112 7481 10115
rect 7432 10084 7481 10112
rect 7432 10072 7438 10084
rect 7469 10081 7481 10084
rect 7515 10081 7527 10115
rect 7469 10075 7527 10081
rect 8021 10115 8079 10121
rect 8021 10081 8033 10115
rect 8067 10112 8079 10115
rect 8294 10112 8300 10124
rect 8067 10084 8300 10112
rect 8067 10081 8079 10084
rect 8021 10075 8079 10081
rect 8294 10072 8300 10084
rect 8352 10112 8358 10124
rect 11532 10121 11560 10152
rect 15378 10140 15384 10152
rect 15436 10140 15442 10192
rect 17221 10183 17279 10189
rect 17221 10149 17233 10183
rect 17267 10180 17279 10183
rect 17957 10183 18015 10189
rect 17957 10180 17969 10183
rect 17267 10152 17969 10180
rect 17267 10149 17279 10152
rect 17221 10143 17279 10149
rect 17957 10149 17969 10152
rect 18003 10149 18015 10183
rect 17957 10143 18015 10149
rect 18414 10140 18420 10192
rect 18472 10140 18478 10192
rect 19242 10140 19248 10192
rect 19300 10180 19306 10192
rect 19300 10152 19932 10180
rect 19300 10140 19306 10152
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 8352 10084 9689 10112
rect 8352 10072 8358 10084
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 10413 10115 10471 10121
rect 10413 10081 10425 10115
rect 10459 10112 10471 10115
rect 11517 10115 11575 10121
rect 11517 10112 11529 10115
rect 10459 10084 11529 10112
rect 10459 10081 10471 10084
rect 10413 10075 10471 10081
rect 11517 10081 11529 10084
rect 11563 10081 11575 10115
rect 11517 10075 11575 10081
rect 13354 10072 13360 10124
rect 13412 10112 13418 10124
rect 13725 10115 13783 10121
rect 13725 10112 13737 10115
rect 13412 10084 13737 10112
rect 13412 10072 13418 10084
rect 13725 10081 13737 10084
rect 13771 10081 13783 10115
rect 13725 10075 13783 10081
rect 14918 10072 14924 10124
rect 14976 10072 14982 10124
rect 15654 10072 15660 10124
rect 15712 10112 15718 10124
rect 15841 10115 15899 10121
rect 15841 10112 15853 10115
rect 15712 10084 15853 10112
rect 15712 10072 15718 10084
rect 15841 10081 15853 10084
rect 15887 10081 15899 10115
rect 15841 10075 15899 10081
rect 16022 10072 16028 10124
rect 16080 10112 16086 10124
rect 16577 10115 16635 10121
rect 16577 10112 16589 10115
rect 16080 10084 16589 10112
rect 16080 10072 16086 10084
rect 16577 10081 16589 10084
rect 16623 10081 16635 10115
rect 16577 10075 16635 10081
rect 16761 10115 16819 10121
rect 16761 10081 16773 10115
rect 16807 10112 16819 10115
rect 17034 10112 17040 10124
rect 16807 10084 17040 10112
rect 16807 10081 16819 10084
rect 16761 10075 16819 10081
rect 17034 10072 17040 10084
rect 17092 10072 17098 10124
rect 18506 10072 18512 10124
rect 18564 10072 18570 10124
rect 18601 10115 18659 10121
rect 18601 10081 18613 10115
rect 18647 10112 18659 10115
rect 18647 10084 19840 10112
rect 18647 10081 18659 10084
rect 18601 10075 18659 10081
rect 6917 10047 6975 10053
rect 6917 10044 6929 10047
rect 6236 10016 6929 10044
rect 6236 10004 6242 10016
rect 6917 10013 6929 10016
rect 6963 10013 6975 10047
rect 6917 10007 6975 10013
rect 7009 10047 7067 10053
rect 7009 10013 7021 10047
rect 7055 10013 7067 10047
rect 7009 10007 7067 10013
rect 7650 10004 7656 10056
rect 7708 10004 7714 10056
rect 9582 10004 9588 10056
rect 9640 10004 9646 10056
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10044 10563 10047
rect 10594 10044 10600 10056
rect 10551 10016 10600 10044
rect 10551 10013 10563 10016
rect 10505 10007 10563 10013
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 11609 10047 11667 10053
rect 11609 10013 11621 10047
rect 11655 10044 11667 10047
rect 11698 10044 11704 10056
rect 11655 10016 11704 10044
rect 11655 10013 11667 10016
rect 11609 10007 11667 10013
rect 11698 10004 11704 10016
rect 11756 10004 11762 10056
rect 13446 10004 13452 10056
rect 13504 10004 13510 10056
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10044 13599 10047
rect 14458 10047 14516 10053
rect 14458 10044 14470 10047
rect 13587 10016 14470 10044
rect 13587 10013 13599 10016
rect 13541 10007 13599 10013
rect 14458 10013 14470 10016
rect 14504 10044 14516 10047
rect 14504 10016 14780 10044
rect 14504 10013 14516 10016
rect 14458 10007 14516 10013
rect 3007 9948 4476 9976
rect 3007 9945 3019 9948
rect 2961 9939 3019 9945
rect 4448 9920 4476 9948
rect 4706 9936 4712 9988
rect 4764 9936 4770 9988
rect 5626 9936 5632 9988
rect 5684 9976 5690 9988
rect 7837 9979 7895 9985
rect 7837 9976 7849 9979
rect 5684 9948 7849 9976
rect 5684 9936 5690 9948
rect 7837 9945 7849 9948
rect 7883 9945 7895 9979
rect 7837 9939 7895 9945
rect 10778 9936 10784 9988
rect 10836 9976 10842 9988
rect 12237 9979 12295 9985
rect 12237 9976 12249 9979
rect 10836 9948 12249 9976
rect 10836 9936 10842 9948
rect 12237 9945 12249 9948
rect 12283 9976 12295 9979
rect 12342 9976 12348 9988
rect 12283 9948 12348 9976
rect 12283 9945 12295 9948
rect 12237 9939 12295 9945
rect 12342 9936 12348 9948
rect 12400 9936 12406 9988
rect 12434 9936 12440 9988
rect 12492 9936 12498 9988
rect 13357 9979 13415 9985
rect 13357 9945 13369 9979
rect 13403 9976 13415 9979
rect 14752 9976 14780 10016
rect 14826 10004 14832 10056
rect 14884 10044 14890 10056
rect 15194 10044 15200 10056
rect 14884 10016 15200 10044
rect 14884 10004 14890 10016
rect 15194 10004 15200 10016
rect 15252 10004 15258 10056
rect 15470 10004 15476 10056
rect 15528 10004 15534 10056
rect 15746 10004 15752 10056
rect 15804 10004 15810 10056
rect 18046 10004 18052 10056
rect 18104 10044 18110 10056
rect 18616 10044 18644 10075
rect 18104 10016 18644 10044
rect 18104 10004 18110 10016
rect 19426 10004 19432 10056
rect 19484 10004 19490 10056
rect 19812 10053 19840 10084
rect 19613 10047 19671 10053
rect 19613 10013 19625 10047
rect 19659 10013 19671 10047
rect 19613 10007 19671 10013
rect 19705 10047 19763 10053
rect 19705 10013 19717 10047
rect 19751 10013 19763 10047
rect 19705 10007 19763 10013
rect 19797 10047 19855 10053
rect 19797 10013 19809 10047
rect 19843 10013 19855 10047
rect 19797 10007 19855 10013
rect 15286 9976 15292 9988
rect 13403 9948 13676 9976
rect 14752 9948 15292 9976
rect 13403 9945 13415 9948
rect 13357 9939 13415 9945
rect 1762 9868 1768 9920
rect 1820 9908 1826 9920
rect 2159 9911 2217 9917
rect 2159 9908 2171 9911
rect 1820 9880 2171 9908
rect 1820 9868 1826 9880
rect 2159 9877 2171 9880
rect 2205 9908 2217 9911
rect 3142 9908 3148 9920
rect 2205 9880 3148 9908
rect 2205 9877 2217 9880
rect 2159 9871 2217 9877
rect 3142 9868 3148 9880
rect 3200 9868 3206 9920
rect 4430 9868 4436 9920
rect 4488 9868 4494 9920
rect 6178 9868 6184 9920
rect 6236 9908 6242 9920
rect 6362 9908 6368 9920
rect 6236 9880 6368 9908
rect 6236 9868 6242 9880
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 7742 9868 7748 9920
rect 7800 9868 7806 9920
rect 9490 9868 9496 9920
rect 9548 9868 9554 9920
rect 10502 9868 10508 9920
rect 10560 9908 10566 9920
rect 10689 9911 10747 9917
rect 10689 9908 10701 9911
rect 10560 9880 10701 9908
rect 10560 9868 10566 9880
rect 10689 9877 10701 9880
rect 10735 9908 10747 9911
rect 10962 9908 10968 9920
rect 10735 9880 10968 9908
rect 10735 9877 10747 9880
rect 10689 9871 10747 9877
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 13648 9908 13676 9948
rect 15286 9936 15292 9948
rect 15344 9976 15350 9988
rect 15838 9976 15844 9988
rect 15344 9948 15844 9976
rect 15344 9936 15350 9948
rect 15838 9936 15844 9948
rect 15896 9936 15902 9988
rect 16574 9936 16580 9988
rect 16632 9976 16638 9988
rect 16853 9979 16911 9985
rect 16853 9976 16865 9979
rect 16632 9948 16865 9976
rect 16632 9936 16638 9948
rect 16853 9945 16865 9948
rect 16899 9945 16911 9979
rect 16853 9939 16911 9945
rect 17954 9936 17960 9988
rect 18012 9976 18018 9988
rect 19628 9976 19656 10007
rect 18012 9948 19656 9976
rect 19720 9976 19748 10007
rect 19904 9976 19932 10152
rect 19720 9948 19932 9976
rect 18012 9936 18018 9948
rect 14461 9911 14519 9917
rect 14461 9908 14473 9911
rect 13648 9880 14473 9908
rect 14461 9877 14473 9880
rect 14507 9908 14519 9911
rect 15102 9908 15108 9920
rect 14507 9880 15108 9908
rect 14507 9877 14519 9880
rect 14461 9871 14519 9877
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 15930 9868 15936 9920
rect 15988 9908 15994 9920
rect 20346 9908 20352 9920
rect 15988 9880 20352 9908
rect 15988 9868 15994 9880
rect 20346 9868 20352 9880
rect 20404 9868 20410 9920
rect 1104 9818 22976 9840
rect 1104 9766 6378 9818
rect 6430 9766 6442 9818
rect 6494 9766 6506 9818
rect 6558 9766 6570 9818
rect 6622 9766 6634 9818
rect 6686 9766 11806 9818
rect 11858 9766 11870 9818
rect 11922 9766 11934 9818
rect 11986 9766 11998 9818
rect 12050 9766 12062 9818
rect 12114 9766 17234 9818
rect 17286 9766 17298 9818
rect 17350 9766 17362 9818
rect 17414 9766 17426 9818
rect 17478 9766 17490 9818
rect 17542 9766 22662 9818
rect 22714 9766 22726 9818
rect 22778 9766 22790 9818
rect 22842 9766 22854 9818
rect 22906 9766 22918 9818
rect 22970 9766 22976 9818
rect 1104 9744 22976 9766
rect 1854 9664 1860 9716
rect 1912 9664 1918 9716
rect 2222 9664 2228 9716
rect 2280 9704 2286 9716
rect 5718 9704 5724 9716
rect 2280 9676 5724 9704
rect 2280 9664 2286 9676
rect 5718 9664 5724 9676
rect 5776 9704 5782 9716
rect 6730 9713 6736 9716
rect 6717 9707 6736 9713
rect 5776 9676 6684 9704
rect 5776 9664 5782 9676
rect 2041 9639 2099 9645
rect 2041 9605 2053 9639
rect 2087 9636 2099 9639
rect 2406 9636 2412 9648
rect 2087 9608 2412 9636
rect 2087 9605 2099 9608
rect 2041 9599 2099 9605
rect 2406 9596 2412 9608
rect 2464 9596 2470 9648
rect 5626 9596 5632 9648
rect 5684 9596 5690 9648
rect 6656 9636 6684 9676
rect 6717 9673 6729 9707
rect 6717 9667 6736 9673
rect 6730 9664 6736 9667
rect 6788 9664 6794 9716
rect 8205 9707 8263 9713
rect 8205 9673 8217 9707
rect 8251 9704 8263 9707
rect 8570 9704 8576 9716
rect 8251 9676 8576 9704
rect 8251 9673 8263 9676
rect 8205 9667 8263 9673
rect 8570 9664 8576 9676
rect 8628 9664 8634 9716
rect 9217 9707 9275 9713
rect 9217 9673 9229 9707
rect 9263 9704 9275 9707
rect 9490 9704 9496 9716
rect 9263 9676 9496 9704
rect 9263 9673 9275 9676
rect 9217 9667 9275 9673
rect 9490 9664 9496 9676
rect 9548 9664 9554 9716
rect 10778 9664 10784 9716
rect 10836 9664 10842 9716
rect 12434 9704 12440 9716
rect 11900 9676 12440 9704
rect 6917 9639 6975 9645
rect 6917 9636 6929 9639
rect 6656 9608 6929 9636
rect 6917 9605 6929 9608
rect 6963 9605 6975 9639
rect 6917 9599 6975 9605
rect 7282 9596 7288 9648
rect 7340 9636 7346 9648
rect 7926 9636 7932 9648
rect 7340 9608 7932 9636
rect 7340 9596 7346 9608
rect 7926 9596 7932 9608
rect 7984 9596 7990 9648
rect 8294 9596 8300 9648
rect 8352 9596 8358 9648
rect 10597 9639 10655 9645
rect 10597 9605 10609 9639
rect 10643 9636 10655 9639
rect 10796 9636 10824 9664
rect 11900 9645 11928 9676
rect 12434 9664 12440 9676
rect 12492 9704 12498 9716
rect 16114 9704 16120 9716
rect 12492 9676 16120 9704
rect 12492 9664 12498 9676
rect 16114 9664 16120 9676
rect 16172 9664 16178 9716
rect 16224 9676 16436 9704
rect 11885 9639 11943 9645
rect 11885 9636 11897 9639
rect 10643 9608 10824 9636
rect 10980 9608 11897 9636
rect 10643 9605 10655 9608
rect 10597 9599 10655 9605
rect 10980 9580 11008 9608
rect 11885 9605 11897 9608
rect 11931 9605 11943 9639
rect 11885 9599 11943 9605
rect 13541 9639 13599 9645
rect 13541 9605 13553 9639
rect 13587 9636 13599 9639
rect 15194 9636 15200 9648
rect 13587 9608 15200 9636
rect 13587 9605 13599 9608
rect 13541 9599 13599 9605
rect 15194 9596 15200 9608
rect 15252 9636 15258 9648
rect 16022 9636 16028 9648
rect 15252 9608 16028 9636
rect 15252 9596 15258 9608
rect 16022 9596 16028 9608
rect 16080 9596 16086 9648
rect 16224 9636 16252 9676
rect 16132 9608 16252 9636
rect 1762 9528 1768 9580
rect 1820 9528 1826 9580
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9568 5871 9571
rect 7742 9568 7748 9580
rect 5859 9540 7748 9568
rect 5859 9537 5871 9540
rect 5813 9531 5871 9537
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 8202 9568 8208 9580
rect 8067 9540 8208 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 9125 9571 9183 9577
rect 9125 9568 9137 9571
rect 8312 9540 9137 9568
rect 8110 9460 8116 9512
rect 8168 9460 8174 9512
rect 2038 9392 2044 9444
rect 2096 9392 2102 9444
rect 5997 9435 6055 9441
rect 5997 9401 6009 9435
rect 6043 9432 6055 9435
rect 6043 9404 6776 9432
rect 6043 9401 6055 9404
rect 5997 9395 6055 9401
rect 6270 9324 6276 9376
rect 6328 9364 6334 9376
rect 6748 9373 6776 9404
rect 7282 9392 7288 9444
rect 7340 9432 7346 9444
rect 8312 9432 8340 9540
rect 9125 9537 9137 9540
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9568 9367 9571
rect 9582 9568 9588 9580
rect 9355 9540 9588 9568
rect 9355 9537 9367 9540
rect 9309 9531 9367 9537
rect 9582 9528 9588 9540
rect 9640 9528 9646 9580
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 10873 9571 10931 9577
rect 10873 9537 10885 9571
rect 10919 9568 10931 9571
rect 10962 9568 10968 9580
rect 10919 9540 10968 9568
rect 10919 9537 10931 9540
rect 10873 9531 10931 9537
rect 10796 9500 10824 9531
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 11422 9528 11428 9580
rect 11480 9568 11486 9580
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 11480 9540 11713 9568
rect 11480 9528 11486 9540
rect 11701 9537 11713 9540
rect 11747 9568 11759 9571
rect 11977 9571 12035 9577
rect 11747 9540 11928 9568
rect 11747 9537 11759 9540
rect 11701 9531 11759 9537
rect 11900 9500 11928 9540
rect 11977 9537 11989 9571
rect 12023 9568 12035 9571
rect 12342 9568 12348 9580
rect 12023 9540 12348 9568
rect 12023 9537 12035 9540
rect 11977 9531 12035 9537
rect 12342 9528 12348 9540
rect 12400 9528 12406 9580
rect 13262 9528 13268 9580
rect 13320 9528 13326 9580
rect 13725 9571 13783 9577
rect 13725 9537 13737 9571
rect 13771 9568 13783 9571
rect 13998 9568 14004 9580
rect 13771 9540 14004 9568
rect 13771 9537 13783 9540
rect 13725 9531 13783 9537
rect 13998 9528 14004 9540
rect 14056 9568 14062 9580
rect 14826 9568 14832 9580
rect 14056 9540 14832 9568
rect 14056 9528 14062 9540
rect 14826 9528 14832 9540
rect 14884 9528 14890 9580
rect 15930 9528 15936 9580
rect 15988 9528 15994 9580
rect 12250 9500 12256 9512
rect 10796 9472 11836 9500
rect 11900 9472 12256 9500
rect 7340 9404 8340 9432
rect 7340 9392 7346 9404
rect 10594 9392 10600 9444
rect 10652 9392 10658 9444
rect 11698 9392 11704 9444
rect 11756 9392 11762 9444
rect 11808 9432 11836 9472
rect 12250 9460 12256 9472
rect 12308 9500 12314 9512
rect 15470 9500 15476 9512
rect 12308 9472 15476 9500
rect 12308 9460 12314 9472
rect 15470 9460 15476 9472
rect 15528 9460 15534 9512
rect 15841 9503 15899 9509
rect 15841 9469 15853 9503
rect 15887 9500 15899 9503
rect 16132 9500 16160 9608
rect 16298 9596 16304 9648
rect 16356 9596 16362 9648
rect 16408 9636 16436 9676
rect 18782 9664 18788 9716
rect 18840 9664 18846 9716
rect 17954 9636 17960 9648
rect 16408 9608 17960 9636
rect 17954 9596 17960 9608
rect 18012 9596 18018 9648
rect 18800 9636 18828 9664
rect 18800 9608 19012 9636
rect 16209 9571 16267 9577
rect 16209 9537 16221 9571
rect 16255 9568 16267 9571
rect 18690 9568 18696 9580
rect 16255 9540 18696 9568
rect 16255 9537 16267 9540
rect 16209 9531 16267 9537
rect 15887 9472 16160 9500
rect 15887 9469 15899 9472
rect 15841 9463 15899 9469
rect 12526 9432 12532 9444
rect 11808 9404 12532 9432
rect 12526 9392 12532 9404
rect 12584 9432 12590 9444
rect 13354 9432 13360 9444
rect 12584 9404 13360 9432
rect 12584 9392 12590 9404
rect 13354 9392 13360 9404
rect 13412 9432 13418 9444
rect 13412 9404 15792 9432
rect 13412 9392 13418 9404
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 6328 9336 6561 9364
rect 6328 9324 6334 9336
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 6549 9327 6607 9333
rect 6733 9367 6791 9373
rect 6733 9333 6745 9367
rect 6779 9333 6791 9367
rect 6733 9327 6791 9333
rect 13446 9324 13452 9376
rect 13504 9364 13510 9376
rect 15657 9367 15715 9373
rect 15657 9364 15669 9367
rect 13504 9336 15669 9364
rect 13504 9324 13510 9336
rect 15657 9333 15669 9336
rect 15703 9333 15715 9367
rect 15764 9364 15792 9404
rect 16224 9364 16252 9531
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 18785 9571 18843 9577
rect 18785 9537 18797 9571
rect 18831 9568 18843 9571
rect 18874 9568 18880 9580
rect 18831 9540 18880 9568
rect 18831 9537 18843 9540
rect 18785 9531 18843 9537
rect 18874 9528 18880 9540
rect 18932 9528 18938 9580
rect 18984 9577 19012 9608
rect 18969 9571 19027 9577
rect 18969 9537 18981 9571
rect 19015 9537 19027 9571
rect 18969 9531 19027 9537
rect 16390 9460 16396 9512
rect 16448 9500 16454 9512
rect 18509 9503 18567 9509
rect 18509 9500 18521 9503
rect 16448 9472 18521 9500
rect 16448 9460 16454 9472
rect 18509 9469 18521 9472
rect 18555 9469 18567 9503
rect 18509 9463 18567 9469
rect 15764 9336 16252 9364
rect 15657 9327 15715 9333
rect 1104 9274 22816 9296
rect 1104 9222 3664 9274
rect 3716 9222 3728 9274
rect 3780 9222 3792 9274
rect 3844 9222 3856 9274
rect 3908 9222 3920 9274
rect 3972 9222 9092 9274
rect 9144 9222 9156 9274
rect 9208 9222 9220 9274
rect 9272 9222 9284 9274
rect 9336 9222 9348 9274
rect 9400 9222 14520 9274
rect 14572 9222 14584 9274
rect 14636 9222 14648 9274
rect 14700 9222 14712 9274
rect 14764 9222 14776 9274
rect 14828 9222 19948 9274
rect 20000 9222 20012 9274
rect 20064 9222 20076 9274
rect 20128 9222 20140 9274
rect 20192 9222 20204 9274
rect 20256 9222 22816 9274
rect 1104 9200 22816 9222
rect 2041 9163 2099 9169
rect 2041 9129 2053 9163
rect 2087 9160 2099 9163
rect 2406 9160 2412 9172
rect 2087 9132 2412 9160
rect 2087 9129 2099 9132
rect 2041 9123 2099 9129
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 7653 9163 7711 9169
rect 7653 9129 7665 9163
rect 7699 9160 7711 9163
rect 7742 9160 7748 9172
rect 7699 9132 7748 9160
rect 7699 9129 7711 9132
rect 7653 9123 7711 9129
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 13170 9120 13176 9172
rect 13228 9120 13234 9172
rect 13354 9120 13360 9172
rect 13412 9120 13418 9172
rect 15746 9120 15752 9172
rect 15804 9120 15810 9172
rect 16114 9120 16120 9172
rect 16172 9120 16178 9172
rect 18877 9163 18935 9169
rect 18877 9129 18889 9163
rect 18923 9160 18935 9163
rect 19426 9160 19432 9172
rect 18923 9132 19432 9160
rect 18923 9129 18935 9132
rect 18877 9123 18935 9129
rect 19426 9120 19432 9132
rect 19484 9120 19490 9172
rect 2409 9027 2467 9033
rect 2409 8993 2421 9027
rect 2455 9024 2467 9027
rect 2590 9024 2596 9036
rect 2455 8996 2596 9024
rect 2455 8993 2467 8996
rect 2409 8987 2467 8993
rect 2590 8984 2596 8996
rect 2648 9024 2654 9036
rect 4338 9024 4344 9036
rect 2648 8996 4344 9024
rect 2648 8984 2654 8996
rect 4338 8984 4344 8996
rect 4396 9024 4402 9036
rect 4433 9027 4491 9033
rect 4433 9024 4445 9027
rect 4396 8996 4445 9024
rect 4396 8984 4402 8996
rect 4433 8993 4445 8996
rect 4479 9024 4491 9027
rect 5442 9024 5448 9036
rect 4479 8996 5448 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 5442 8984 5448 8996
rect 5500 9024 5506 9036
rect 7282 9024 7288 9036
rect 5500 8996 7288 9024
rect 5500 8984 5506 8996
rect 7282 8984 7288 8996
rect 7340 8984 7346 9036
rect 13354 9024 13360 9036
rect 12452 8996 13360 9024
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8925 2283 8959
rect 2225 8919 2283 8925
rect 2240 8888 2268 8919
rect 4246 8916 4252 8968
rect 4304 8916 4310 8968
rect 7466 8916 7472 8968
rect 7524 8916 7530 8968
rect 12452 8965 12480 8996
rect 13354 8984 13360 8996
rect 13412 8984 13418 9036
rect 18417 9027 18475 9033
rect 18417 8993 18429 9027
rect 18463 9024 18475 9027
rect 19334 9024 19340 9036
rect 18463 8996 19340 9024
rect 18463 8993 18475 8996
rect 18417 8987 18475 8993
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8925 12495 8959
rect 12437 8919 12495 8925
rect 12618 8916 12624 8968
rect 12676 8916 12682 8968
rect 15286 8916 15292 8968
rect 15344 8956 15350 8968
rect 15933 8959 15991 8965
rect 15933 8956 15945 8959
rect 15344 8928 15945 8956
rect 15344 8916 15350 8928
rect 15933 8925 15945 8928
rect 15979 8925 15991 8959
rect 15933 8919 15991 8925
rect 16206 8916 16212 8968
rect 16264 8956 16270 8968
rect 16301 8959 16359 8965
rect 16301 8956 16313 8959
rect 16264 8928 16313 8956
rect 16264 8916 16270 8928
rect 16301 8925 16313 8928
rect 16347 8925 16359 8959
rect 16301 8919 16359 8925
rect 18322 8916 18328 8968
rect 18380 8956 18386 8968
rect 18509 8959 18567 8965
rect 18509 8956 18521 8959
rect 18380 8928 18521 8956
rect 18380 8916 18386 8928
rect 18509 8925 18521 8928
rect 18555 8925 18567 8959
rect 18509 8919 18567 8925
rect 18690 8916 18696 8968
rect 18748 8916 18754 8968
rect 5994 8888 6000 8900
rect 2240 8860 6000 8888
rect 5994 8848 6000 8860
rect 6052 8848 6058 8900
rect 12158 8848 12164 8900
rect 12216 8888 12222 8900
rect 13341 8891 13399 8897
rect 12216 8860 13308 8888
rect 12216 8848 12222 8860
rect 4065 8823 4123 8829
rect 4065 8789 4077 8823
rect 4111 8820 4123 8823
rect 4154 8820 4160 8832
rect 4111 8792 4160 8820
rect 4111 8789 4123 8792
rect 4065 8783 4123 8789
rect 4154 8780 4160 8792
rect 4212 8780 4218 8832
rect 12250 8780 12256 8832
rect 12308 8820 12314 8832
rect 12529 8823 12587 8829
rect 12529 8820 12541 8823
rect 12308 8792 12541 8820
rect 12308 8780 12314 8792
rect 12529 8789 12541 8792
rect 12575 8789 12587 8823
rect 13280 8820 13308 8860
rect 13341 8857 13353 8891
rect 13387 8888 13399 8891
rect 13446 8888 13452 8900
rect 13387 8860 13452 8888
rect 13387 8857 13399 8860
rect 13341 8851 13399 8857
rect 13446 8848 13452 8860
rect 13504 8848 13510 8900
rect 13541 8891 13599 8897
rect 13541 8857 13553 8891
rect 13587 8888 13599 8891
rect 16390 8888 16396 8900
rect 13587 8860 16396 8888
rect 13587 8857 13599 8860
rect 13541 8851 13599 8857
rect 13556 8820 13584 8851
rect 16390 8848 16396 8860
rect 16448 8848 16454 8900
rect 13280 8792 13584 8820
rect 12529 8783 12587 8789
rect 1104 8730 22976 8752
rect 1104 8678 6378 8730
rect 6430 8678 6442 8730
rect 6494 8678 6506 8730
rect 6558 8678 6570 8730
rect 6622 8678 6634 8730
rect 6686 8678 11806 8730
rect 11858 8678 11870 8730
rect 11922 8678 11934 8730
rect 11986 8678 11998 8730
rect 12050 8678 12062 8730
rect 12114 8678 17234 8730
rect 17286 8678 17298 8730
rect 17350 8678 17362 8730
rect 17414 8678 17426 8730
rect 17478 8678 17490 8730
rect 17542 8678 22662 8730
rect 22714 8678 22726 8730
rect 22778 8678 22790 8730
rect 22842 8678 22854 8730
rect 22906 8678 22918 8730
rect 22970 8678 22976 8730
rect 1104 8656 22976 8678
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 4614 8616 4620 8628
rect 4295 8588 4620 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 6822 8625 6828 8628
rect 6818 8616 6828 8625
rect 6783 8588 6828 8616
rect 6818 8579 6828 8588
rect 6822 8576 6828 8579
rect 6880 8576 6886 8628
rect 8481 8619 8539 8625
rect 8481 8616 8493 8619
rect 7484 8588 8493 8616
rect 4338 8548 4344 8560
rect 3620 8520 4344 8548
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8480 3019 8483
rect 3142 8480 3148 8492
rect 3007 8452 3148 8480
rect 3007 8449 3019 8452
rect 2961 8443 3019 8449
rect 3142 8440 3148 8452
rect 3200 8480 3206 8492
rect 3510 8480 3516 8492
rect 3200 8452 3516 8480
rect 3200 8440 3206 8452
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 3620 8489 3648 8520
rect 4338 8508 4344 8520
rect 4396 8508 4402 8560
rect 7374 8548 7380 8560
rect 6656 8520 7380 8548
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 3789 8483 3847 8489
rect 3789 8449 3801 8483
rect 3835 8449 3847 8483
rect 3789 8443 3847 8449
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8449 3939 8483
rect 3881 8443 3939 8449
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8480 4031 8483
rect 4154 8480 4160 8492
rect 4019 8452 4160 8480
rect 4019 8449 4031 8452
rect 3973 8443 4031 8449
rect 3053 8415 3111 8421
rect 3053 8381 3065 8415
rect 3099 8412 3111 8415
rect 3804 8412 3832 8443
rect 3099 8384 3832 8412
rect 3099 8381 3111 8384
rect 3053 8375 3111 8381
rect 3418 8304 3424 8356
rect 3476 8344 3482 8356
rect 3896 8344 3924 8443
rect 4154 8440 4160 8452
rect 4212 8440 4218 8492
rect 4890 8440 4896 8492
rect 4948 8440 4954 8492
rect 5902 8440 5908 8492
rect 5960 8480 5966 8492
rect 6656 8489 6684 8520
rect 7374 8508 7380 8520
rect 7432 8508 7438 8560
rect 6641 8483 6699 8489
rect 6641 8480 6653 8483
rect 5960 8452 6653 8480
rect 5960 8440 5966 8452
rect 6641 8449 6653 8452
rect 6687 8449 6699 8483
rect 6641 8443 6699 8449
rect 6730 8440 6736 8492
rect 6788 8440 6794 8492
rect 6914 8440 6920 8492
rect 6972 8440 6978 8492
rect 7282 8440 7288 8492
rect 7340 8480 7346 8492
rect 7484 8489 7512 8588
rect 8481 8585 8493 8588
rect 8527 8585 8539 8619
rect 8481 8579 8539 8585
rect 10689 8619 10747 8625
rect 10689 8585 10701 8619
rect 10735 8585 10747 8619
rect 10689 8579 10747 8585
rect 10704 8548 10732 8579
rect 11606 8576 11612 8628
rect 11664 8616 11670 8628
rect 11885 8619 11943 8625
rect 11885 8616 11897 8619
rect 11664 8588 11897 8616
rect 11664 8576 11670 8588
rect 11885 8585 11897 8588
rect 11931 8585 11943 8619
rect 11885 8579 11943 8585
rect 12069 8619 12127 8625
rect 12069 8585 12081 8619
rect 12115 8616 12127 8619
rect 12158 8616 12164 8628
rect 12115 8588 12164 8616
rect 12115 8585 12127 8588
rect 12069 8579 12127 8585
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 13630 8576 13636 8628
rect 13688 8616 13694 8628
rect 17865 8619 17923 8625
rect 13688 8588 15700 8616
rect 13688 8576 13694 8588
rect 7576 8520 10732 8548
rect 7576 8489 7604 8520
rect 11146 8508 11152 8560
rect 11204 8508 11210 8560
rect 12618 8508 12624 8560
rect 12676 8548 12682 8560
rect 15194 8548 15200 8560
rect 12676 8520 15200 8548
rect 12676 8508 12682 8520
rect 7469 8483 7527 8489
rect 7469 8480 7481 8483
rect 7340 8452 7481 8480
rect 7340 8440 7346 8452
rect 7469 8449 7481 8452
rect 7515 8449 7527 8483
rect 7469 8443 7527 8449
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 8757 8483 8815 8489
rect 8757 8449 8769 8483
rect 8803 8480 8815 8483
rect 9582 8480 9588 8492
rect 8803 8452 9588 8480
rect 8803 8449 8815 8452
rect 8757 8443 8815 8449
rect 4706 8372 4712 8424
rect 4764 8412 4770 8424
rect 5920 8412 5948 8440
rect 4764 8384 5948 8412
rect 4764 8372 4770 8384
rect 5994 8372 6000 8424
rect 6052 8412 6058 8424
rect 7760 8412 7788 8443
rect 9582 8440 9588 8452
rect 9640 8440 9646 8492
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8480 9735 8483
rect 11422 8480 11428 8492
rect 9723 8452 11428 8480
rect 9723 8449 9735 8452
rect 9677 8443 9735 8449
rect 11422 8440 11428 8452
rect 11480 8440 11486 8492
rect 12912 8489 12940 8520
rect 13832 8489 13860 8520
rect 15194 8508 15200 8520
rect 15252 8508 15258 8560
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8449 13139 8483
rect 13081 8443 13139 8449
rect 13817 8483 13875 8489
rect 13817 8449 13829 8483
rect 13863 8449 13875 8483
rect 13817 8443 13875 8449
rect 6052 8384 7788 8412
rect 6052 8372 6058 8384
rect 8478 8372 8484 8424
rect 8536 8412 8542 8424
rect 9309 8415 9367 8421
rect 9309 8412 9321 8415
rect 8536 8384 9321 8412
rect 8536 8372 8542 8384
rect 9309 8381 9321 8384
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 9398 8372 9404 8424
rect 9456 8372 9462 8424
rect 9766 8372 9772 8424
rect 9824 8412 9830 8424
rect 9824 8384 10079 8412
rect 9824 8372 9830 8384
rect 3476 8316 3924 8344
rect 3476 8304 3482 8316
rect 7466 8304 7472 8356
rect 7524 8344 7530 8356
rect 7653 8347 7711 8353
rect 7653 8344 7665 8347
rect 7524 8316 7665 8344
rect 7524 8304 7530 8316
rect 7653 8313 7665 8316
rect 7699 8313 7711 8347
rect 7653 8307 7711 8313
rect 7929 8347 7987 8353
rect 7929 8313 7941 8347
rect 7975 8344 7987 8347
rect 9490 8344 9496 8356
rect 7975 8316 9496 8344
rect 7975 8313 7987 8316
rect 7929 8307 7987 8313
rect 9490 8304 9496 8316
rect 9548 8304 9554 8356
rect 5074 8236 5080 8288
rect 5132 8236 5138 8288
rect 8938 8236 8944 8288
rect 8996 8276 9002 8288
rect 9398 8276 9404 8288
rect 8996 8248 9404 8276
rect 8996 8236 9002 8248
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 9950 8236 9956 8288
rect 10008 8236 10014 8288
rect 10051 8276 10079 8384
rect 10686 8372 10692 8424
rect 10744 8372 10750 8424
rect 13096 8412 13124 8443
rect 14366 8440 14372 8492
rect 14424 8480 14430 8492
rect 14461 8483 14519 8489
rect 14461 8480 14473 8483
rect 14424 8452 14473 8480
rect 14424 8440 14430 8452
rect 14461 8449 14473 8452
rect 14507 8449 14519 8483
rect 14461 8443 14519 8449
rect 14645 8483 14703 8489
rect 14645 8449 14657 8483
rect 14691 8480 14703 8483
rect 14918 8480 14924 8492
rect 14691 8452 14924 8480
rect 14691 8449 14703 8452
rect 14645 8443 14703 8449
rect 14918 8440 14924 8452
rect 14976 8440 14982 8492
rect 15672 8489 15700 8588
rect 17865 8585 17877 8619
rect 17911 8616 17923 8619
rect 17954 8616 17960 8628
rect 17911 8588 17960 8616
rect 17911 8585 17923 8588
rect 17865 8579 17923 8585
rect 17954 8576 17960 8588
rect 18012 8576 18018 8628
rect 16482 8548 16488 8560
rect 16132 8520 16488 8548
rect 16132 8489 16160 8520
rect 16482 8508 16488 8520
rect 16540 8508 16546 8560
rect 18322 8548 18328 8560
rect 17788 8520 18328 8548
rect 17788 8489 17816 8520
rect 18322 8508 18328 8520
rect 18380 8508 18386 8560
rect 15657 8483 15715 8489
rect 15657 8449 15669 8483
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8449 16175 8483
rect 17773 8483 17831 8489
rect 17773 8480 17785 8483
rect 16117 8443 16175 8449
rect 16408 8452 17785 8480
rect 13354 8412 13360 8424
rect 13096 8384 13360 8412
rect 13354 8372 13360 8384
rect 13412 8412 13418 8424
rect 14553 8415 14611 8421
rect 14553 8412 14565 8415
rect 13412 8384 14565 8412
rect 13412 8372 13418 8384
rect 14553 8381 14565 8384
rect 14599 8381 14611 8415
rect 14553 8375 14611 8381
rect 15470 8372 15476 8424
rect 15528 8412 15534 8424
rect 15749 8415 15807 8421
rect 15749 8412 15761 8415
rect 15528 8384 15761 8412
rect 15528 8372 15534 8384
rect 15749 8381 15761 8384
rect 15795 8381 15807 8415
rect 15749 8375 15807 8381
rect 10704 8344 10732 8372
rect 10781 8347 10839 8353
rect 10781 8344 10793 8347
rect 10704 8316 10793 8344
rect 10781 8313 10793 8316
rect 10827 8313 10839 8347
rect 10781 8307 10839 8313
rect 12250 8304 12256 8356
rect 12308 8344 12314 8356
rect 12437 8347 12495 8353
rect 12437 8344 12449 8347
rect 12308 8316 12449 8344
rect 12308 8304 12314 8316
rect 12437 8313 12449 8316
rect 12483 8313 12495 8347
rect 12989 8347 13047 8353
rect 12989 8344 13001 8347
rect 12437 8307 12495 8313
rect 12544 8316 13001 8344
rect 10962 8276 10968 8288
rect 10051 8248 10968 8276
rect 10962 8236 10968 8248
rect 11020 8236 11026 8288
rect 12069 8279 12127 8285
rect 12069 8245 12081 8279
rect 12115 8276 12127 8279
rect 12544 8276 12572 8316
rect 12989 8313 13001 8316
rect 13035 8313 13047 8347
rect 12989 8307 13047 8313
rect 13998 8304 14004 8356
rect 14056 8344 14062 8356
rect 16132 8344 16160 8443
rect 14056 8316 16160 8344
rect 14056 8304 14062 8316
rect 12115 8248 12572 8276
rect 12115 8245 12127 8248
rect 12069 8239 12127 8245
rect 13906 8236 13912 8288
rect 13964 8236 13970 8288
rect 15010 8236 15016 8288
rect 15068 8276 15074 8288
rect 16408 8276 16436 8452
rect 17773 8449 17785 8452
rect 17819 8449 17831 8483
rect 17773 8443 17831 8449
rect 17957 8483 18015 8489
rect 17957 8449 17969 8483
rect 18003 8449 18015 8483
rect 17957 8443 18015 8449
rect 16482 8372 16488 8424
rect 16540 8412 16546 8424
rect 17972 8412 18000 8443
rect 18230 8440 18236 8492
rect 18288 8480 18294 8492
rect 18417 8483 18475 8489
rect 18417 8480 18429 8483
rect 18288 8452 18429 8480
rect 18288 8440 18294 8452
rect 18417 8449 18429 8452
rect 18463 8480 18475 8483
rect 19058 8480 19064 8492
rect 18463 8452 19064 8480
rect 18463 8449 18475 8452
rect 18417 8443 18475 8449
rect 19058 8440 19064 8452
rect 19116 8440 19122 8492
rect 19153 8415 19211 8421
rect 19153 8412 19165 8415
rect 16540 8384 19165 8412
rect 16540 8372 16546 8384
rect 19153 8381 19165 8384
rect 19199 8381 19211 8415
rect 19613 8415 19671 8421
rect 19613 8412 19625 8415
rect 19153 8375 19211 8381
rect 19260 8384 19625 8412
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 18601 8347 18659 8353
rect 18601 8344 18613 8347
rect 16632 8316 18613 8344
rect 16632 8304 16638 8316
rect 18601 8313 18613 8316
rect 18647 8344 18659 8347
rect 18782 8344 18788 8356
rect 18647 8316 18788 8344
rect 18647 8313 18659 8316
rect 18601 8307 18659 8313
rect 18782 8304 18788 8316
rect 18840 8344 18846 8356
rect 19260 8344 19288 8384
rect 19613 8381 19625 8384
rect 19659 8381 19671 8415
rect 19613 8375 19671 8381
rect 18840 8316 19288 8344
rect 18840 8304 18846 8316
rect 19334 8304 19340 8356
rect 19392 8304 19398 8356
rect 15068 8248 16436 8276
rect 15068 8236 15074 8248
rect 1104 8186 22816 8208
rect 1104 8134 3664 8186
rect 3716 8134 3728 8186
rect 3780 8134 3792 8186
rect 3844 8134 3856 8186
rect 3908 8134 3920 8186
rect 3972 8134 9092 8186
rect 9144 8134 9156 8186
rect 9208 8134 9220 8186
rect 9272 8134 9284 8186
rect 9336 8134 9348 8186
rect 9400 8134 14520 8186
rect 14572 8134 14584 8186
rect 14636 8134 14648 8186
rect 14700 8134 14712 8186
rect 14764 8134 14776 8186
rect 14828 8134 19948 8186
rect 20000 8134 20012 8186
rect 20064 8134 20076 8186
rect 20128 8134 20140 8186
rect 20192 8134 20204 8186
rect 20256 8134 22816 8186
rect 1104 8112 22816 8134
rect 3237 8075 3295 8081
rect 3237 8041 3249 8075
rect 3283 8041 3295 8075
rect 3237 8035 3295 8041
rect 3252 8004 3280 8035
rect 3418 8032 3424 8084
rect 3476 8032 3482 8084
rect 3510 8032 3516 8084
rect 3568 8072 3574 8084
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 3568 8044 4077 8072
rect 3568 8032 3574 8044
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 4065 8035 4123 8041
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 4890 8072 4896 8084
rect 4304 8044 4896 8072
rect 4304 8032 4310 8044
rect 4890 8032 4896 8044
rect 4948 8032 4954 8084
rect 7377 8075 7435 8081
rect 7377 8041 7389 8075
rect 7423 8041 7435 8075
rect 7377 8035 7435 8041
rect 3252 7976 4568 8004
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 4433 7871 4491 7877
rect 4433 7868 4445 7871
rect 4212 7840 4445 7868
rect 4212 7828 4218 7840
rect 4433 7837 4445 7840
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 4540 7868 4568 7976
rect 7392 7948 7420 8035
rect 7558 8032 7564 8084
rect 7616 8032 7622 8084
rect 8478 8032 8484 8084
rect 8536 8032 8542 8084
rect 9769 8075 9827 8081
rect 9769 8041 9781 8075
rect 9815 8072 9827 8075
rect 9950 8072 9956 8084
rect 9815 8044 9956 8072
rect 9815 8041 9827 8044
rect 9769 8035 9827 8041
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 10965 8075 11023 8081
rect 10965 8041 10977 8075
rect 11011 8072 11023 8075
rect 13446 8072 13452 8084
rect 11011 8044 13452 8072
rect 11011 8041 11023 8044
rect 10965 8035 11023 8041
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 13633 8075 13691 8081
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 15562 8072 15568 8084
rect 13679 8044 15568 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 15562 8032 15568 8044
rect 15620 8032 15626 8084
rect 15657 8075 15715 8081
rect 15657 8041 15669 8075
rect 15703 8072 15715 8075
rect 16298 8072 16304 8084
rect 15703 8044 16304 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 8389 8007 8447 8013
rect 8389 7973 8401 8007
rect 8435 8004 8447 8007
rect 8662 8004 8668 8016
rect 8435 7976 8668 8004
rect 8435 7973 8447 7976
rect 8389 7967 8447 7973
rect 8662 7964 8668 7976
rect 8720 7964 8726 8016
rect 12158 8004 12164 8016
rect 8772 7976 12164 8004
rect 5074 7896 5080 7948
rect 5132 7936 5138 7948
rect 7009 7939 7067 7945
rect 7009 7936 7021 7939
rect 5132 7908 7021 7936
rect 5132 7896 5138 7908
rect 4706 7868 4712 7880
rect 4540 7840 4712 7868
rect 3053 7803 3111 7809
rect 3053 7769 3065 7803
rect 3099 7769 3111 7803
rect 3053 7763 3111 7769
rect 3269 7803 3327 7809
rect 3269 7769 3281 7803
rect 3315 7800 3327 7803
rect 4246 7800 4252 7812
rect 3315 7772 4252 7800
rect 3315 7769 3327 7772
rect 3269 7763 3327 7769
rect 3068 7732 3096 7763
rect 4246 7760 4252 7772
rect 4304 7760 4310 7812
rect 4341 7803 4399 7809
rect 4341 7769 4353 7803
rect 4387 7800 4399 7803
rect 4540 7800 4568 7840
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 5276 7877 5304 7908
rect 7009 7905 7021 7908
rect 7055 7905 7067 7939
rect 7009 7899 7067 7905
rect 7374 7896 7380 7948
rect 7432 7936 7438 7948
rect 8772 7936 8800 7976
rect 12158 7964 12164 7976
rect 12216 7964 12222 8016
rect 13541 8007 13599 8013
rect 13541 8004 13553 8007
rect 12406 7976 13553 8004
rect 9861 7939 9919 7945
rect 7432 7908 8800 7936
rect 8864 7908 9812 7936
rect 7432 7896 7438 7908
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7837 5319 7871
rect 5261 7831 5319 7837
rect 5442 7828 5448 7880
rect 5500 7828 5506 7880
rect 5534 7828 5540 7880
rect 5592 7828 5598 7880
rect 5902 7828 5908 7880
rect 5960 7868 5966 7880
rect 5997 7871 6055 7877
rect 5997 7868 6009 7871
rect 5960 7840 6009 7868
rect 5960 7828 5966 7840
rect 5997 7837 6009 7840
rect 6043 7837 6055 7871
rect 6273 7871 6331 7877
rect 6273 7868 6285 7871
rect 5997 7831 6055 7837
rect 6104 7840 6285 7868
rect 4387 7772 4568 7800
rect 4617 7803 4675 7809
rect 4387 7769 4399 7772
rect 4341 7763 4399 7769
rect 4617 7769 4629 7803
rect 4663 7800 4675 7803
rect 5460 7800 5488 7828
rect 6104 7800 6132 7840
rect 6273 7837 6285 7840
rect 6319 7837 6331 7871
rect 6273 7831 6331 7837
rect 6362 7828 6368 7880
rect 6420 7868 6426 7880
rect 6420 7840 7052 7868
rect 6420 7828 6426 7840
rect 7024 7812 7052 7840
rect 7926 7828 7932 7880
rect 7984 7868 7990 7880
rect 8021 7871 8079 7877
rect 8021 7868 8033 7871
rect 7984 7840 8033 7868
rect 7984 7828 7990 7840
rect 8021 7837 8033 7840
rect 8067 7868 8079 7871
rect 8864 7868 8892 7908
rect 8067 7840 8892 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 9398 7828 9404 7880
rect 9456 7868 9462 7880
rect 9640 7871 9698 7877
rect 9640 7868 9652 7871
rect 9456 7840 9652 7868
rect 9456 7828 9462 7840
rect 9640 7837 9652 7840
rect 9686 7837 9698 7871
rect 9784 7868 9812 7908
rect 9861 7905 9873 7939
rect 9907 7936 9919 7939
rect 12406 7936 12434 7976
rect 13541 7973 13553 7976
rect 13587 7973 13599 8007
rect 13541 7967 13599 7973
rect 9907 7908 12434 7936
rect 9907 7905 9919 7908
rect 9861 7899 9919 7905
rect 12526 7896 12532 7948
rect 12584 7896 12590 7948
rect 13446 7896 13452 7948
rect 13504 7896 13510 7948
rect 15672 7936 15700 8035
rect 16298 8032 16304 8044
rect 16356 8032 16362 8084
rect 18506 8032 18512 8084
rect 18564 8072 18570 8084
rect 18601 8075 18659 8081
rect 18601 8072 18613 8075
rect 18564 8044 18613 8072
rect 18564 8032 18570 8044
rect 18601 8041 18613 8044
rect 18647 8041 18659 8075
rect 18601 8035 18659 8041
rect 19613 8075 19671 8081
rect 19613 8041 19625 8075
rect 19659 8041 19671 8075
rect 19613 8035 19671 8041
rect 16114 7964 16120 8016
rect 16172 8004 16178 8016
rect 17034 8004 17040 8016
rect 16172 7976 17040 8004
rect 16172 7964 16178 7976
rect 17034 7964 17040 7976
rect 17092 7964 17098 8016
rect 18322 7964 18328 8016
rect 18380 8004 18386 8016
rect 19628 8004 19656 8035
rect 18380 7976 19656 8004
rect 18380 7964 18386 7976
rect 18138 7936 18144 7948
rect 13740 7908 15700 7936
rect 16316 7908 18144 7936
rect 10873 7871 10931 7877
rect 10873 7868 10885 7871
rect 9784 7840 10885 7868
rect 9640 7831 9698 7837
rect 10873 7837 10885 7840
rect 10919 7868 10931 7871
rect 10962 7868 10968 7880
rect 10919 7840 10968 7868
rect 10919 7837 10931 7840
rect 10873 7831 10931 7837
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 11054 7828 11060 7880
rect 11112 7868 11118 7880
rect 13740 7877 13768 7908
rect 11241 7871 11299 7877
rect 11241 7868 11253 7871
rect 11112 7840 11253 7868
rect 11112 7828 11118 7840
rect 11241 7837 11253 7840
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14461 7871 14519 7877
rect 14461 7868 14473 7871
rect 13964 7840 14473 7868
rect 13964 7828 13970 7840
rect 14461 7837 14473 7840
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7868 14611 7871
rect 16114 7868 16120 7880
rect 14599 7840 16120 7868
rect 14599 7837 14611 7840
rect 14553 7831 14611 7837
rect 4663 7772 5396 7800
rect 5460 7772 6132 7800
rect 6181 7803 6239 7809
rect 4663 7769 4675 7772
rect 4617 7763 4675 7769
rect 4632 7732 4660 7763
rect 3068 7704 4660 7732
rect 5074 7692 5080 7744
rect 5132 7692 5138 7744
rect 5368 7732 5396 7772
rect 6181 7769 6193 7803
rect 6227 7769 6239 7803
rect 6730 7800 6736 7812
rect 6181 7763 6239 7769
rect 6380 7772 6736 7800
rect 5534 7732 5540 7744
rect 5368 7704 5540 7732
rect 5534 7692 5540 7704
rect 5592 7692 5598 7744
rect 6196 7732 6224 7763
rect 6380 7732 6408 7772
rect 6730 7760 6736 7772
rect 6788 7760 6794 7812
rect 7006 7760 7012 7812
rect 7064 7760 7070 7812
rect 9490 7760 9496 7812
rect 9548 7760 9554 7812
rect 12253 7803 12311 7809
rect 12253 7800 12265 7803
rect 9600 7772 12265 7800
rect 9600 7744 9628 7772
rect 12253 7769 12265 7772
rect 12299 7769 12311 7803
rect 12253 7763 12311 7769
rect 14274 7760 14280 7812
rect 14332 7760 14338 7812
rect 14366 7760 14372 7812
rect 14424 7800 14430 7812
rect 14568 7800 14596 7831
rect 16114 7828 16120 7840
rect 16172 7868 16178 7880
rect 16316 7877 16344 7908
rect 18138 7896 18144 7908
rect 18196 7896 18202 7948
rect 19518 7896 19524 7948
rect 19576 7936 19582 7948
rect 19576 7908 19840 7936
rect 19576 7896 19582 7908
rect 16301 7871 16359 7877
rect 16301 7868 16313 7871
rect 16172 7840 16313 7868
rect 16172 7828 16178 7840
rect 16301 7837 16313 7840
rect 16347 7837 16359 7871
rect 16301 7831 16359 7837
rect 16482 7828 16488 7880
rect 16540 7828 16546 7880
rect 16942 7828 16948 7880
rect 17000 7828 17006 7880
rect 17034 7828 17040 7880
rect 17092 7868 17098 7880
rect 17129 7871 17187 7877
rect 17129 7868 17141 7871
rect 17092 7840 17141 7868
rect 17092 7828 17098 7840
rect 17129 7837 17141 7840
rect 17175 7837 17187 7871
rect 17129 7831 17187 7837
rect 17405 7871 17463 7877
rect 17405 7837 17417 7871
rect 17451 7837 17463 7871
rect 17405 7831 17463 7837
rect 14424 7772 14596 7800
rect 14645 7803 14703 7809
rect 14424 7760 14430 7772
rect 14645 7769 14657 7803
rect 14691 7769 14703 7803
rect 14645 7763 14703 7769
rect 6196 7704 6408 7732
rect 6549 7735 6607 7741
rect 6549 7701 6561 7735
rect 6595 7732 6607 7735
rect 7377 7735 7435 7741
rect 7377 7732 7389 7735
rect 6595 7704 7389 7732
rect 6595 7701 6607 7704
rect 6549 7695 6607 7701
rect 7377 7701 7389 7704
rect 7423 7701 7435 7735
rect 7377 7695 7435 7701
rect 9582 7692 9588 7744
rect 9640 7692 9646 7744
rect 10137 7735 10195 7741
rect 10137 7701 10149 7735
rect 10183 7732 10195 7735
rect 10594 7732 10600 7744
rect 10183 7704 10600 7732
rect 10183 7701 10195 7704
rect 10137 7695 10195 7701
rect 10594 7692 10600 7704
rect 10652 7692 10658 7744
rect 10686 7692 10692 7744
rect 10744 7692 10750 7744
rect 12342 7692 12348 7744
rect 12400 7732 12406 7744
rect 12526 7732 12532 7744
rect 12400 7704 12532 7732
rect 12400 7692 12406 7704
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 14660 7732 14688 7763
rect 15010 7760 15016 7812
rect 15068 7760 15074 7812
rect 15102 7760 15108 7812
rect 15160 7800 15166 7812
rect 15841 7803 15899 7809
rect 15841 7800 15853 7803
rect 15160 7772 15853 7800
rect 15160 7760 15166 7772
rect 15841 7769 15853 7772
rect 15887 7769 15899 7803
rect 16500 7800 16528 7828
rect 15841 7763 15899 7769
rect 15948 7772 16528 7800
rect 14918 7732 14924 7744
rect 14660 7704 14924 7732
rect 14918 7692 14924 7704
rect 14976 7732 14982 7744
rect 15473 7735 15531 7741
rect 15473 7732 15485 7735
rect 14976 7704 15485 7732
rect 14976 7692 14982 7704
rect 15473 7701 15485 7704
rect 15519 7701 15531 7735
rect 15473 7695 15531 7701
rect 15641 7735 15699 7741
rect 15641 7701 15653 7735
rect 15687 7732 15699 7735
rect 15948 7732 15976 7772
rect 16574 7760 16580 7812
rect 16632 7800 16638 7812
rect 17420 7800 17448 7831
rect 18046 7828 18052 7880
rect 18104 7828 18110 7880
rect 18414 7828 18420 7880
rect 18472 7828 18478 7880
rect 18782 7828 18788 7880
rect 18840 7868 18846 7880
rect 19812 7877 19840 7908
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 18840 7840 19625 7868
rect 18840 7828 18846 7840
rect 19613 7837 19625 7840
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 19797 7871 19855 7877
rect 19797 7837 19809 7871
rect 19843 7837 19855 7871
rect 19797 7831 19855 7837
rect 16632 7772 17448 7800
rect 17589 7803 17647 7809
rect 16632 7760 16638 7772
rect 17589 7769 17601 7803
rect 17635 7800 17647 7803
rect 18233 7803 18291 7809
rect 18233 7800 18245 7803
rect 17635 7772 18245 7800
rect 17635 7769 17647 7772
rect 17589 7763 17647 7769
rect 18233 7769 18245 7772
rect 18279 7769 18291 7803
rect 18233 7763 18291 7769
rect 18325 7803 18383 7809
rect 18325 7769 18337 7803
rect 18371 7800 18383 7803
rect 18371 7772 19472 7800
rect 18371 7769 18383 7772
rect 18325 7763 18383 7769
rect 15687 7704 15976 7732
rect 15687 7701 15699 7704
rect 15641 7695 15699 7701
rect 16022 7692 16028 7744
rect 16080 7732 16086 7744
rect 19444 7741 19472 7772
rect 16301 7735 16359 7741
rect 16301 7732 16313 7735
rect 16080 7704 16313 7732
rect 16080 7692 16086 7704
rect 16301 7701 16313 7704
rect 16347 7701 16359 7735
rect 16301 7695 16359 7701
rect 19429 7735 19487 7741
rect 19429 7701 19441 7735
rect 19475 7701 19487 7735
rect 19429 7695 19487 7701
rect 1104 7642 22976 7664
rect 1104 7590 6378 7642
rect 6430 7590 6442 7642
rect 6494 7590 6506 7642
rect 6558 7590 6570 7642
rect 6622 7590 6634 7642
rect 6686 7590 11806 7642
rect 11858 7590 11870 7642
rect 11922 7590 11934 7642
rect 11986 7590 11998 7642
rect 12050 7590 12062 7642
rect 12114 7590 17234 7642
rect 17286 7590 17298 7642
rect 17350 7590 17362 7642
rect 17414 7590 17426 7642
rect 17478 7590 17490 7642
rect 17542 7590 22662 7642
rect 22714 7590 22726 7642
rect 22778 7590 22790 7642
rect 22842 7590 22854 7642
rect 22906 7590 22918 7642
rect 22970 7590 22976 7642
rect 1104 7568 22976 7590
rect 4433 7531 4491 7537
rect 4433 7497 4445 7531
rect 4479 7528 4491 7531
rect 4522 7528 4528 7540
rect 4479 7500 4528 7528
rect 4479 7497 4491 7500
rect 4433 7491 4491 7497
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 4890 7488 4896 7540
rect 4948 7528 4954 7540
rect 6549 7531 6607 7537
rect 6549 7528 6561 7531
rect 4948 7500 6561 7528
rect 4948 7488 4954 7500
rect 6549 7497 6561 7500
rect 6595 7497 6607 7531
rect 6549 7491 6607 7497
rect 6914 7488 6920 7540
rect 6972 7528 6978 7540
rect 7377 7531 7435 7537
rect 7377 7528 7389 7531
rect 6972 7500 7389 7528
rect 6972 7488 6978 7500
rect 7377 7497 7389 7500
rect 7423 7497 7435 7531
rect 7377 7491 7435 7497
rect 9398 7488 9404 7540
rect 9456 7488 9462 7540
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 10137 7531 10195 7537
rect 10137 7528 10149 7531
rect 10100 7500 10149 7528
rect 10100 7488 10106 7500
rect 10137 7497 10149 7500
rect 10183 7497 10195 7531
rect 10137 7491 10195 7497
rect 10594 7488 10600 7540
rect 10652 7528 10658 7540
rect 17589 7531 17647 7537
rect 10652 7500 13400 7528
rect 10652 7488 10658 7500
rect 4249 7463 4307 7469
rect 4249 7429 4261 7463
rect 4295 7460 4307 7463
rect 4338 7460 4344 7472
rect 4295 7432 4344 7460
rect 4295 7429 4307 7432
rect 4249 7423 4307 7429
rect 4338 7420 4344 7432
rect 4396 7460 4402 7472
rect 7282 7460 7288 7472
rect 4396 7432 7288 7460
rect 4396 7420 4402 7432
rect 7282 7420 7288 7432
rect 7340 7420 7346 7472
rect 8478 7460 8484 7472
rect 7668 7432 8484 7460
rect 3418 7352 3424 7404
rect 3476 7392 3482 7404
rect 3881 7395 3939 7401
rect 3881 7392 3893 7395
rect 3476 7364 3893 7392
rect 3476 7352 3482 7364
rect 3881 7361 3893 7364
rect 3927 7361 3939 7395
rect 3881 7355 3939 7361
rect 6730 7352 6736 7404
rect 6788 7392 6794 7404
rect 7668 7401 7696 7432
rect 8478 7420 8484 7432
rect 8536 7420 8542 7472
rect 10321 7463 10379 7469
rect 10321 7429 10333 7463
rect 10367 7460 10379 7463
rect 11701 7463 11759 7469
rect 11701 7460 11713 7463
rect 10367 7432 11713 7460
rect 10367 7429 10379 7432
rect 10321 7423 10379 7429
rect 11701 7429 11713 7432
rect 11747 7429 11759 7463
rect 12069 7463 12127 7469
rect 11701 7423 11759 7429
rect 11808 7432 12020 7460
rect 7653 7395 7711 7401
rect 7653 7392 7665 7395
rect 6788 7364 7665 7392
rect 6788 7352 6794 7364
rect 7653 7361 7665 7364
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 7926 7352 7932 7404
rect 7984 7392 7990 7404
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 7984 7364 8125 7392
rect 7984 7352 7990 7364
rect 8113 7361 8125 7364
rect 8159 7392 8171 7395
rect 8941 7395 8999 7401
rect 8941 7392 8953 7395
rect 8159 7364 8953 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 8941 7361 8953 7364
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7392 9459 7395
rect 10686 7392 10692 7404
rect 9447 7364 10692 7392
rect 9447 7361 9459 7364
rect 9401 7355 9459 7361
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 11146 7352 11152 7404
rect 11204 7392 11210 7404
rect 11808 7392 11836 7432
rect 11204 7364 11836 7392
rect 11885 7395 11943 7401
rect 11204 7352 11210 7364
rect 11885 7361 11897 7395
rect 11931 7361 11943 7395
rect 11992 7392 12020 7432
rect 12069 7429 12081 7463
rect 12115 7460 12127 7463
rect 12342 7460 12348 7472
rect 12115 7432 12348 7460
rect 12115 7429 12127 7432
rect 12069 7423 12127 7429
rect 12342 7420 12348 7432
rect 12400 7420 12406 7472
rect 13372 7460 13400 7500
rect 13740 7500 17540 7528
rect 13740 7460 13768 7500
rect 13372 7432 13768 7460
rect 13906 7420 13912 7472
rect 13964 7460 13970 7472
rect 13964 7432 14872 7460
rect 13964 7420 13970 7432
rect 12161 7395 12219 7401
rect 12161 7392 12173 7395
rect 11992 7364 12173 7392
rect 11885 7355 11943 7361
rect 12161 7361 12173 7364
rect 12207 7392 12219 7395
rect 14274 7392 14280 7404
rect 12207 7364 14280 7392
rect 12207 7361 12219 7364
rect 12161 7355 12219 7361
rect 6917 7327 6975 7333
rect 6917 7293 6929 7327
rect 6963 7324 6975 7327
rect 7006 7324 7012 7336
rect 6963 7296 7012 7324
rect 6963 7293 6975 7296
rect 6917 7287 6975 7293
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 7374 7284 7380 7336
rect 7432 7284 7438 7336
rect 7466 7284 7472 7336
rect 7524 7324 7530 7336
rect 7561 7327 7619 7333
rect 7561 7324 7573 7327
rect 7524 7296 7573 7324
rect 7524 7284 7530 7296
rect 7561 7293 7573 7296
rect 7607 7324 7619 7327
rect 11900 7324 11928 7355
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 12250 7324 12256 7336
rect 7607 7296 10732 7324
rect 11900 7296 12256 7324
rect 7607 7293 7619 7296
rect 7561 7287 7619 7293
rect 5074 7256 5080 7268
rect 4264 7228 5080 7256
rect 4264 7197 4292 7228
rect 5074 7216 5080 7228
rect 5132 7216 5138 7268
rect 8205 7259 8263 7265
rect 8205 7225 8217 7259
rect 8251 7256 8263 7259
rect 9582 7256 9588 7268
rect 8251 7228 9588 7256
rect 8251 7225 8263 7228
rect 8205 7219 8263 7225
rect 9582 7216 9588 7228
rect 9640 7216 9646 7268
rect 10704 7265 10732 7296
rect 12250 7284 12256 7296
rect 12308 7284 12314 7336
rect 13998 7284 14004 7336
rect 14056 7284 14062 7336
rect 14844 7324 14872 7432
rect 15838 7420 15844 7472
rect 15896 7460 15902 7472
rect 15993 7463 16051 7469
rect 15993 7460 16005 7463
rect 15896 7432 16005 7460
rect 15896 7420 15902 7432
rect 15993 7429 16005 7432
rect 16039 7429 16051 7463
rect 15993 7423 16051 7429
rect 16209 7463 16267 7469
rect 16209 7429 16221 7463
rect 16255 7460 16267 7463
rect 16390 7460 16396 7472
rect 16255 7432 16396 7460
rect 16255 7429 16267 7432
rect 16209 7423 16267 7429
rect 16390 7420 16396 7432
rect 16448 7420 16454 7472
rect 16942 7420 16948 7472
rect 17000 7460 17006 7472
rect 17512 7460 17540 7500
rect 17589 7497 17601 7531
rect 17635 7528 17647 7531
rect 18046 7528 18052 7540
rect 17635 7500 18052 7528
rect 17635 7497 17647 7500
rect 17589 7491 17647 7497
rect 18046 7488 18052 7500
rect 18104 7488 18110 7540
rect 18414 7488 18420 7540
rect 18472 7488 18478 7540
rect 19242 7528 19248 7540
rect 18616 7500 19248 7528
rect 18616 7460 18644 7500
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 19518 7460 19524 7472
rect 17000 7432 17448 7460
rect 17512 7432 18644 7460
rect 18708 7432 19524 7460
rect 17000 7420 17006 7432
rect 16574 7352 16580 7404
rect 16632 7392 16638 7404
rect 17420 7401 17448 7432
rect 17221 7395 17279 7401
rect 17221 7392 17233 7395
rect 16632 7364 17233 7392
rect 16632 7352 16638 7364
rect 17221 7361 17233 7364
rect 17267 7361 17279 7395
rect 17221 7355 17279 7361
rect 17313 7395 17371 7401
rect 17313 7361 17325 7395
rect 17359 7361 17371 7395
rect 17313 7355 17371 7361
rect 17405 7395 17463 7401
rect 17405 7361 17417 7395
rect 17451 7361 17463 7395
rect 17405 7355 17463 7361
rect 14844 7296 15884 7324
rect 10689 7259 10747 7265
rect 10689 7225 10701 7259
rect 10735 7256 10747 7259
rect 15010 7256 15016 7268
rect 10735 7228 15016 7256
rect 10735 7225 10747 7228
rect 10689 7219 10747 7225
rect 15010 7216 15016 7228
rect 15068 7216 15074 7268
rect 15856 7265 15884 7296
rect 17034 7284 17040 7336
rect 17092 7324 17098 7336
rect 17328 7324 17356 7355
rect 18322 7352 18328 7404
rect 18380 7392 18386 7404
rect 18708 7401 18736 7432
rect 19518 7420 19524 7432
rect 19576 7420 19582 7472
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 18380 7364 18613 7392
rect 18380 7352 18386 7364
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 18693 7395 18751 7401
rect 18693 7361 18705 7395
rect 18739 7361 18751 7395
rect 18693 7355 18751 7361
rect 18782 7352 18788 7404
rect 18840 7352 18846 7404
rect 17092 7296 17356 7324
rect 17092 7284 17098 7296
rect 15841 7259 15899 7265
rect 15841 7225 15853 7259
rect 15887 7225 15899 7259
rect 15841 7219 15899 7225
rect 4249 7191 4307 7197
rect 4249 7157 4261 7191
rect 4295 7157 4307 7191
rect 4249 7151 4307 7157
rect 8662 7148 8668 7200
rect 8720 7188 8726 7200
rect 9079 7191 9137 7197
rect 9079 7188 9091 7191
rect 8720 7160 9091 7188
rect 8720 7148 8726 7160
rect 9079 7157 9091 7160
rect 9125 7157 9137 7191
rect 9079 7151 9137 7157
rect 9214 7148 9220 7200
rect 9272 7148 9278 7200
rect 10321 7191 10379 7197
rect 10321 7157 10333 7191
rect 10367 7188 10379 7191
rect 12158 7188 12164 7200
rect 10367 7160 12164 7188
rect 10367 7157 10379 7160
rect 10321 7151 10379 7157
rect 12158 7148 12164 7160
rect 12216 7148 12222 7200
rect 13446 7148 13452 7200
rect 13504 7188 13510 7200
rect 13725 7191 13783 7197
rect 13725 7188 13737 7191
rect 13504 7160 13737 7188
rect 13504 7148 13510 7160
rect 13725 7157 13737 7160
rect 13771 7157 13783 7191
rect 13725 7151 13783 7157
rect 14185 7191 14243 7197
rect 14185 7157 14197 7191
rect 14231 7188 14243 7191
rect 15286 7188 15292 7200
rect 14231 7160 15292 7188
rect 14231 7157 14243 7160
rect 14185 7151 14243 7157
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 16022 7148 16028 7200
rect 16080 7148 16086 7200
rect 1104 7098 22816 7120
rect 1104 7046 3664 7098
rect 3716 7046 3728 7098
rect 3780 7046 3792 7098
rect 3844 7046 3856 7098
rect 3908 7046 3920 7098
rect 3972 7046 9092 7098
rect 9144 7046 9156 7098
rect 9208 7046 9220 7098
rect 9272 7046 9284 7098
rect 9336 7046 9348 7098
rect 9400 7046 14520 7098
rect 14572 7046 14584 7098
rect 14636 7046 14648 7098
rect 14700 7046 14712 7098
rect 14764 7046 14776 7098
rect 14828 7046 19948 7098
rect 20000 7046 20012 7098
rect 20064 7046 20076 7098
rect 20128 7046 20140 7098
rect 20192 7046 20204 7098
rect 20256 7046 22816 7098
rect 1104 7024 22816 7046
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 9766 6984 9772 6996
rect 5592 6956 9772 6984
rect 5592 6944 5598 6956
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 15838 6944 15844 6996
rect 15896 6944 15902 6996
rect 10962 6876 10968 6928
rect 11020 6916 11026 6928
rect 18230 6916 18236 6928
rect 11020 6888 18236 6916
rect 11020 6876 11026 6888
rect 18230 6876 18236 6888
rect 18288 6876 18294 6928
rect 16025 6783 16083 6789
rect 16025 6749 16037 6783
rect 16071 6780 16083 6783
rect 16114 6780 16120 6792
rect 16071 6752 16120 6780
rect 16071 6749 16083 6752
rect 16025 6743 16083 6749
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6780 16267 6783
rect 16482 6780 16488 6792
rect 16255 6752 16488 6780
rect 16255 6749 16267 6752
rect 16209 6743 16267 6749
rect 16482 6740 16488 6752
rect 16540 6740 16546 6792
rect 1104 6554 22976 6576
rect 1104 6502 6378 6554
rect 6430 6502 6442 6554
rect 6494 6502 6506 6554
rect 6558 6502 6570 6554
rect 6622 6502 6634 6554
rect 6686 6502 11806 6554
rect 11858 6502 11870 6554
rect 11922 6502 11934 6554
rect 11986 6502 11998 6554
rect 12050 6502 12062 6554
rect 12114 6502 17234 6554
rect 17286 6502 17298 6554
rect 17350 6502 17362 6554
rect 17414 6502 17426 6554
rect 17478 6502 17490 6554
rect 17542 6502 22662 6554
rect 22714 6502 22726 6554
rect 22778 6502 22790 6554
rect 22842 6502 22854 6554
rect 22906 6502 22918 6554
rect 22970 6502 22976 6554
rect 1104 6480 22976 6502
rect 1104 6010 22816 6032
rect 1104 5958 3664 6010
rect 3716 5958 3728 6010
rect 3780 5958 3792 6010
rect 3844 5958 3856 6010
rect 3908 5958 3920 6010
rect 3972 5958 9092 6010
rect 9144 5958 9156 6010
rect 9208 5958 9220 6010
rect 9272 5958 9284 6010
rect 9336 5958 9348 6010
rect 9400 5958 14520 6010
rect 14572 5958 14584 6010
rect 14636 5958 14648 6010
rect 14700 5958 14712 6010
rect 14764 5958 14776 6010
rect 14828 5958 19948 6010
rect 20000 5958 20012 6010
rect 20064 5958 20076 6010
rect 20128 5958 20140 6010
rect 20192 5958 20204 6010
rect 20256 5958 22816 6010
rect 1104 5936 22816 5958
rect 1104 5466 22976 5488
rect 1104 5414 6378 5466
rect 6430 5414 6442 5466
rect 6494 5414 6506 5466
rect 6558 5414 6570 5466
rect 6622 5414 6634 5466
rect 6686 5414 11806 5466
rect 11858 5414 11870 5466
rect 11922 5414 11934 5466
rect 11986 5414 11998 5466
rect 12050 5414 12062 5466
rect 12114 5414 17234 5466
rect 17286 5414 17298 5466
rect 17350 5414 17362 5466
rect 17414 5414 17426 5466
rect 17478 5414 17490 5466
rect 17542 5414 22662 5466
rect 22714 5414 22726 5466
rect 22778 5414 22790 5466
rect 22842 5414 22854 5466
rect 22906 5414 22918 5466
rect 22970 5414 22976 5466
rect 1104 5392 22976 5414
rect 1104 4922 22816 4944
rect 1104 4870 3664 4922
rect 3716 4870 3728 4922
rect 3780 4870 3792 4922
rect 3844 4870 3856 4922
rect 3908 4870 3920 4922
rect 3972 4870 9092 4922
rect 9144 4870 9156 4922
rect 9208 4870 9220 4922
rect 9272 4870 9284 4922
rect 9336 4870 9348 4922
rect 9400 4870 14520 4922
rect 14572 4870 14584 4922
rect 14636 4870 14648 4922
rect 14700 4870 14712 4922
rect 14764 4870 14776 4922
rect 14828 4870 19948 4922
rect 20000 4870 20012 4922
rect 20064 4870 20076 4922
rect 20128 4870 20140 4922
rect 20192 4870 20204 4922
rect 20256 4870 22816 4922
rect 1104 4848 22816 4870
rect 1104 4378 22976 4400
rect 1104 4326 6378 4378
rect 6430 4326 6442 4378
rect 6494 4326 6506 4378
rect 6558 4326 6570 4378
rect 6622 4326 6634 4378
rect 6686 4326 11806 4378
rect 11858 4326 11870 4378
rect 11922 4326 11934 4378
rect 11986 4326 11998 4378
rect 12050 4326 12062 4378
rect 12114 4326 17234 4378
rect 17286 4326 17298 4378
rect 17350 4326 17362 4378
rect 17414 4326 17426 4378
rect 17478 4326 17490 4378
rect 17542 4326 22662 4378
rect 22714 4326 22726 4378
rect 22778 4326 22790 4378
rect 22842 4326 22854 4378
rect 22906 4326 22918 4378
rect 22970 4326 22976 4378
rect 1104 4304 22976 4326
rect 1104 3834 22816 3856
rect 1104 3782 3664 3834
rect 3716 3782 3728 3834
rect 3780 3782 3792 3834
rect 3844 3782 3856 3834
rect 3908 3782 3920 3834
rect 3972 3782 9092 3834
rect 9144 3782 9156 3834
rect 9208 3782 9220 3834
rect 9272 3782 9284 3834
rect 9336 3782 9348 3834
rect 9400 3782 14520 3834
rect 14572 3782 14584 3834
rect 14636 3782 14648 3834
rect 14700 3782 14712 3834
rect 14764 3782 14776 3834
rect 14828 3782 19948 3834
rect 20000 3782 20012 3834
rect 20064 3782 20076 3834
rect 20128 3782 20140 3834
rect 20192 3782 20204 3834
rect 20256 3782 22816 3834
rect 1104 3760 22816 3782
rect 1104 3290 22976 3312
rect 1104 3238 6378 3290
rect 6430 3238 6442 3290
rect 6494 3238 6506 3290
rect 6558 3238 6570 3290
rect 6622 3238 6634 3290
rect 6686 3238 11806 3290
rect 11858 3238 11870 3290
rect 11922 3238 11934 3290
rect 11986 3238 11998 3290
rect 12050 3238 12062 3290
rect 12114 3238 17234 3290
rect 17286 3238 17298 3290
rect 17350 3238 17362 3290
rect 17414 3238 17426 3290
rect 17478 3238 17490 3290
rect 17542 3238 22662 3290
rect 22714 3238 22726 3290
rect 22778 3238 22790 3290
rect 22842 3238 22854 3290
rect 22906 3238 22918 3290
rect 22970 3238 22976 3290
rect 1104 3216 22976 3238
rect 1104 2746 22816 2768
rect 1104 2694 3664 2746
rect 3716 2694 3728 2746
rect 3780 2694 3792 2746
rect 3844 2694 3856 2746
rect 3908 2694 3920 2746
rect 3972 2694 9092 2746
rect 9144 2694 9156 2746
rect 9208 2694 9220 2746
rect 9272 2694 9284 2746
rect 9336 2694 9348 2746
rect 9400 2694 14520 2746
rect 14572 2694 14584 2746
rect 14636 2694 14648 2746
rect 14700 2694 14712 2746
rect 14764 2694 14776 2746
rect 14828 2694 19948 2746
rect 20000 2694 20012 2746
rect 20064 2694 20076 2746
rect 20128 2694 20140 2746
rect 20192 2694 20204 2746
rect 20256 2694 22816 2746
rect 1104 2672 22816 2694
rect 10870 2592 10876 2644
rect 10928 2632 10934 2644
rect 10928 2604 16574 2632
rect 10928 2592 10934 2604
rect 6086 2524 6092 2576
rect 6144 2564 6150 2576
rect 6144 2536 14412 2564
rect 6144 2524 6150 2536
rect 8846 2456 8852 2508
rect 8904 2496 8910 2508
rect 8904 2468 14320 2496
rect 8904 2456 8910 2468
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2428 2283 2431
rect 4982 2428 4988 2440
rect 2271 2400 4988 2428
rect 2271 2397 2283 2400
rect 2225 2391 2283 2397
rect 4982 2388 4988 2400
rect 5040 2388 5046 2440
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2428 5227 2431
rect 5902 2428 5908 2440
rect 5215 2400 5908 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 5902 2388 5908 2400
rect 5960 2388 5966 2440
rect 8113 2431 8171 2437
rect 8113 2397 8125 2431
rect 8159 2428 8171 2431
rect 8386 2428 8392 2440
rect 8159 2400 8392 2428
rect 8159 2397 8171 2400
rect 8113 2391 8171 2397
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 8570 2388 8576 2440
rect 8628 2428 8634 2440
rect 14292 2437 14320 2468
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 8628 2400 10609 2428
rect 8628 2388 8634 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 14277 2431 14335 2437
rect 14277 2397 14289 2431
rect 14323 2397 14335 2431
rect 14384 2428 14412 2536
rect 16546 2496 16574 2604
rect 16546 2468 19472 2496
rect 19444 2437 19472 2468
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 14384 2400 16865 2428
rect 14277 2391 14335 2397
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 20990 2388 20996 2440
rect 21048 2388 21054 2440
rect 1670 2320 1676 2372
rect 1728 2360 1734 2372
rect 1949 2363 2007 2369
rect 1949 2360 1961 2363
rect 1728 2332 1961 2360
rect 1728 2320 1734 2332
rect 1949 2329 1961 2332
rect 1995 2329 2007 2363
rect 1949 2323 2007 2329
rect 4614 2320 4620 2372
rect 4672 2360 4678 2372
rect 4893 2363 4951 2369
rect 4893 2360 4905 2363
rect 4672 2332 4905 2360
rect 4672 2320 4678 2332
rect 4893 2329 4905 2332
rect 4939 2329 4951 2363
rect 4893 2323 4951 2329
rect 7558 2320 7564 2372
rect 7616 2360 7622 2372
rect 7837 2363 7895 2369
rect 7837 2360 7849 2363
rect 7616 2332 7849 2360
rect 7616 2320 7622 2332
rect 7837 2329 7849 2332
rect 7883 2329 7895 2363
rect 7837 2323 7895 2329
rect 10502 2320 10508 2372
rect 10560 2360 10566 2372
rect 10873 2363 10931 2369
rect 10873 2360 10885 2363
rect 10560 2332 10885 2360
rect 10560 2320 10566 2332
rect 10873 2329 10885 2332
rect 10919 2329 10931 2363
rect 10873 2323 10931 2329
rect 13814 2320 13820 2372
rect 13872 2360 13878 2372
rect 14553 2363 14611 2369
rect 14553 2360 14565 2363
rect 13872 2332 14565 2360
rect 13872 2320 13878 2332
rect 14553 2329 14565 2332
rect 14599 2329 14611 2363
rect 14553 2323 14611 2329
rect 16574 2320 16580 2372
rect 16632 2360 16638 2372
rect 17129 2363 17187 2369
rect 17129 2360 17141 2363
rect 16632 2332 17141 2360
rect 16632 2320 16638 2332
rect 17129 2329 17141 2332
rect 17175 2329 17187 2363
rect 17129 2323 17187 2329
rect 19334 2320 19340 2372
rect 19392 2360 19398 2372
rect 19705 2363 19763 2369
rect 19705 2360 19717 2363
rect 19392 2332 19717 2360
rect 19392 2320 19398 2332
rect 19705 2329 19717 2332
rect 19751 2329 19763 2363
rect 19705 2323 19763 2329
rect 21269 2363 21327 2369
rect 21269 2329 21281 2363
rect 21315 2360 21327 2363
rect 22278 2360 22284 2372
rect 21315 2332 22284 2360
rect 21315 2329 21327 2332
rect 21269 2323 21327 2329
rect 22278 2320 22284 2332
rect 22336 2320 22342 2372
rect 1104 2202 22976 2224
rect 1104 2150 6378 2202
rect 6430 2150 6442 2202
rect 6494 2150 6506 2202
rect 6558 2150 6570 2202
rect 6622 2150 6634 2202
rect 6686 2150 11806 2202
rect 11858 2150 11870 2202
rect 11922 2150 11934 2202
rect 11986 2150 11998 2202
rect 12050 2150 12062 2202
rect 12114 2150 17234 2202
rect 17286 2150 17298 2202
rect 17350 2150 17362 2202
rect 17414 2150 17426 2202
rect 17478 2150 17490 2202
rect 17542 2150 22662 2202
rect 22714 2150 22726 2202
rect 22778 2150 22790 2202
rect 22842 2150 22854 2202
rect 22906 2150 22918 2202
rect 22970 2150 22976 2202
rect 1104 2128 22976 2150
<< via1 >>
rect 6378 21734 6430 21786
rect 6442 21734 6494 21786
rect 6506 21734 6558 21786
rect 6570 21734 6622 21786
rect 6634 21734 6686 21786
rect 11806 21734 11858 21786
rect 11870 21734 11922 21786
rect 11934 21734 11986 21786
rect 11998 21734 12050 21786
rect 12062 21734 12114 21786
rect 17234 21734 17286 21786
rect 17298 21734 17350 21786
rect 17362 21734 17414 21786
rect 17426 21734 17478 21786
rect 17490 21734 17542 21786
rect 22662 21734 22714 21786
rect 22726 21734 22778 21786
rect 22790 21734 22842 21786
rect 22854 21734 22906 21786
rect 22918 21734 22970 21786
rect 12164 21607 12216 21616
rect 12164 21573 12173 21607
rect 12173 21573 12207 21607
rect 12207 21573 12216 21607
rect 12164 21564 12216 21573
rect 16488 21564 16540 21616
rect 19984 21564 20036 21616
rect 16396 21496 16448 21548
rect 16120 21428 16172 21480
rect 15384 21360 15436 21412
rect 17132 21360 17184 21412
rect 19708 21428 19760 21480
rect 1860 21292 1912 21344
rect 10232 21292 10284 21344
rect 15936 21292 15988 21344
rect 19432 21335 19484 21344
rect 19432 21301 19441 21335
rect 19441 21301 19475 21335
rect 19475 21301 19484 21335
rect 19432 21292 19484 21301
rect 19800 21292 19852 21344
rect 20352 21335 20404 21344
rect 20352 21301 20361 21335
rect 20361 21301 20395 21335
rect 20395 21301 20404 21335
rect 20352 21292 20404 21301
rect 3664 21190 3716 21242
rect 3728 21190 3780 21242
rect 3792 21190 3844 21242
rect 3856 21190 3908 21242
rect 3920 21190 3972 21242
rect 9092 21190 9144 21242
rect 9156 21190 9208 21242
rect 9220 21190 9272 21242
rect 9284 21190 9336 21242
rect 9348 21190 9400 21242
rect 14520 21190 14572 21242
rect 14584 21190 14636 21242
rect 14648 21190 14700 21242
rect 14712 21190 14764 21242
rect 14776 21190 14828 21242
rect 19948 21190 20000 21242
rect 20012 21190 20064 21242
rect 20076 21190 20128 21242
rect 20140 21190 20192 21242
rect 20204 21190 20256 21242
rect 2964 20952 3016 21004
rect 2688 20816 2740 20868
rect 2964 20859 3016 20868
rect 2964 20825 2973 20859
rect 2973 20825 3007 20859
rect 3007 20825 3016 20859
rect 2964 20816 3016 20825
rect 4252 20816 4304 20868
rect 6000 20884 6052 20936
rect 7012 20884 7064 20936
rect 3976 20748 4028 20800
rect 6920 20748 6972 20800
rect 16396 21088 16448 21140
rect 17224 21088 17276 21140
rect 10232 21063 10284 21072
rect 10232 21029 10241 21063
rect 10241 21029 10275 21063
rect 10275 21029 10284 21063
rect 10232 21020 10284 21029
rect 13820 21020 13872 21072
rect 12164 20884 12216 20936
rect 15476 20927 15528 20936
rect 15476 20893 15485 20927
rect 15485 20893 15519 20927
rect 15519 20893 15528 20927
rect 15476 20884 15528 20893
rect 9128 20859 9180 20868
rect 9128 20825 9137 20859
rect 9137 20825 9171 20859
rect 9171 20825 9180 20859
rect 9128 20816 9180 20825
rect 9312 20859 9364 20868
rect 9312 20825 9321 20859
rect 9321 20825 9355 20859
rect 9355 20825 9364 20859
rect 9312 20816 9364 20825
rect 16028 20816 16080 20868
rect 16304 20927 16356 20936
rect 16304 20893 16313 20927
rect 16313 20893 16347 20927
rect 16347 20893 16356 20927
rect 16304 20884 16356 20893
rect 16488 20884 16540 20936
rect 17316 21063 17368 21072
rect 17316 21029 17325 21063
rect 17325 21029 17359 21063
rect 17359 21029 17368 21063
rect 17316 21020 17368 21029
rect 17960 20995 18012 21004
rect 17960 20961 17969 20995
rect 17969 20961 18003 20995
rect 18003 20961 18012 20995
rect 17960 20952 18012 20961
rect 17224 20816 17276 20868
rect 18236 20927 18288 20936
rect 18236 20893 18245 20927
rect 18245 20893 18279 20927
rect 18279 20893 18288 20927
rect 18236 20884 18288 20893
rect 19708 20927 19760 20936
rect 19708 20893 19717 20927
rect 19717 20893 19751 20927
rect 19751 20893 19760 20927
rect 19708 20884 19760 20893
rect 19892 20884 19944 20936
rect 20444 20816 20496 20868
rect 9956 20748 10008 20800
rect 16488 20748 16540 20800
rect 18696 20748 18748 20800
rect 18788 20748 18840 20800
rect 6378 20646 6430 20698
rect 6442 20646 6494 20698
rect 6506 20646 6558 20698
rect 6570 20646 6622 20698
rect 6634 20646 6686 20698
rect 11806 20646 11858 20698
rect 11870 20646 11922 20698
rect 11934 20646 11986 20698
rect 11998 20646 12050 20698
rect 12062 20646 12114 20698
rect 17234 20646 17286 20698
rect 17298 20646 17350 20698
rect 17362 20646 17414 20698
rect 17426 20646 17478 20698
rect 17490 20646 17542 20698
rect 22662 20646 22714 20698
rect 22726 20646 22778 20698
rect 22790 20646 22842 20698
rect 22854 20646 22906 20698
rect 22918 20646 22970 20698
rect 1860 20587 1912 20596
rect 1860 20553 1869 20587
rect 1869 20553 1903 20587
rect 1903 20553 1912 20587
rect 1860 20544 1912 20553
rect 2964 20544 3016 20596
rect 4252 20544 4304 20596
rect 9128 20544 9180 20596
rect 13820 20587 13872 20596
rect 13820 20553 13829 20587
rect 13829 20553 13863 20587
rect 13863 20553 13872 20587
rect 13820 20544 13872 20553
rect 17960 20544 18012 20596
rect 18236 20544 18288 20596
rect 1768 20451 1820 20460
rect 1768 20417 1777 20451
rect 1777 20417 1811 20451
rect 1811 20417 1820 20451
rect 1768 20408 1820 20417
rect 6920 20476 6972 20528
rect 9956 20519 10008 20528
rect 9956 20485 9990 20519
rect 9990 20485 10008 20519
rect 9956 20476 10008 20485
rect 3056 20408 3108 20460
rect 7012 20451 7064 20460
rect 7012 20417 7021 20451
rect 7021 20417 7055 20451
rect 7055 20417 7064 20451
rect 7012 20408 7064 20417
rect 6000 20340 6052 20392
rect 9312 20408 9364 20460
rect 14372 20408 14424 20460
rect 15384 20408 15436 20460
rect 15936 20451 15988 20460
rect 15936 20417 15945 20451
rect 15945 20417 15979 20451
rect 15979 20417 15988 20451
rect 15936 20408 15988 20417
rect 16488 20408 16540 20460
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 17224 20451 17276 20460
rect 17224 20417 17233 20451
rect 17233 20417 17267 20451
rect 17267 20417 17276 20451
rect 17224 20408 17276 20417
rect 20444 20476 20496 20528
rect 19432 20408 19484 20460
rect 2688 20272 2740 20324
rect 2228 20204 2280 20256
rect 2872 20247 2924 20256
rect 2872 20213 2881 20247
rect 2881 20213 2915 20247
rect 2915 20213 2924 20247
rect 2872 20204 2924 20213
rect 3976 20204 4028 20256
rect 9496 20340 9548 20392
rect 12164 20340 12216 20392
rect 18972 20383 19024 20392
rect 18972 20349 18981 20383
rect 18981 20349 19015 20383
rect 19015 20349 19024 20383
rect 18972 20340 19024 20349
rect 15200 20272 15252 20324
rect 18696 20272 18748 20324
rect 16120 20247 16172 20256
rect 16120 20213 16129 20247
rect 16129 20213 16163 20247
rect 16163 20213 16172 20247
rect 16120 20204 16172 20213
rect 3664 20102 3716 20154
rect 3728 20102 3780 20154
rect 3792 20102 3844 20154
rect 3856 20102 3908 20154
rect 3920 20102 3972 20154
rect 9092 20102 9144 20154
rect 9156 20102 9208 20154
rect 9220 20102 9272 20154
rect 9284 20102 9336 20154
rect 9348 20102 9400 20154
rect 14520 20102 14572 20154
rect 14584 20102 14636 20154
rect 14648 20102 14700 20154
rect 14712 20102 14764 20154
rect 14776 20102 14828 20154
rect 19948 20102 20000 20154
rect 20012 20102 20064 20154
rect 20076 20102 20128 20154
rect 20140 20102 20192 20154
rect 20204 20102 20256 20154
rect 3056 20043 3108 20052
rect 3056 20009 3065 20043
rect 3065 20009 3099 20043
rect 3099 20009 3108 20043
rect 3056 20000 3108 20009
rect 16028 20043 16080 20052
rect 16028 20009 16037 20043
rect 16037 20009 16071 20043
rect 16071 20009 16080 20043
rect 16028 20000 16080 20009
rect 1768 19932 1820 19984
rect 17040 19932 17092 19984
rect 1860 19864 1912 19916
rect 2228 19839 2280 19848
rect 2228 19805 2237 19839
rect 2237 19805 2271 19839
rect 2271 19805 2280 19839
rect 2228 19796 2280 19805
rect 2872 19796 2924 19848
rect 6000 19796 6052 19848
rect 11704 19796 11756 19848
rect 12164 19839 12216 19848
rect 12164 19805 12173 19839
rect 12173 19805 12207 19839
rect 12207 19805 12216 19839
rect 12164 19796 12216 19805
rect 13360 19796 13412 19848
rect 2504 19728 2556 19780
rect 2964 19728 3016 19780
rect 4528 19728 4580 19780
rect 14280 19728 14332 19780
rect 14372 19771 14424 19780
rect 14372 19737 14381 19771
rect 14381 19737 14415 19771
rect 14415 19737 14424 19771
rect 14372 19728 14424 19737
rect 15200 19771 15252 19780
rect 15200 19737 15209 19771
rect 15209 19737 15243 19771
rect 15243 19737 15252 19771
rect 15200 19728 15252 19737
rect 16396 19864 16448 19916
rect 17224 19796 17276 19848
rect 2412 19703 2464 19712
rect 2412 19669 2421 19703
rect 2421 19669 2455 19703
rect 2455 19669 2464 19703
rect 2412 19660 2464 19669
rect 4068 19660 4120 19712
rect 8300 19660 8352 19712
rect 15108 19660 15160 19712
rect 16396 19771 16448 19780
rect 16396 19737 16405 19771
rect 16405 19737 16439 19771
rect 16439 19737 16448 19771
rect 16396 19728 16448 19737
rect 6378 19558 6430 19610
rect 6442 19558 6494 19610
rect 6506 19558 6558 19610
rect 6570 19558 6622 19610
rect 6634 19558 6686 19610
rect 11806 19558 11858 19610
rect 11870 19558 11922 19610
rect 11934 19558 11986 19610
rect 11998 19558 12050 19610
rect 12062 19558 12114 19610
rect 17234 19558 17286 19610
rect 17298 19558 17350 19610
rect 17362 19558 17414 19610
rect 17426 19558 17478 19610
rect 17490 19558 17542 19610
rect 22662 19558 22714 19610
rect 22726 19558 22778 19610
rect 22790 19558 22842 19610
rect 22854 19558 22906 19610
rect 22918 19558 22970 19610
rect 2412 19388 2464 19440
rect 1860 19320 1912 19372
rect 2688 19320 2740 19372
rect 6000 19363 6052 19372
rect 6000 19329 6009 19363
rect 6009 19329 6043 19363
rect 6043 19329 6052 19363
rect 6000 19320 6052 19329
rect 7012 19320 7064 19372
rect 16120 19456 16172 19508
rect 13360 19388 13412 19440
rect 13544 19388 13596 19440
rect 9772 19363 9824 19372
rect 9772 19329 9806 19363
rect 9806 19329 9824 19363
rect 9772 19320 9824 19329
rect 17040 19388 17092 19440
rect 9496 19295 9548 19304
rect 9496 19261 9505 19295
rect 9505 19261 9539 19295
rect 9539 19261 9548 19295
rect 9496 19252 9548 19261
rect 11704 19252 11756 19304
rect 16580 19320 16632 19372
rect 18696 19388 18748 19440
rect 18604 19320 18656 19372
rect 18972 19320 19024 19372
rect 15476 19252 15528 19304
rect 16028 19252 16080 19304
rect 16488 19252 16540 19304
rect 17132 19295 17184 19304
rect 17132 19261 17141 19295
rect 17141 19261 17175 19295
rect 17175 19261 17184 19295
rect 17132 19252 17184 19261
rect 14280 19184 14332 19236
rect 4620 19159 4672 19168
rect 4620 19125 4629 19159
rect 4629 19125 4663 19159
rect 4663 19125 4672 19159
rect 4620 19116 4672 19125
rect 8392 19116 8444 19168
rect 16396 19116 16448 19168
rect 19340 19252 19392 19304
rect 18696 19159 18748 19168
rect 18696 19125 18705 19159
rect 18705 19125 18739 19159
rect 18739 19125 18748 19159
rect 18696 19116 18748 19125
rect 19616 19159 19668 19168
rect 19616 19125 19625 19159
rect 19625 19125 19659 19159
rect 19659 19125 19668 19159
rect 19616 19116 19668 19125
rect 3664 19014 3716 19066
rect 3728 19014 3780 19066
rect 3792 19014 3844 19066
rect 3856 19014 3908 19066
rect 3920 19014 3972 19066
rect 9092 19014 9144 19066
rect 9156 19014 9208 19066
rect 9220 19014 9272 19066
rect 9284 19014 9336 19066
rect 9348 19014 9400 19066
rect 14520 19014 14572 19066
rect 14584 19014 14636 19066
rect 14648 19014 14700 19066
rect 14712 19014 14764 19066
rect 14776 19014 14828 19066
rect 19948 19014 20000 19066
rect 20012 19014 20064 19066
rect 20076 19014 20128 19066
rect 20140 19014 20192 19066
rect 20204 19014 20256 19066
rect 4528 18955 4580 18964
rect 4528 18921 4537 18955
rect 4537 18921 4571 18955
rect 4571 18921 4580 18955
rect 4528 18912 4580 18921
rect 9680 18912 9732 18964
rect 15108 18912 15160 18964
rect 16580 18955 16632 18964
rect 16580 18921 16589 18955
rect 16589 18921 16623 18955
rect 16623 18921 16632 18955
rect 16580 18912 16632 18921
rect 6000 18776 6052 18828
rect 2688 18708 2740 18760
rect 4620 18708 4672 18760
rect 8116 18751 8168 18760
rect 8116 18717 8125 18751
rect 8125 18717 8159 18751
rect 8159 18717 8168 18751
rect 8116 18708 8168 18717
rect 8392 18708 8444 18760
rect 13544 18776 13596 18828
rect 4068 18640 4120 18692
rect 11704 18708 11756 18760
rect 15292 18708 15344 18760
rect 15660 18708 15712 18760
rect 16488 18708 16540 18760
rect 18604 18708 18656 18760
rect 18696 18751 18748 18760
rect 18696 18717 18705 18751
rect 18705 18717 18739 18751
rect 18739 18717 18748 18751
rect 18696 18708 18748 18717
rect 20444 18776 20496 18828
rect 17040 18640 17092 18692
rect 19616 18751 19668 18760
rect 19616 18717 19625 18751
rect 19625 18717 19659 18751
rect 19659 18717 19668 18751
rect 19616 18708 19668 18717
rect 20996 18640 21048 18692
rect 3424 18615 3476 18624
rect 3424 18581 3433 18615
rect 3433 18581 3467 18615
rect 3467 18581 3476 18615
rect 3424 18572 3476 18581
rect 9588 18572 9640 18624
rect 15752 18572 15804 18624
rect 17132 18572 17184 18624
rect 18512 18615 18564 18624
rect 18512 18581 18521 18615
rect 18521 18581 18555 18615
rect 18555 18581 18564 18615
rect 18512 18572 18564 18581
rect 19616 18615 19668 18624
rect 19616 18581 19625 18615
rect 19625 18581 19659 18615
rect 19659 18581 19668 18615
rect 19616 18572 19668 18581
rect 6378 18470 6430 18522
rect 6442 18470 6494 18522
rect 6506 18470 6558 18522
rect 6570 18470 6622 18522
rect 6634 18470 6686 18522
rect 11806 18470 11858 18522
rect 11870 18470 11922 18522
rect 11934 18470 11986 18522
rect 11998 18470 12050 18522
rect 12062 18470 12114 18522
rect 17234 18470 17286 18522
rect 17298 18470 17350 18522
rect 17362 18470 17414 18522
rect 17426 18470 17478 18522
rect 17490 18470 17542 18522
rect 22662 18470 22714 18522
rect 22726 18470 22778 18522
rect 22790 18470 22842 18522
rect 22854 18470 22906 18522
rect 22918 18470 22970 18522
rect 4068 18411 4120 18420
rect 4068 18377 4077 18411
rect 4077 18377 4111 18411
rect 4111 18377 4120 18411
rect 4068 18368 4120 18377
rect 15292 18411 15344 18420
rect 15292 18377 15301 18411
rect 15301 18377 15335 18411
rect 15335 18377 15344 18411
rect 15292 18368 15344 18377
rect 2688 18300 2740 18352
rect 3424 18300 3476 18352
rect 1860 18207 1912 18216
rect 1860 18173 1869 18207
rect 1869 18173 1903 18207
rect 1903 18173 1912 18207
rect 1860 18164 1912 18173
rect 2596 18096 2648 18148
rect 4620 18232 4672 18284
rect 18512 18343 18564 18352
rect 18512 18309 18521 18343
rect 18521 18309 18555 18343
rect 18555 18309 18564 18343
rect 18512 18300 18564 18309
rect 19432 18343 19484 18352
rect 19432 18309 19441 18343
rect 19441 18309 19475 18343
rect 19475 18309 19484 18343
rect 19432 18300 19484 18309
rect 6000 18232 6052 18284
rect 8116 18232 8168 18284
rect 15476 18275 15528 18284
rect 15476 18241 15485 18275
rect 15485 18241 15519 18275
rect 15519 18241 15528 18275
rect 15476 18232 15528 18241
rect 15752 18275 15804 18284
rect 15752 18241 15761 18275
rect 15761 18241 15795 18275
rect 15795 18241 15804 18275
rect 15752 18232 15804 18241
rect 20444 18232 20496 18284
rect 12256 18164 12308 18216
rect 16028 18164 16080 18216
rect 18788 18207 18840 18216
rect 18788 18173 18797 18207
rect 18797 18173 18831 18207
rect 18831 18173 18840 18207
rect 18788 18164 18840 18173
rect 16212 18096 16264 18148
rect 3240 18028 3292 18080
rect 15660 18071 15712 18080
rect 15660 18037 15669 18071
rect 15669 18037 15703 18071
rect 15703 18037 15712 18071
rect 15660 18028 15712 18037
rect 18236 18071 18288 18080
rect 18236 18037 18245 18071
rect 18245 18037 18279 18071
rect 18279 18037 18288 18071
rect 18236 18028 18288 18037
rect 3664 17926 3716 17978
rect 3728 17926 3780 17978
rect 3792 17926 3844 17978
rect 3856 17926 3908 17978
rect 3920 17926 3972 17978
rect 9092 17926 9144 17978
rect 9156 17926 9208 17978
rect 9220 17926 9272 17978
rect 9284 17926 9336 17978
rect 9348 17926 9400 17978
rect 14520 17926 14572 17978
rect 14584 17926 14636 17978
rect 14648 17926 14700 17978
rect 14712 17926 14764 17978
rect 14776 17926 14828 17978
rect 19948 17926 20000 17978
rect 20012 17926 20064 17978
rect 20076 17926 20128 17978
rect 20140 17926 20192 17978
rect 20204 17926 20256 17978
rect 1860 17620 1912 17672
rect 2320 17620 2372 17672
rect 4620 17824 4672 17876
rect 6000 17824 6052 17876
rect 9680 17824 9732 17876
rect 11704 17867 11756 17876
rect 11704 17833 11713 17867
rect 11713 17833 11747 17867
rect 11747 17833 11756 17867
rect 11704 17824 11756 17833
rect 15476 17867 15528 17876
rect 15476 17833 15485 17867
rect 15485 17833 15519 17867
rect 15519 17833 15528 17867
rect 15476 17824 15528 17833
rect 3056 17663 3108 17672
rect 3056 17629 3065 17663
rect 3065 17629 3099 17663
rect 3099 17629 3108 17663
rect 3056 17620 3108 17629
rect 2504 17552 2556 17604
rect 10600 17552 10652 17604
rect 15200 17620 15252 17672
rect 15660 17620 15712 17672
rect 16212 17663 16264 17672
rect 16212 17629 16221 17663
rect 16221 17629 16255 17663
rect 16255 17629 16264 17663
rect 16212 17620 16264 17629
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 16396 17552 16448 17604
rect 18788 17552 18840 17604
rect 19248 17552 19300 17604
rect 19800 17595 19852 17604
rect 19800 17561 19809 17595
rect 19809 17561 19843 17595
rect 19843 17561 19852 17595
rect 19800 17552 19852 17561
rect 1952 17484 2004 17536
rect 2596 17484 2648 17536
rect 2872 17484 2924 17536
rect 12900 17484 12952 17536
rect 15752 17484 15804 17536
rect 16948 17484 17000 17536
rect 6378 17382 6430 17434
rect 6442 17382 6494 17434
rect 6506 17382 6558 17434
rect 6570 17382 6622 17434
rect 6634 17382 6686 17434
rect 11806 17382 11858 17434
rect 11870 17382 11922 17434
rect 11934 17382 11986 17434
rect 11998 17382 12050 17434
rect 12062 17382 12114 17434
rect 17234 17382 17286 17434
rect 17298 17382 17350 17434
rect 17362 17382 17414 17434
rect 17426 17382 17478 17434
rect 17490 17382 17542 17434
rect 22662 17382 22714 17434
rect 22726 17382 22778 17434
rect 22790 17382 22842 17434
rect 22854 17382 22906 17434
rect 22918 17382 22970 17434
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 2872 17280 2924 17332
rect 2320 17187 2372 17196
rect 2320 17153 2329 17187
rect 2329 17153 2363 17187
rect 2363 17153 2372 17187
rect 2320 17144 2372 17153
rect 3056 17187 3108 17196
rect 3056 17153 3065 17187
rect 3065 17153 3099 17187
rect 3099 17153 3108 17187
rect 3056 17144 3108 17153
rect 3240 17187 3292 17196
rect 3240 17153 3249 17187
rect 3249 17153 3283 17187
rect 3283 17153 3292 17187
rect 15200 17212 15252 17264
rect 19248 17280 19300 17332
rect 19340 17255 19392 17264
rect 19340 17221 19349 17255
rect 19349 17221 19383 17255
rect 19383 17221 19392 17255
rect 19340 17212 19392 17221
rect 19800 17212 19852 17264
rect 3240 17144 3292 17153
rect 2504 17076 2556 17128
rect 6000 17187 6052 17196
rect 6000 17153 6009 17187
rect 6009 17153 6043 17187
rect 6043 17153 6052 17187
rect 6000 17144 6052 17153
rect 7012 17144 7064 17196
rect 7472 17144 7524 17196
rect 11704 17144 11756 17196
rect 12900 17187 12952 17196
rect 12900 17153 12909 17187
rect 12909 17153 12943 17187
rect 12943 17153 12952 17187
rect 12900 17144 12952 17153
rect 16488 17144 16540 17196
rect 18236 17144 18288 17196
rect 18696 17144 18748 17196
rect 19524 17144 19576 17196
rect 19616 17144 19668 17196
rect 9680 17119 9732 17128
rect 9680 17085 9689 17119
rect 9689 17085 9723 17119
rect 9723 17085 9732 17119
rect 9680 17076 9732 17085
rect 14924 17008 14976 17060
rect 17684 17119 17736 17128
rect 17684 17085 17693 17119
rect 17693 17085 17727 17119
rect 17727 17085 17736 17119
rect 17684 17076 17736 17085
rect 20996 17187 21048 17196
rect 20996 17153 21005 17187
rect 21005 17153 21039 17187
rect 21039 17153 21048 17187
rect 20996 17144 21048 17153
rect 18236 17008 18288 17060
rect 3148 16983 3200 16992
rect 3148 16949 3157 16983
rect 3157 16949 3191 16983
rect 3191 16949 3200 16983
rect 3148 16940 3200 16949
rect 4988 16940 5040 16992
rect 8760 16983 8812 16992
rect 8760 16949 8769 16983
rect 8769 16949 8803 16983
rect 8803 16949 8812 16983
rect 8760 16940 8812 16949
rect 19708 16940 19760 16992
rect 20904 16983 20956 16992
rect 20904 16949 20913 16983
rect 20913 16949 20947 16983
rect 20947 16949 20956 16983
rect 20904 16940 20956 16949
rect 3664 16838 3716 16890
rect 3728 16838 3780 16890
rect 3792 16838 3844 16890
rect 3856 16838 3908 16890
rect 3920 16838 3972 16890
rect 9092 16838 9144 16890
rect 9156 16838 9208 16890
rect 9220 16838 9272 16890
rect 9284 16838 9336 16890
rect 9348 16838 9400 16890
rect 14520 16838 14572 16890
rect 14584 16838 14636 16890
rect 14648 16838 14700 16890
rect 14712 16838 14764 16890
rect 14776 16838 14828 16890
rect 19948 16838 20000 16890
rect 20012 16838 20064 16890
rect 20076 16838 20128 16890
rect 20140 16838 20192 16890
rect 20204 16838 20256 16890
rect 1952 16600 2004 16652
rect 6000 16736 6052 16788
rect 16488 16779 16540 16788
rect 16488 16745 16497 16779
rect 16497 16745 16531 16779
rect 16531 16745 16540 16779
rect 16488 16736 16540 16745
rect 18696 16779 18748 16788
rect 18696 16745 18705 16779
rect 18705 16745 18739 16779
rect 18739 16745 18748 16779
rect 18696 16736 18748 16745
rect 1768 16464 1820 16516
rect 3148 16532 3200 16584
rect 3240 16575 3292 16584
rect 3240 16541 3249 16575
rect 3249 16541 3283 16575
rect 3283 16541 3292 16575
rect 3240 16532 3292 16541
rect 3884 16532 3936 16584
rect 7012 16643 7064 16652
rect 7012 16609 7021 16643
rect 7021 16609 7055 16643
rect 7055 16609 7064 16643
rect 7012 16600 7064 16609
rect 9680 16600 9732 16652
rect 11704 16600 11756 16652
rect 16120 16643 16172 16652
rect 16120 16609 16129 16643
rect 16129 16609 16163 16643
rect 16163 16609 16172 16643
rect 16120 16600 16172 16609
rect 17684 16643 17736 16652
rect 17684 16609 17693 16643
rect 17693 16609 17727 16643
rect 17727 16609 17736 16643
rect 17684 16600 17736 16609
rect 16028 16575 16080 16584
rect 16028 16541 16037 16575
rect 16037 16541 16071 16575
rect 16071 16541 16080 16575
rect 16028 16532 16080 16541
rect 2412 16439 2464 16448
rect 2412 16405 2421 16439
rect 2421 16405 2455 16439
rect 2455 16405 2464 16439
rect 2412 16396 2464 16405
rect 3884 16396 3936 16448
rect 5816 16396 5868 16448
rect 8392 16439 8444 16448
rect 8392 16405 8401 16439
rect 8401 16405 8435 16439
rect 8435 16405 8444 16439
rect 8392 16396 8444 16405
rect 12164 16464 12216 16516
rect 14924 16464 14976 16516
rect 17224 16532 17276 16584
rect 19248 16600 19300 16652
rect 19616 16600 19668 16652
rect 18236 16575 18288 16584
rect 18236 16541 18245 16575
rect 18245 16541 18279 16575
rect 18279 16541 18288 16575
rect 18236 16532 18288 16541
rect 18328 16575 18380 16584
rect 18328 16541 18337 16575
rect 18337 16541 18371 16575
rect 18371 16541 18380 16575
rect 18328 16532 18380 16541
rect 18512 16575 18564 16584
rect 18512 16541 18521 16575
rect 18521 16541 18555 16575
rect 18555 16541 18564 16575
rect 18512 16532 18564 16541
rect 19432 16575 19484 16584
rect 19432 16541 19441 16575
rect 19441 16541 19475 16575
rect 19475 16541 19484 16575
rect 19432 16532 19484 16541
rect 19708 16575 19760 16584
rect 19708 16541 19717 16575
rect 19717 16541 19751 16575
rect 19751 16541 19760 16575
rect 19708 16532 19760 16541
rect 19616 16464 19668 16516
rect 15016 16396 15068 16448
rect 6378 16294 6430 16346
rect 6442 16294 6494 16346
rect 6506 16294 6558 16346
rect 6570 16294 6622 16346
rect 6634 16294 6686 16346
rect 11806 16294 11858 16346
rect 11870 16294 11922 16346
rect 11934 16294 11986 16346
rect 11998 16294 12050 16346
rect 12062 16294 12114 16346
rect 17234 16294 17286 16346
rect 17298 16294 17350 16346
rect 17362 16294 17414 16346
rect 17426 16294 17478 16346
rect 17490 16294 17542 16346
rect 22662 16294 22714 16346
rect 22726 16294 22778 16346
rect 22790 16294 22842 16346
rect 22854 16294 22906 16346
rect 22918 16294 22970 16346
rect 1768 16235 1820 16244
rect 1768 16201 1777 16235
rect 1777 16201 1811 16235
rect 1811 16201 1820 16235
rect 1768 16192 1820 16201
rect 2412 16192 2464 16244
rect 2964 16192 3016 16244
rect 2320 16124 2372 16176
rect 2596 16124 2648 16176
rect 3240 16192 3292 16244
rect 4068 16192 4120 16244
rect 2504 16056 2556 16108
rect 3148 16124 3200 16176
rect 2872 16099 2924 16108
rect 2872 16065 2881 16099
rect 2881 16065 2915 16099
rect 2915 16065 2924 16099
rect 2872 16056 2924 16065
rect 8300 16124 8352 16176
rect 2136 15988 2188 16040
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 17132 16099 17184 16108
rect 17132 16065 17141 16099
rect 17141 16065 17175 16099
rect 17175 16065 17184 16099
rect 17132 16056 17184 16065
rect 18512 16124 18564 16176
rect 19340 16056 19392 16108
rect 19524 16099 19576 16108
rect 19524 16065 19533 16099
rect 19533 16065 19567 16099
rect 19567 16065 19576 16099
rect 19524 16056 19576 16065
rect 20904 16056 20956 16108
rect 12348 15988 12400 16040
rect 16764 15988 16816 16040
rect 18604 15988 18656 16040
rect 2688 15963 2740 15972
rect 2688 15929 2697 15963
rect 2697 15929 2731 15963
rect 2731 15929 2740 15963
rect 2688 15920 2740 15929
rect 2964 15920 3016 15972
rect 7472 15920 7524 15972
rect 16120 15920 16172 15972
rect 18328 15920 18380 15972
rect 9680 15852 9732 15904
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 10600 15852 10652 15861
rect 16856 15852 16908 15904
rect 3664 15750 3716 15802
rect 3728 15750 3780 15802
rect 3792 15750 3844 15802
rect 3856 15750 3908 15802
rect 3920 15750 3972 15802
rect 9092 15750 9144 15802
rect 9156 15750 9208 15802
rect 9220 15750 9272 15802
rect 9284 15750 9336 15802
rect 9348 15750 9400 15802
rect 14520 15750 14572 15802
rect 14584 15750 14636 15802
rect 14648 15750 14700 15802
rect 14712 15750 14764 15802
rect 14776 15750 14828 15802
rect 19948 15750 20000 15802
rect 20012 15750 20064 15802
rect 20076 15750 20128 15802
rect 20140 15750 20192 15802
rect 20204 15750 20256 15802
rect 2136 15691 2188 15700
rect 2136 15657 2145 15691
rect 2145 15657 2179 15691
rect 2179 15657 2188 15691
rect 2136 15648 2188 15657
rect 16764 15648 16816 15700
rect 17132 15648 17184 15700
rect 2504 15580 2556 15632
rect 20076 15580 20128 15632
rect 2320 15555 2372 15564
rect 2320 15521 2329 15555
rect 2329 15521 2363 15555
rect 2363 15521 2372 15555
rect 2320 15512 2372 15521
rect 2596 15555 2648 15564
rect 2596 15521 2605 15555
rect 2605 15521 2639 15555
rect 2639 15521 2648 15555
rect 2596 15512 2648 15521
rect 3056 15512 3108 15564
rect 4068 15512 4120 15564
rect 1952 15444 2004 15496
rect 2688 15444 2740 15496
rect 9588 15487 9640 15496
rect 9588 15453 9597 15487
rect 9597 15453 9631 15487
rect 9631 15453 9640 15487
rect 9588 15444 9640 15453
rect 9680 15444 9732 15496
rect 12348 15487 12400 15496
rect 12348 15453 12357 15487
rect 12357 15453 12391 15487
rect 12391 15453 12400 15487
rect 12348 15444 12400 15453
rect 15384 15444 15436 15496
rect 16028 15444 16080 15496
rect 15108 15376 15160 15428
rect 16488 15419 16540 15428
rect 16488 15385 16497 15419
rect 16497 15385 16531 15419
rect 16531 15385 16540 15419
rect 16488 15376 16540 15385
rect 18328 15444 18380 15496
rect 19340 15444 19392 15496
rect 19708 15419 19760 15428
rect 19708 15385 19717 15419
rect 19717 15385 19751 15419
rect 19751 15385 19760 15419
rect 19708 15376 19760 15385
rect 10876 15308 10928 15360
rect 15568 15308 15620 15360
rect 17592 15308 17644 15360
rect 18788 15308 18840 15360
rect 6378 15206 6430 15258
rect 6442 15206 6494 15258
rect 6506 15206 6558 15258
rect 6570 15206 6622 15258
rect 6634 15206 6686 15258
rect 11806 15206 11858 15258
rect 11870 15206 11922 15258
rect 11934 15206 11986 15258
rect 11998 15206 12050 15258
rect 12062 15206 12114 15258
rect 17234 15206 17286 15258
rect 17298 15206 17350 15258
rect 17362 15206 17414 15258
rect 17426 15206 17478 15258
rect 17490 15206 17542 15258
rect 22662 15206 22714 15258
rect 22726 15206 22778 15258
rect 22790 15206 22842 15258
rect 22854 15206 22906 15258
rect 22918 15206 22970 15258
rect 2504 15104 2556 15156
rect 2596 15036 2648 15088
rect 2412 14968 2464 15020
rect 2872 15104 2924 15156
rect 8116 15104 8168 15156
rect 15108 15104 15160 15156
rect 17132 15104 17184 15156
rect 18880 15104 18932 15156
rect 19524 15104 19576 15156
rect 12164 15036 12216 15088
rect 3516 15011 3568 15020
rect 3516 14977 3525 15011
rect 3525 14977 3559 15011
rect 3559 14977 3568 15011
rect 3516 14968 3568 14977
rect 4068 14968 4120 15020
rect 13728 14968 13780 15020
rect 7656 14943 7708 14952
rect 7656 14909 7665 14943
rect 7665 14909 7699 14943
rect 7699 14909 7708 14943
rect 7656 14900 7708 14909
rect 12348 14943 12400 14952
rect 12348 14909 12357 14943
rect 12357 14909 12391 14943
rect 12391 14909 12400 14943
rect 12348 14900 12400 14909
rect 13636 14900 13688 14952
rect 15568 15011 15620 15020
rect 15568 14977 15577 15011
rect 15577 14977 15611 15011
rect 15611 14977 15620 15011
rect 15568 14968 15620 14977
rect 16120 14968 16172 15020
rect 16764 14968 16816 15020
rect 17960 14968 18012 15020
rect 18052 14968 18104 15020
rect 18512 15011 18564 15020
rect 18512 14977 18521 15011
rect 18521 14977 18555 15011
rect 18555 14977 18564 15011
rect 18512 14968 18564 14977
rect 19340 15011 19392 15020
rect 19340 14977 19349 15011
rect 19349 14977 19383 15011
rect 19383 14977 19392 15011
rect 19340 14968 19392 14977
rect 20076 15011 20128 15020
rect 20076 14977 20085 15011
rect 20085 14977 20119 15011
rect 20119 14977 20128 15011
rect 20076 14968 20128 14977
rect 15384 14832 15436 14884
rect 16488 14900 16540 14952
rect 5632 14764 5684 14816
rect 6000 14764 6052 14816
rect 8852 14764 8904 14816
rect 18788 14832 18840 14884
rect 19248 14943 19300 14952
rect 19248 14909 19257 14943
rect 19257 14909 19291 14943
rect 19291 14909 19300 14943
rect 19248 14900 19300 14909
rect 19524 14900 19576 14952
rect 19432 14832 19484 14884
rect 19800 14832 19852 14884
rect 16856 14807 16908 14816
rect 16856 14773 16865 14807
rect 16865 14773 16899 14807
rect 16899 14773 16908 14807
rect 16856 14764 16908 14773
rect 3664 14662 3716 14714
rect 3728 14662 3780 14714
rect 3792 14662 3844 14714
rect 3856 14662 3908 14714
rect 3920 14662 3972 14714
rect 9092 14662 9144 14714
rect 9156 14662 9208 14714
rect 9220 14662 9272 14714
rect 9284 14662 9336 14714
rect 9348 14662 9400 14714
rect 14520 14662 14572 14714
rect 14584 14662 14636 14714
rect 14648 14662 14700 14714
rect 14712 14662 14764 14714
rect 14776 14662 14828 14714
rect 19948 14662 20000 14714
rect 20012 14662 20064 14714
rect 20076 14662 20128 14714
rect 20140 14662 20192 14714
rect 20204 14662 20256 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 4068 14560 4120 14612
rect 12256 14560 12308 14612
rect 13360 14560 13412 14612
rect 16488 14560 16540 14612
rect 17040 14560 17092 14612
rect 18604 14560 18656 14612
rect 19616 14603 19668 14612
rect 19616 14569 19625 14603
rect 19625 14569 19659 14603
rect 19659 14569 19668 14603
rect 19616 14560 19668 14569
rect 19800 14603 19852 14612
rect 19800 14569 19809 14603
rect 19809 14569 19843 14603
rect 19843 14569 19852 14603
rect 19800 14560 19852 14569
rect 2136 14492 2188 14544
rect 2504 14356 2556 14408
rect 5632 14399 5684 14408
rect 5632 14365 5641 14399
rect 5641 14365 5675 14399
rect 5675 14365 5684 14399
rect 5632 14356 5684 14365
rect 8208 14356 8260 14408
rect 9588 14356 9640 14408
rect 11060 14356 11112 14408
rect 12348 14399 12400 14408
rect 12348 14365 12357 14399
rect 12357 14365 12391 14399
rect 12391 14365 12400 14399
rect 12348 14356 12400 14365
rect 17592 14492 17644 14544
rect 18788 14492 18840 14544
rect 20260 14492 20312 14544
rect 16672 14424 16724 14476
rect 16764 14399 16816 14408
rect 16764 14365 16773 14399
rect 16773 14365 16807 14399
rect 16807 14365 16816 14399
rect 16764 14356 16816 14365
rect 4620 14288 4672 14340
rect 7564 14288 7616 14340
rect 4160 14220 4212 14272
rect 5908 14220 5960 14272
rect 9772 14220 9824 14272
rect 10692 14220 10744 14272
rect 14648 14288 14700 14340
rect 15752 14288 15804 14340
rect 15660 14220 15712 14272
rect 16028 14263 16080 14272
rect 16028 14229 16037 14263
rect 16037 14229 16071 14263
rect 16071 14229 16080 14263
rect 16028 14220 16080 14229
rect 16856 14288 16908 14340
rect 17040 14399 17092 14408
rect 17040 14365 17049 14399
rect 17049 14365 17083 14399
rect 17083 14365 17092 14399
rect 17040 14356 17092 14365
rect 17960 14356 18012 14408
rect 18604 14399 18656 14408
rect 18604 14365 18613 14399
rect 18613 14365 18647 14399
rect 18647 14365 18656 14399
rect 18604 14356 18656 14365
rect 18788 14356 18840 14408
rect 19524 14356 19576 14408
rect 20444 14288 20496 14340
rect 17592 14263 17644 14272
rect 17592 14229 17601 14263
rect 17601 14229 17635 14263
rect 17635 14229 17644 14263
rect 17592 14220 17644 14229
rect 18696 14220 18748 14272
rect 19800 14220 19852 14272
rect 6378 14118 6430 14170
rect 6442 14118 6494 14170
rect 6506 14118 6558 14170
rect 6570 14118 6622 14170
rect 6634 14118 6686 14170
rect 11806 14118 11858 14170
rect 11870 14118 11922 14170
rect 11934 14118 11986 14170
rect 11998 14118 12050 14170
rect 12062 14118 12114 14170
rect 17234 14118 17286 14170
rect 17298 14118 17350 14170
rect 17362 14118 17414 14170
rect 17426 14118 17478 14170
rect 17490 14118 17542 14170
rect 22662 14118 22714 14170
rect 22726 14118 22778 14170
rect 22790 14118 22842 14170
rect 22854 14118 22906 14170
rect 22918 14118 22970 14170
rect 3516 14016 3568 14068
rect 11060 14016 11112 14068
rect 15568 14016 15620 14068
rect 20996 14016 21048 14068
rect 2044 13880 2096 13932
rect 5632 13948 5684 14000
rect 7656 13948 7708 14000
rect 8208 13948 8260 14000
rect 13912 13948 13964 14000
rect 15752 13948 15804 14000
rect 4528 13923 4580 13932
rect 4528 13889 4562 13923
rect 4562 13889 4580 13923
rect 4528 13880 4580 13889
rect 7288 13923 7340 13932
rect 7288 13889 7297 13923
rect 7297 13889 7331 13923
rect 7331 13889 7340 13923
rect 7288 13880 7340 13889
rect 6828 13812 6880 13864
rect 10048 13923 10100 13932
rect 10048 13889 10082 13923
rect 10082 13889 10100 13923
rect 10048 13880 10100 13889
rect 9772 13855 9824 13864
rect 9772 13821 9781 13855
rect 9781 13821 9815 13855
rect 9815 13821 9824 13855
rect 9772 13812 9824 13821
rect 12348 13812 12400 13864
rect 13636 13880 13688 13932
rect 14648 13923 14700 13932
rect 14648 13889 14657 13923
rect 14657 13889 14691 13923
rect 14691 13889 14700 13923
rect 14648 13880 14700 13889
rect 15200 13880 15252 13932
rect 15844 13923 15896 13932
rect 15844 13889 15853 13923
rect 15853 13889 15887 13923
rect 15887 13889 15896 13923
rect 15844 13880 15896 13889
rect 16028 13880 16080 13932
rect 16488 13880 16540 13932
rect 18696 13923 18748 13932
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 20352 13880 20404 13932
rect 5724 13676 5776 13728
rect 8668 13719 8720 13728
rect 8668 13685 8677 13719
rect 8677 13685 8711 13719
rect 8711 13685 8720 13719
rect 8668 13676 8720 13685
rect 11152 13719 11204 13728
rect 11152 13685 11161 13719
rect 11161 13685 11195 13719
rect 11195 13685 11204 13719
rect 11152 13676 11204 13685
rect 13912 13787 13964 13796
rect 13912 13753 13921 13787
rect 13921 13753 13955 13787
rect 13955 13753 13964 13787
rect 13912 13744 13964 13753
rect 15384 13855 15436 13864
rect 15384 13821 15393 13855
rect 15393 13821 15427 13855
rect 15427 13821 15436 13855
rect 15384 13812 15436 13821
rect 16212 13855 16264 13864
rect 16212 13821 16221 13855
rect 16221 13821 16255 13855
rect 16255 13821 16264 13855
rect 16212 13812 16264 13821
rect 16672 13812 16724 13864
rect 16948 13855 17000 13864
rect 16948 13821 16957 13855
rect 16957 13821 16991 13855
rect 16991 13821 17000 13855
rect 16948 13812 17000 13821
rect 18880 13855 18932 13864
rect 18880 13821 18889 13855
rect 18889 13821 18923 13855
rect 18923 13821 18932 13855
rect 18880 13812 18932 13821
rect 18972 13855 19024 13864
rect 18972 13821 18981 13855
rect 18981 13821 19015 13855
rect 19015 13821 19024 13855
rect 18972 13812 19024 13821
rect 19524 13812 19576 13864
rect 3664 13574 3716 13626
rect 3728 13574 3780 13626
rect 3792 13574 3844 13626
rect 3856 13574 3908 13626
rect 3920 13574 3972 13626
rect 9092 13574 9144 13626
rect 9156 13574 9208 13626
rect 9220 13574 9272 13626
rect 9284 13574 9336 13626
rect 9348 13574 9400 13626
rect 14520 13574 14572 13626
rect 14584 13574 14636 13626
rect 14648 13574 14700 13626
rect 14712 13574 14764 13626
rect 14776 13574 14828 13626
rect 19948 13574 20000 13626
rect 20012 13574 20064 13626
rect 20076 13574 20128 13626
rect 20140 13574 20192 13626
rect 20204 13574 20256 13626
rect 5632 13472 5684 13524
rect 7288 13472 7340 13524
rect 19708 13447 19760 13456
rect 19708 13413 19717 13447
rect 19717 13413 19751 13447
rect 19751 13413 19760 13447
rect 19708 13404 19760 13413
rect 10600 13268 10652 13320
rect 16764 13336 16816 13388
rect 19432 13336 19484 13388
rect 19892 13336 19944 13388
rect 16948 13268 17000 13320
rect 18052 13311 18104 13320
rect 18052 13277 18061 13311
rect 18061 13277 18095 13311
rect 18095 13277 18104 13311
rect 18052 13268 18104 13277
rect 18972 13268 19024 13320
rect 12348 13200 12400 13252
rect 16856 13200 16908 13252
rect 19248 13200 19300 13252
rect 16212 13175 16264 13184
rect 16212 13141 16221 13175
rect 16221 13141 16255 13175
rect 16255 13141 16264 13175
rect 16212 13132 16264 13141
rect 16580 13175 16632 13184
rect 16580 13141 16589 13175
rect 16589 13141 16623 13175
rect 16623 13141 16632 13175
rect 16580 13132 16632 13141
rect 18696 13175 18748 13184
rect 18696 13141 18705 13175
rect 18705 13141 18739 13175
rect 18739 13141 18748 13175
rect 18696 13132 18748 13141
rect 18972 13132 19024 13184
rect 6378 13030 6430 13082
rect 6442 13030 6494 13082
rect 6506 13030 6558 13082
rect 6570 13030 6622 13082
rect 6634 13030 6686 13082
rect 11806 13030 11858 13082
rect 11870 13030 11922 13082
rect 11934 13030 11986 13082
rect 11998 13030 12050 13082
rect 12062 13030 12114 13082
rect 17234 13030 17286 13082
rect 17298 13030 17350 13082
rect 17362 13030 17414 13082
rect 17426 13030 17478 13082
rect 17490 13030 17542 13082
rect 22662 13030 22714 13082
rect 22726 13030 22778 13082
rect 22790 13030 22842 13082
rect 22854 13030 22906 13082
rect 22918 13030 22970 13082
rect 8300 12860 8352 12912
rect 19892 12971 19944 12980
rect 19892 12937 19901 12971
rect 19901 12937 19935 12971
rect 19935 12937 19944 12971
rect 19892 12928 19944 12937
rect 19064 12860 19116 12912
rect 19524 12860 19576 12912
rect 4252 12792 4304 12844
rect 5632 12792 5684 12844
rect 11612 12792 11664 12844
rect 15200 12792 15252 12844
rect 16212 12792 16264 12844
rect 19616 12792 19668 12844
rect 4436 12588 4488 12640
rect 9772 12767 9824 12776
rect 9772 12733 9781 12767
rect 9781 12733 9815 12767
rect 9815 12733 9824 12767
rect 9772 12724 9824 12733
rect 12348 12724 12400 12776
rect 15384 12724 15436 12776
rect 18604 12724 18656 12776
rect 8208 12588 8260 12640
rect 9588 12588 9640 12640
rect 16856 12656 16908 12708
rect 18512 12656 18564 12708
rect 11060 12588 11112 12640
rect 13268 12588 13320 12640
rect 16580 12588 16632 12640
rect 18144 12588 18196 12640
rect 18696 12588 18748 12640
rect 18972 12631 19024 12640
rect 18972 12597 18981 12631
rect 18981 12597 19015 12631
rect 19015 12597 19024 12631
rect 18972 12588 19024 12597
rect 19340 12588 19392 12640
rect 19892 12588 19944 12640
rect 3664 12486 3716 12538
rect 3728 12486 3780 12538
rect 3792 12486 3844 12538
rect 3856 12486 3908 12538
rect 3920 12486 3972 12538
rect 9092 12486 9144 12538
rect 9156 12486 9208 12538
rect 9220 12486 9272 12538
rect 9284 12486 9336 12538
rect 9348 12486 9400 12538
rect 14520 12486 14572 12538
rect 14584 12486 14636 12538
rect 14648 12486 14700 12538
rect 14712 12486 14764 12538
rect 14776 12486 14828 12538
rect 19948 12486 20000 12538
rect 20012 12486 20064 12538
rect 20076 12486 20128 12538
rect 20140 12486 20192 12538
rect 20204 12486 20256 12538
rect 5724 12384 5776 12436
rect 6184 12384 6236 12436
rect 15292 12384 15344 12436
rect 15844 12316 15896 12368
rect 16948 12316 17000 12368
rect 1952 12180 2004 12232
rect 2228 12223 2280 12232
rect 2228 12189 2237 12223
rect 2237 12189 2271 12223
rect 2271 12189 2280 12223
rect 2228 12180 2280 12189
rect 3148 12248 3200 12300
rect 11060 12248 11112 12300
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 5632 12223 5684 12232
rect 5632 12189 5641 12223
rect 5641 12189 5675 12223
rect 5675 12189 5684 12223
rect 5632 12180 5684 12189
rect 8208 12180 8260 12232
rect 10324 12180 10376 12232
rect 15660 12248 15712 12300
rect 12348 12180 12400 12232
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 16580 12248 16632 12300
rect 17868 12248 17920 12300
rect 2780 12112 2832 12164
rect 6736 12112 6788 12164
rect 11244 12112 11296 12164
rect 13912 12112 13964 12164
rect 4160 12044 4212 12096
rect 7380 12044 7432 12096
rect 10508 12044 10560 12096
rect 13636 12044 13688 12096
rect 18328 12248 18380 12300
rect 19616 12291 19668 12300
rect 19616 12257 19625 12291
rect 19625 12257 19659 12291
rect 19659 12257 19668 12291
rect 19616 12248 19668 12257
rect 19892 12291 19944 12300
rect 19892 12257 19901 12291
rect 19901 12257 19935 12291
rect 19935 12257 19944 12291
rect 19892 12248 19944 12257
rect 18236 12112 18288 12164
rect 18604 12112 18656 12164
rect 19432 12112 19484 12164
rect 18512 12044 18564 12096
rect 19156 12044 19208 12096
rect 19340 12044 19392 12096
rect 19892 12044 19944 12096
rect 6378 11942 6430 11994
rect 6442 11942 6494 11994
rect 6506 11942 6558 11994
rect 6570 11942 6622 11994
rect 6634 11942 6686 11994
rect 11806 11942 11858 11994
rect 11870 11942 11922 11994
rect 11934 11942 11986 11994
rect 11998 11942 12050 11994
rect 12062 11942 12114 11994
rect 17234 11942 17286 11994
rect 17298 11942 17350 11994
rect 17362 11942 17414 11994
rect 17426 11942 17478 11994
rect 17490 11942 17542 11994
rect 22662 11942 22714 11994
rect 22726 11942 22778 11994
rect 22790 11942 22842 11994
rect 22854 11942 22906 11994
rect 22918 11942 22970 11994
rect 2596 11840 2648 11892
rect 2780 11840 2832 11892
rect 16856 11883 16908 11892
rect 16856 11849 16865 11883
rect 16865 11849 16899 11883
rect 16899 11849 16908 11883
rect 16856 11840 16908 11849
rect 18328 11840 18380 11892
rect 19340 11840 19392 11892
rect 19524 11883 19576 11892
rect 19524 11849 19533 11883
rect 19533 11849 19567 11883
rect 19567 11849 19576 11883
rect 19524 11840 19576 11849
rect 2688 11704 2740 11756
rect 4160 11772 4212 11824
rect 3148 11747 3200 11756
rect 3148 11713 3157 11747
rect 3157 11713 3191 11747
rect 3191 11713 3200 11747
rect 3148 11704 3200 11713
rect 5632 11772 5684 11824
rect 2596 11636 2648 11688
rect 4160 11636 4212 11688
rect 8208 11704 8260 11756
rect 8576 11747 8628 11756
rect 8576 11713 8610 11747
rect 8610 11713 8628 11747
rect 8576 11704 8628 11713
rect 12348 11704 12400 11756
rect 13176 11704 13228 11756
rect 15660 11747 15712 11756
rect 15660 11713 15669 11747
rect 15669 11713 15703 11747
rect 15703 11713 15712 11747
rect 15660 11704 15712 11713
rect 15200 11636 15252 11688
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 17592 11704 17644 11756
rect 18236 11704 18288 11756
rect 18972 11747 19024 11756
rect 18972 11713 18981 11747
rect 18981 11713 19015 11747
rect 19015 11713 19024 11747
rect 18972 11704 19024 11713
rect 19156 11747 19208 11756
rect 19156 11713 19165 11747
rect 19165 11713 19199 11747
rect 19199 11713 19208 11747
rect 19156 11704 19208 11713
rect 19616 11747 19668 11756
rect 19616 11713 19625 11747
rect 19625 11713 19659 11747
rect 19659 11713 19668 11747
rect 19616 11704 19668 11713
rect 15476 11568 15528 11620
rect 16488 11568 16540 11620
rect 6000 11500 6052 11552
rect 9680 11543 9732 11552
rect 9680 11509 9689 11543
rect 9689 11509 9723 11543
rect 9723 11509 9732 11543
rect 9680 11500 9732 11509
rect 15568 11500 15620 11552
rect 3664 11398 3716 11450
rect 3728 11398 3780 11450
rect 3792 11398 3844 11450
rect 3856 11398 3908 11450
rect 3920 11398 3972 11450
rect 9092 11398 9144 11450
rect 9156 11398 9208 11450
rect 9220 11398 9272 11450
rect 9284 11398 9336 11450
rect 9348 11398 9400 11450
rect 14520 11398 14572 11450
rect 14584 11398 14636 11450
rect 14648 11398 14700 11450
rect 14712 11398 14764 11450
rect 14776 11398 14828 11450
rect 19948 11398 20000 11450
rect 20012 11398 20064 11450
rect 20076 11398 20128 11450
rect 20140 11398 20192 11450
rect 20204 11398 20256 11450
rect 7472 11228 7524 11280
rect 15568 11228 15620 11280
rect 16304 11228 16356 11280
rect 5632 11160 5684 11212
rect 15660 11160 15712 11212
rect 18604 11160 18656 11212
rect 17868 11092 17920 11144
rect 18328 11135 18380 11144
rect 18328 11101 18337 11135
rect 18337 11101 18371 11135
rect 18371 11101 18380 11135
rect 18328 11092 18380 11101
rect 5908 11024 5960 11076
rect 17040 11024 17092 11076
rect 6378 10854 6430 10906
rect 6442 10854 6494 10906
rect 6506 10854 6558 10906
rect 6570 10854 6622 10906
rect 6634 10854 6686 10906
rect 11806 10854 11858 10906
rect 11870 10854 11922 10906
rect 11934 10854 11986 10906
rect 11998 10854 12050 10906
rect 12062 10854 12114 10906
rect 17234 10854 17286 10906
rect 17298 10854 17350 10906
rect 17362 10854 17414 10906
rect 17426 10854 17478 10906
rect 17490 10854 17542 10906
rect 22662 10854 22714 10906
rect 22726 10854 22778 10906
rect 22790 10854 22842 10906
rect 22854 10854 22906 10906
rect 22918 10854 22970 10906
rect 2044 10684 2096 10736
rect 2596 10752 2648 10804
rect 4344 10752 4396 10804
rect 5632 10752 5684 10804
rect 6644 10752 6696 10804
rect 8300 10752 8352 10804
rect 13912 10752 13964 10804
rect 4160 10684 4212 10736
rect 2320 10616 2372 10668
rect 3516 10659 3568 10668
rect 3516 10625 3525 10659
rect 3525 10625 3559 10659
rect 3559 10625 3568 10659
rect 3516 10616 3568 10625
rect 4436 10616 4488 10668
rect 2044 10523 2096 10532
rect 2044 10489 2053 10523
rect 2053 10489 2087 10523
rect 2087 10489 2096 10523
rect 2044 10480 2096 10489
rect 6184 10480 6236 10532
rect 5908 10455 5960 10464
rect 5908 10421 5917 10455
rect 5917 10421 5951 10455
rect 5951 10421 5960 10455
rect 5908 10412 5960 10421
rect 7748 10684 7800 10736
rect 6644 10616 6696 10668
rect 7656 10616 7708 10668
rect 9680 10684 9732 10736
rect 7288 10548 7340 10600
rect 7380 10591 7432 10600
rect 7380 10557 7389 10591
rect 7389 10557 7423 10591
rect 7423 10557 7432 10591
rect 7380 10548 7432 10557
rect 8484 10659 8536 10668
rect 8484 10625 8493 10659
rect 8493 10625 8527 10659
rect 8527 10625 8536 10659
rect 8484 10616 8536 10625
rect 9588 10616 9640 10668
rect 13084 10659 13136 10668
rect 13084 10625 13093 10659
rect 13093 10625 13127 10659
rect 13127 10625 13136 10659
rect 13084 10616 13136 10625
rect 13452 10616 13504 10668
rect 15292 10616 15344 10668
rect 15752 10616 15804 10668
rect 13360 10591 13412 10600
rect 13360 10557 13369 10591
rect 13369 10557 13403 10591
rect 13403 10557 13412 10591
rect 13360 10548 13412 10557
rect 8300 10480 8352 10532
rect 9496 10480 9548 10532
rect 14924 10480 14976 10532
rect 15660 10548 15712 10600
rect 16580 10616 16632 10668
rect 18236 10659 18288 10668
rect 18236 10625 18245 10659
rect 18245 10625 18279 10659
rect 18279 10625 18288 10659
rect 18236 10616 18288 10625
rect 18604 10659 18656 10668
rect 18604 10625 18613 10659
rect 18613 10625 18647 10659
rect 18647 10625 18656 10659
rect 18604 10616 18656 10625
rect 18696 10659 18748 10668
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 19340 10616 19392 10668
rect 20444 10616 20496 10668
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 16212 10480 16264 10532
rect 6644 10455 6696 10464
rect 6644 10421 6653 10455
rect 6653 10421 6687 10455
rect 6687 10421 6696 10455
rect 6644 10412 6696 10421
rect 8116 10412 8168 10464
rect 13820 10412 13872 10464
rect 15660 10455 15712 10464
rect 15660 10421 15669 10455
rect 15669 10421 15703 10455
rect 15703 10421 15712 10455
rect 15660 10412 15712 10421
rect 16948 10412 17000 10464
rect 18972 10455 19024 10464
rect 18972 10421 18981 10455
rect 18981 10421 19015 10455
rect 19015 10421 19024 10455
rect 18972 10412 19024 10421
rect 3664 10310 3716 10362
rect 3728 10310 3780 10362
rect 3792 10310 3844 10362
rect 3856 10310 3908 10362
rect 3920 10310 3972 10362
rect 9092 10310 9144 10362
rect 9156 10310 9208 10362
rect 9220 10310 9272 10362
rect 9284 10310 9336 10362
rect 9348 10310 9400 10362
rect 14520 10310 14572 10362
rect 14584 10310 14636 10362
rect 14648 10310 14700 10362
rect 14712 10310 14764 10362
rect 14776 10310 14828 10362
rect 19948 10310 20000 10362
rect 20012 10310 20064 10362
rect 20076 10310 20128 10362
rect 20140 10310 20192 10362
rect 20204 10310 20256 10362
rect 2320 10251 2372 10260
rect 2320 10217 2329 10251
rect 2329 10217 2363 10251
rect 2363 10217 2372 10251
rect 2320 10208 2372 10217
rect 2688 10208 2740 10260
rect 2412 10140 2464 10192
rect 2688 10072 2740 10124
rect 1860 9936 1912 9988
rect 3516 10140 3568 10192
rect 5632 10208 5684 10260
rect 6736 10208 6788 10260
rect 8484 10208 8536 10260
rect 10324 10251 10376 10260
rect 10324 10217 10333 10251
rect 10333 10217 10367 10251
rect 10367 10217 10376 10251
rect 10324 10208 10376 10217
rect 11244 10251 11296 10260
rect 11244 10217 11253 10251
rect 11253 10217 11287 10251
rect 11287 10217 11296 10251
rect 11244 10208 11296 10217
rect 12256 10251 12308 10260
rect 12256 10217 12265 10251
rect 12265 10217 12299 10251
rect 12299 10217 12308 10251
rect 12256 10208 12308 10217
rect 12348 10208 12400 10260
rect 13084 10208 13136 10260
rect 13820 10208 13872 10260
rect 18972 10208 19024 10260
rect 19800 10208 19852 10260
rect 4160 10072 4212 10124
rect 4344 10004 4396 10056
rect 5724 10047 5776 10056
rect 5724 10013 5733 10047
rect 5733 10013 5767 10047
rect 5767 10013 5776 10047
rect 5724 10004 5776 10013
rect 5908 10047 5960 10056
rect 5908 10013 5917 10047
rect 5917 10013 5951 10047
rect 5951 10013 5960 10047
rect 5908 10004 5960 10013
rect 6644 10072 6696 10124
rect 6184 10004 6236 10056
rect 7380 10072 7432 10124
rect 8300 10072 8352 10124
rect 15384 10140 15436 10192
rect 18420 10183 18472 10192
rect 18420 10149 18429 10183
rect 18429 10149 18463 10183
rect 18463 10149 18472 10183
rect 18420 10140 18472 10149
rect 19248 10140 19300 10192
rect 13360 10072 13412 10124
rect 14924 10115 14976 10124
rect 14924 10081 14933 10115
rect 14933 10081 14967 10115
rect 14967 10081 14976 10115
rect 14924 10072 14976 10081
rect 15660 10072 15712 10124
rect 16028 10072 16080 10124
rect 17040 10072 17092 10124
rect 18512 10115 18564 10124
rect 18512 10081 18521 10115
rect 18521 10081 18555 10115
rect 18555 10081 18564 10115
rect 18512 10072 18564 10081
rect 7656 10047 7708 10056
rect 7656 10013 7665 10047
rect 7665 10013 7699 10047
rect 7699 10013 7708 10047
rect 7656 10004 7708 10013
rect 9588 10047 9640 10056
rect 9588 10013 9597 10047
rect 9597 10013 9631 10047
rect 9631 10013 9640 10047
rect 9588 10004 9640 10013
rect 10600 10004 10652 10056
rect 11704 10004 11756 10056
rect 13452 10047 13504 10056
rect 13452 10013 13461 10047
rect 13461 10013 13495 10047
rect 13495 10013 13504 10047
rect 13452 10004 13504 10013
rect 4712 9979 4764 9988
rect 4712 9945 4721 9979
rect 4721 9945 4755 9979
rect 4755 9945 4764 9979
rect 4712 9936 4764 9945
rect 5632 9936 5684 9988
rect 10784 9979 10836 9988
rect 10784 9945 10793 9979
rect 10793 9945 10827 9979
rect 10827 9945 10836 9979
rect 10784 9936 10836 9945
rect 12348 9936 12400 9988
rect 12440 9979 12492 9988
rect 12440 9945 12449 9979
rect 12449 9945 12483 9979
rect 12483 9945 12492 9979
rect 12440 9936 12492 9945
rect 14832 10047 14884 10056
rect 14832 10013 14841 10047
rect 14841 10013 14875 10047
rect 14875 10013 14884 10047
rect 14832 10004 14884 10013
rect 15200 10004 15252 10056
rect 15476 10047 15528 10056
rect 15476 10013 15485 10047
rect 15485 10013 15519 10047
rect 15519 10013 15528 10047
rect 15476 10004 15528 10013
rect 15752 10047 15804 10056
rect 15752 10013 15761 10047
rect 15761 10013 15795 10047
rect 15795 10013 15804 10047
rect 15752 10004 15804 10013
rect 18052 10004 18104 10056
rect 19432 10047 19484 10056
rect 19432 10013 19441 10047
rect 19441 10013 19475 10047
rect 19475 10013 19484 10047
rect 19432 10004 19484 10013
rect 1768 9868 1820 9920
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 4436 9868 4488 9920
rect 6184 9868 6236 9920
rect 6368 9868 6420 9920
rect 7748 9911 7800 9920
rect 7748 9877 7757 9911
rect 7757 9877 7791 9911
rect 7791 9877 7800 9911
rect 7748 9868 7800 9877
rect 9496 9911 9548 9920
rect 9496 9877 9505 9911
rect 9505 9877 9539 9911
rect 9539 9877 9548 9911
rect 9496 9868 9548 9877
rect 10508 9868 10560 9920
rect 10968 9868 11020 9920
rect 15292 9936 15344 9988
rect 15844 9936 15896 9988
rect 16580 9936 16632 9988
rect 17960 9936 18012 9988
rect 15108 9868 15160 9920
rect 15936 9911 15988 9920
rect 15936 9877 15945 9911
rect 15945 9877 15979 9911
rect 15979 9877 15988 9911
rect 15936 9868 15988 9877
rect 20352 9868 20404 9920
rect 6378 9766 6430 9818
rect 6442 9766 6494 9818
rect 6506 9766 6558 9818
rect 6570 9766 6622 9818
rect 6634 9766 6686 9818
rect 11806 9766 11858 9818
rect 11870 9766 11922 9818
rect 11934 9766 11986 9818
rect 11998 9766 12050 9818
rect 12062 9766 12114 9818
rect 17234 9766 17286 9818
rect 17298 9766 17350 9818
rect 17362 9766 17414 9818
rect 17426 9766 17478 9818
rect 17490 9766 17542 9818
rect 22662 9766 22714 9818
rect 22726 9766 22778 9818
rect 22790 9766 22842 9818
rect 22854 9766 22906 9818
rect 22918 9766 22970 9818
rect 1860 9707 1912 9716
rect 1860 9673 1869 9707
rect 1869 9673 1903 9707
rect 1903 9673 1912 9707
rect 1860 9664 1912 9673
rect 2228 9664 2280 9716
rect 5724 9664 5776 9716
rect 6736 9707 6788 9716
rect 2412 9596 2464 9648
rect 5632 9639 5684 9648
rect 5632 9605 5641 9639
rect 5641 9605 5675 9639
rect 5675 9605 5684 9639
rect 5632 9596 5684 9605
rect 6736 9673 6763 9707
rect 6763 9673 6788 9707
rect 6736 9664 6788 9673
rect 8576 9664 8628 9716
rect 9496 9664 9548 9716
rect 10784 9664 10836 9716
rect 7288 9596 7340 9648
rect 7932 9639 7984 9648
rect 7932 9605 7941 9639
rect 7941 9605 7975 9639
rect 7975 9605 7984 9639
rect 7932 9596 7984 9605
rect 8300 9639 8352 9648
rect 8300 9605 8309 9639
rect 8309 9605 8343 9639
rect 8343 9605 8352 9639
rect 8300 9596 8352 9605
rect 12440 9664 12492 9716
rect 16120 9664 16172 9716
rect 15200 9596 15252 9648
rect 16028 9596 16080 9648
rect 1768 9571 1820 9580
rect 1768 9537 1777 9571
rect 1777 9537 1811 9571
rect 1811 9537 1820 9571
rect 1768 9528 1820 9537
rect 7748 9528 7800 9580
rect 8208 9528 8260 9580
rect 8116 9503 8168 9512
rect 8116 9469 8125 9503
rect 8125 9469 8159 9503
rect 8159 9469 8168 9503
rect 8116 9460 8168 9469
rect 2044 9435 2096 9444
rect 2044 9401 2053 9435
rect 2053 9401 2087 9435
rect 2087 9401 2096 9435
rect 2044 9392 2096 9401
rect 6276 9324 6328 9376
rect 7288 9392 7340 9444
rect 9588 9528 9640 9580
rect 10968 9528 11020 9580
rect 11428 9528 11480 9580
rect 12348 9528 12400 9580
rect 13268 9571 13320 9580
rect 13268 9537 13277 9571
rect 13277 9537 13311 9571
rect 13311 9537 13320 9571
rect 13268 9528 13320 9537
rect 14004 9528 14056 9580
rect 14832 9528 14884 9580
rect 15936 9571 15988 9580
rect 15936 9537 15945 9571
rect 15945 9537 15979 9571
rect 15979 9537 15988 9571
rect 15936 9528 15988 9537
rect 10600 9435 10652 9444
rect 10600 9401 10609 9435
rect 10609 9401 10643 9435
rect 10643 9401 10652 9435
rect 10600 9392 10652 9401
rect 11704 9435 11756 9444
rect 11704 9401 11713 9435
rect 11713 9401 11747 9435
rect 11747 9401 11756 9435
rect 11704 9392 11756 9401
rect 12256 9460 12308 9512
rect 15476 9460 15528 9512
rect 16304 9639 16356 9648
rect 16304 9605 16313 9639
rect 16313 9605 16347 9639
rect 16347 9605 16356 9639
rect 16304 9596 16356 9605
rect 18788 9664 18840 9716
rect 17960 9596 18012 9648
rect 12532 9392 12584 9444
rect 13360 9392 13412 9444
rect 13452 9324 13504 9376
rect 18696 9528 18748 9580
rect 18880 9528 18932 9580
rect 16396 9460 16448 9512
rect 3664 9222 3716 9274
rect 3728 9222 3780 9274
rect 3792 9222 3844 9274
rect 3856 9222 3908 9274
rect 3920 9222 3972 9274
rect 9092 9222 9144 9274
rect 9156 9222 9208 9274
rect 9220 9222 9272 9274
rect 9284 9222 9336 9274
rect 9348 9222 9400 9274
rect 14520 9222 14572 9274
rect 14584 9222 14636 9274
rect 14648 9222 14700 9274
rect 14712 9222 14764 9274
rect 14776 9222 14828 9274
rect 19948 9222 20000 9274
rect 20012 9222 20064 9274
rect 20076 9222 20128 9274
rect 20140 9222 20192 9274
rect 20204 9222 20256 9274
rect 2412 9120 2464 9172
rect 7748 9120 7800 9172
rect 13176 9163 13228 9172
rect 13176 9129 13185 9163
rect 13185 9129 13219 9163
rect 13219 9129 13228 9163
rect 13176 9120 13228 9129
rect 13360 9163 13412 9172
rect 13360 9129 13369 9163
rect 13369 9129 13403 9163
rect 13403 9129 13412 9163
rect 13360 9120 13412 9129
rect 15752 9163 15804 9172
rect 15752 9129 15761 9163
rect 15761 9129 15795 9163
rect 15795 9129 15804 9163
rect 15752 9120 15804 9129
rect 16120 9163 16172 9172
rect 16120 9129 16129 9163
rect 16129 9129 16163 9163
rect 16163 9129 16172 9163
rect 16120 9120 16172 9129
rect 19432 9120 19484 9172
rect 2596 8984 2648 9036
rect 4344 8984 4396 9036
rect 5448 8984 5500 9036
rect 7288 9027 7340 9036
rect 7288 8993 7297 9027
rect 7297 8993 7331 9027
rect 7331 8993 7340 9027
rect 7288 8984 7340 8993
rect 4252 8959 4304 8968
rect 4252 8925 4261 8959
rect 4261 8925 4295 8959
rect 4295 8925 4304 8959
rect 4252 8916 4304 8925
rect 7472 8959 7524 8968
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 13360 8984 13412 9036
rect 19340 8984 19392 9036
rect 12624 8959 12676 8968
rect 12624 8925 12633 8959
rect 12633 8925 12667 8959
rect 12667 8925 12676 8959
rect 12624 8916 12676 8925
rect 15292 8916 15344 8968
rect 16212 8916 16264 8968
rect 18328 8916 18380 8968
rect 18696 8959 18748 8968
rect 18696 8925 18705 8959
rect 18705 8925 18739 8959
rect 18739 8925 18748 8959
rect 18696 8916 18748 8925
rect 6000 8848 6052 8900
rect 12164 8848 12216 8900
rect 4160 8780 4212 8832
rect 12256 8780 12308 8832
rect 13452 8848 13504 8900
rect 16396 8848 16448 8900
rect 6378 8678 6430 8730
rect 6442 8678 6494 8730
rect 6506 8678 6558 8730
rect 6570 8678 6622 8730
rect 6634 8678 6686 8730
rect 11806 8678 11858 8730
rect 11870 8678 11922 8730
rect 11934 8678 11986 8730
rect 11998 8678 12050 8730
rect 12062 8678 12114 8730
rect 17234 8678 17286 8730
rect 17298 8678 17350 8730
rect 17362 8678 17414 8730
rect 17426 8678 17478 8730
rect 17490 8678 17542 8730
rect 22662 8678 22714 8730
rect 22726 8678 22778 8730
rect 22790 8678 22842 8730
rect 22854 8678 22906 8730
rect 22918 8678 22970 8730
rect 4620 8576 4672 8628
rect 6828 8619 6880 8628
rect 6828 8585 6830 8619
rect 6830 8585 6864 8619
rect 6864 8585 6880 8619
rect 6828 8576 6880 8585
rect 3148 8440 3200 8492
rect 3516 8440 3568 8492
rect 4344 8508 4396 8560
rect 3424 8304 3476 8356
rect 4160 8440 4212 8492
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 5908 8440 5960 8492
rect 7380 8508 7432 8560
rect 6736 8483 6788 8492
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 7288 8440 7340 8492
rect 11612 8576 11664 8628
rect 12164 8576 12216 8628
rect 13636 8576 13688 8628
rect 11152 8551 11204 8560
rect 11152 8517 11161 8551
rect 11161 8517 11195 8551
rect 11195 8517 11204 8551
rect 11152 8508 11204 8517
rect 12624 8508 12676 8560
rect 4712 8415 4764 8424
rect 4712 8381 4721 8415
rect 4721 8381 4755 8415
rect 4755 8381 4764 8415
rect 4712 8372 4764 8381
rect 6000 8372 6052 8424
rect 9588 8440 9640 8492
rect 11428 8440 11480 8492
rect 15200 8508 15252 8560
rect 8484 8372 8536 8424
rect 9404 8415 9456 8424
rect 9404 8381 9413 8415
rect 9413 8381 9447 8415
rect 9447 8381 9456 8415
rect 9404 8372 9456 8381
rect 9772 8415 9824 8424
rect 9772 8381 9781 8415
rect 9781 8381 9815 8415
rect 9815 8381 9824 8415
rect 9772 8372 9824 8381
rect 7472 8304 7524 8356
rect 9496 8304 9548 8356
rect 5080 8279 5132 8288
rect 5080 8245 5089 8279
rect 5089 8245 5123 8279
rect 5123 8245 5132 8279
rect 5080 8236 5132 8245
rect 8944 8236 8996 8288
rect 9404 8236 9456 8288
rect 9956 8279 10008 8288
rect 9956 8245 9965 8279
rect 9965 8245 9999 8279
rect 9999 8245 10008 8279
rect 9956 8236 10008 8245
rect 10692 8372 10744 8424
rect 14372 8440 14424 8492
rect 14924 8440 14976 8492
rect 17960 8576 18012 8628
rect 16488 8508 16540 8560
rect 18328 8508 18380 8560
rect 13360 8372 13412 8424
rect 15476 8372 15528 8424
rect 12256 8304 12308 8356
rect 10968 8236 11020 8288
rect 14004 8304 14056 8356
rect 13912 8279 13964 8288
rect 13912 8245 13921 8279
rect 13921 8245 13955 8279
rect 13955 8245 13964 8279
rect 13912 8236 13964 8245
rect 15016 8236 15068 8288
rect 16488 8372 16540 8424
rect 18236 8440 18288 8492
rect 19064 8440 19116 8492
rect 16580 8304 16632 8356
rect 18788 8304 18840 8356
rect 19340 8347 19392 8356
rect 19340 8313 19349 8347
rect 19349 8313 19383 8347
rect 19383 8313 19392 8347
rect 19340 8304 19392 8313
rect 3664 8134 3716 8186
rect 3728 8134 3780 8186
rect 3792 8134 3844 8186
rect 3856 8134 3908 8186
rect 3920 8134 3972 8186
rect 9092 8134 9144 8186
rect 9156 8134 9208 8186
rect 9220 8134 9272 8186
rect 9284 8134 9336 8186
rect 9348 8134 9400 8186
rect 14520 8134 14572 8186
rect 14584 8134 14636 8186
rect 14648 8134 14700 8186
rect 14712 8134 14764 8186
rect 14776 8134 14828 8186
rect 19948 8134 20000 8186
rect 20012 8134 20064 8186
rect 20076 8134 20128 8186
rect 20140 8134 20192 8186
rect 20204 8134 20256 8186
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 3516 8032 3568 8084
rect 4252 8032 4304 8084
rect 4896 8032 4948 8084
rect 4160 7828 4212 7880
rect 7564 8075 7616 8084
rect 7564 8041 7573 8075
rect 7573 8041 7607 8075
rect 7607 8041 7616 8075
rect 7564 8032 7616 8041
rect 8484 8075 8536 8084
rect 8484 8041 8493 8075
rect 8493 8041 8527 8075
rect 8527 8041 8536 8075
rect 8484 8032 8536 8041
rect 9956 8032 10008 8084
rect 13452 8032 13504 8084
rect 15568 8032 15620 8084
rect 8668 7964 8720 8016
rect 5080 7896 5132 7948
rect 4252 7803 4304 7812
rect 4252 7769 4261 7803
rect 4261 7769 4295 7803
rect 4295 7769 4304 7803
rect 4252 7760 4304 7769
rect 4712 7828 4764 7880
rect 7380 7896 7432 7948
rect 12164 7964 12216 8016
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 5540 7871 5592 7880
rect 5540 7837 5549 7871
rect 5549 7837 5583 7871
rect 5583 7837 5592 7871
rect 5540 7828 5592 7837
rect 5908 7828 5960 7880
rect 6368 7871 6420 7880
rect 6368 7837 6377 7871
rect 6377 7837 6411 7871
rect 6411 7837 6420 7871
rect 6368 7828 6420 7837
rect 7932 7828 7984 7880
rect 9404 7828 9456 7880
rect 12532 7939 12584 7948
rect 12532 7905 12541 7939
rect 12541 7905 12575 7939
rect 12575 7905 12584 7939
rect 12532 7896 12584 7905
rect 13452 7939 13504 7948
rect 13452 7905 13461 7939
rect 13461 7905 13495 7939
rect 13495 7905 13504 7939
rect 13452 7896 13504 7905
rect 16304 8032 16356 8084
rect 18512 8032 18564 8084
rect 16120 7964 16172 8016
rect 17040 7964 17092 8016
rect 18328 7964 18380 8016
rect 10968 7828 11020 7880
rect 11060 7828 11112 7880
rect 13912 7828 13964 7880
rect 5080 7735 5132 7744
rect 5080 7701 5089 7735
rect 5089 7701 5123 7735
rect 5123 7701 5132 7735
rect 5080 7692 5132 7701
rect 5540 7692 5592 7744
rect 6736 7760 6788 7812
rect 7012 7760 7064 7812
rect 9496 7803 9548 7812
rect 9496 7769 9505 7803
rect 9505 7769 9539 7803
rect 9539 7769 9548 7803
rect 9496 7760 9548 7769
rect 14280 7803 14332 7812
rect 14280 7769 14289 7803
rect 14289 7769 14323 7803
rect 14323 7769 14332 7803
rect 14280 7760 14332 7769
rect 14372 7760 14424 7812
rect 16120 7828 16172 7880
rect 18144 7896 18196 7948
rect 19524 7896 19576 7948
rect 16488 7871 16540 7880
rect 16488 7837 16497 7871
rect 16497 7837 16531 7871
rect 16531 7837 16540 7871
rect 16488 7828 16540 7837
rect 16948 7871 17000 7880
rect 16948 7837 16957 7871
rect 16957 7837 16991 7871
rect 16991 7837 17000 7871
rect 16948 7828 17000 7837
rect 17040 7828 17092 7880
rect 9588 7692 9640 7744
rect 10600 7692 10652 7744
rect 10692 7735 10744 7744
rect 10692 7701 10701 7735
rect 10701 7701 10735 7735
rect 10735 7701 10744 7735
rect 10692 7692 10744 7701
rect 12348 7692 12400 7744
rect 12532 7692 12584 7744
rect 15016 7803 15068 7812
rect 15016 7769 15025 7803
rect 15025 7769 15059 7803
rect 15059 7769 15068 7803
rect 15016 7760 15068 7769
rect 15108 7760 15160 7812
rect 14924 7692 14976 7744
rect 16580 7760 16632 7812
rect 18052 7871 18104 7880
rect 18052 7837 18061 7871
rect 18061 7837 18095 7871
rect 18095 7837 18104 7871
rect 18052 7828 18104 7837
rect 18420 7871 18472 7880
rect 18420 7837 18429 7871
rect 18429 7837 18463 7871
rect 18463 7837 18472 7871
rect 18420 7828 18472 7837
rect 18788 7828 18840 7880
rect 16028 7692 16080 7744
rect 6378 7590 6430 7642
rect 6442 7590 6494 7642
rect 6506 7590 6558 7642
rect 6570 7590 6622 7642
rect 6634 7590 6686 7642
rect 11806 7590 11858 7642
rect 11870 7590 11922 7642
rect 11934 7590 11986 7642
rect 11998 7590 12050 7642
rect 12062 7590 12114 7642
rect 17234 7590 17286 7642
rect 17298 7590 17350 7642
rect 17362 7590 17414 7642
rect 17426 7590 17478 7642
rect 17490 7590 17542 7642
rect 22662 7590 22714 7642
rect 22726 7590 22778 7642
rect 22790 7590 22842 7642
rect 22854 7590 22906 7642
rect 22918 7590 22970 7642
rect 4528 7488 4580 7540
rect 4896 7488 4948 7540
rect 6920 7488 6972 7540
rect 9404 7531 9456 7540
rect 9404 7497 9413 7531
rect 9413 7497 9447 7531
rect 9447 7497 9456 7531
rect 9404 7488 9456 7497
rect 10048 7488 10100 7540
rect 10600 7488 10652 7540
rect 4344 7420 4396 7472
rect 7288 7420 7340 7472
rect 3424 7352 3476 7404
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 8484 7420 8536 7472
rect 6736 7352 6788 7361
rect 7932 7352 7984 7404
rect 10692 7352 10744 7404
rect 11152 7352 11204 7404
rect 12348 7420 12400 7472
rect 13912 7420 13964 7472
rect 14280 7395 14332 7404
rect 7012 7284 7064 7336
rect 7380 7327 7432 7336
rect 7380 7293 7389 7327
rect 7389 7293 7423 7327
rect 7423 7293 7432 7327
rect 7380 7284 7432 7293
rect 7472 7284 7524 7336
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 5080 7216 5132 7268
rect 9588 7216 9640 7268
rect 12256 7284 12308 7336
rect 14004 7327 14056 7336
rect 14004 7293 14013 7327
rect 14013 7293 14047 7327
rect 14047 7293 14056 7327
rect 14004 7284 14056 7293
rect 15844 7420 15896 7472
rect 16396 7420 16448 7472
rect 16948 7420 17000 7472
rect 18052 7488 18104 7540
rect 18420 7531 18472 7540
rect 18420 7497 18429 7531
rect 18429 7497 18463 7531
rect 18463 7497 18472 7531
rect 18420 7488 18472 7497
rect 19248 7488 19300 7540
rect 16580 7352 16632 7404
rect 15016 7216 15068 7268
rect 17040 7284 17092 7336
rect 18328 7352 18380 7404
rect 19524 7420 19576 7472
rect 18788 7395 18840 7404
rect 18788 7361 18797 7395
rect 18797 7361 18831 7395
rect 18831 7361 18840 7395
rect 18788 7352 18840 7361
rect 8668 7148 8720 7200
rect 9220 7191 9272 7200
rect 9220 7157 9229 7191
rect 9229 7157 9263 7191
rect 9263 7157 9272 7191
rect 9220 7148 9272 7157
rect 12164 7148 12216 7200
rect 13452 7148 13504 7200
rect 15292 7148 15344 7200
rect 16028 7191 16080 7200
rect 16028 7157 16037 7191
rect 16037 7157 16071 7191
rect 16071 7157 16080 7191
rect 16028 7148 16080 7157
rect 3664 7046 3716 7098
rect 3728 7046 3780 7098
rect 3792 7046 3844 7098
rect 3856 7046 3908 7098
rect 3920 7046 3972 7098
rect 9092 7046 9144 7098
rect 9156 7046 9208 7098
rect 9220 7046 9272 7098
rect 9284 7046 9336 7098
rect 9348 7046 9400 7098
rect 14520 7046 14572 7098
rect 14584 7046 14636 7098
rect 14648 7046 14700 7098
rect 14712 7046 14764 7098
rect 14776 7046 14828 7098
rect 19948 7046 20000 7098
rect 20012 7046 20064 7098
rect 20076 7046 20128 7098
rect 20140 7046 20192 7098
rect 20204 7046 20256 7098
rect 5540 6944 5592 6996
rect 9772 6944 9824 6996
rect 15844 6987 15896 6996
rect 15844 6953 15853 6987
rect 15853 6953 15887 6987
rect 15887 6953 15896 6987
rect 15844 6944 15896 6953
rect 10968 6876 11020 6928
rect 18236 6876 18288 6928
rect 16120 6740 16172 6792
rect 16488 6740 16540 6792
rect 6378 6502 6430 6554
rect 6442 6502 6494 6554
rect 6506 6502 6558 6554
rect 6570 6502 6622 6554
rect 6634 6502 6686 6554
rect 11806 6502 11858 6554
rect 11870 6502 11922 6554
rect 11934 6502 11986 6554
rect 11998 6502 12050 6554
rect 12062 6502 12114 6554
rect 17234 6502 17286 6554
rect 17298 6502 17350 6554
rect 17362 6502 17414 6554
rect 17426 6502 17478 6554
rect 17490 6502 17542 6554
rect 22662 6502 22714 6554
rect 22726 6502 22778 6554
rect 22790 6502 22842 6554
rect 22854 6502 22906 6554
rect 22918 6502 22970 6554
rect 3664 5958 3716 6010
rect 3728 5958 3780 6010
rect 3792 5958 3844 6010
rect 3856 5958 3908 6010
rect 3920 5958 3972 6010
rect 9092 5958 9144 6010
rect 9156 5958 9208 6010
rect 9220 5958 9272 6010
rect 9284 5958 9336 6010
rect 9348 5958 9400 6010
rect 14520 5958 14572 6010
rect 14584 5958 14636 6010
rect 14648 5958 14700 6010
rect 14712 5958 14764 6010
rect 14776 5958 14828 6010
rect 19948 5958 20000 6010
rect 20012 5958 20064 6010
rect 20076 5958 20128 6010
rect 20140 5958 20192 6010
rect 20204 5958 20256 6010
rect 6378 5414 6430 5466
rect 6442 5414 6494 5466
rect 6506 5414 6558 5466
rect 6570 5414 6622 5466
rect 6634 5414 6686 5466
rect 11806 5414 11858 5466
rect 11870 5414 11922 5466
rect 11934 5414 11986 5466
rect 11998 5414 12050 5466
rect 12062 5414 12114 5466
rect 17234 5414 17286 5466
rect 17298 5414 17350 5466
rect 17362 5414 17414 5466
rect 17426 5414 17478 5466
rect 17490 5414 17542 5466
rect 22662 5414 22714 5466
rect 22726 5414 22778 5466
rect 22790 5414 22842 5466
rect 22854 5414 22906 5466
rect 22918 5414 22970 5466
rect 3664 4870 3716 4922
rect 3728 4870 3780 4922
rect 3792 4870 3844 4922
rect 3856 4870 3908 4922
rect 3920 4870 3972 4922
rect 9092 4870 9144 4922
rect 9156 4870 9208 4922
rect 9220 4870 9272 4922
rect 9284 4870 9336 4922
rect 9348 4870 9400 4922
rect 14520 4870 14572 4922
rect 14584 4870 14636 4922
rect 14648 4870 14700 4922
rect 14712 4870 14764 4922
rect 14776 4870 14828 4922
rect 19948 4870 20000 4922
rect 20012 4870 20064 4922
rect 20076 4870 20128 4922
rect 20140 4870 20192 4922
rect 20204 4870 20256 4922
rect 6378 4326 6430 4378
rect 6442 4326 6494 4378
rect 6506 4326 6558 4378
rect 6570 4326 6622 4378
rect 6634 4326 6686 4378
rect 11806 4326 11858 4378
rect 11870 4326 11922 4378
rect 11934 4326 11986 4378
rect 11998 4326 12050 4378
rect 12062 4326 12114 4378
rect 17234 4326 17286 4378
rect 17298 4326 17350 4378
rect 17362 4326 17414 4378
rect 17426 4326 17478 4378
rect 17490 4326 17542 4378
rect 22662 4326 22714 4378
rect 22726 4326 22778 4378
rect 22790 4326 22842 4378
rect 22854 4326 22906 4378
rect 22918 4326 22970 4378
rect 3664 3782 3716 3834
rect 3728 3782 3780 3834
rect 3792 3782 3844 3834
rect 3856 3782 3908 3834
rect 3920 3782 3972 3834
rect 9092 3782 9144 3834
rect 9156 3782 9208 3834
rect 9220 3782 9272 3834
rect 9284 3782 9336 3834
rect 9348 3782 9400 3834
rect 14520 3782 14572 3834
rect 14584 3782 14636 3834
rect 14648 3782 14700 3834
rect 14712 3782 14764 3834
rect 14776 3782 14828 3834
rect 19948 3782 20000 3834
rect 20012 3782 20064 3834
rect 20076 3782 20128 3834
rect 20140 3782 20192 3834
rect 20204 3782 20256 3834
rect 6378 3238 6430 3290
rect 6442 3238 6494 3290
rect 6506 3238 6558 3290
rect 6570 3238 6622 3290
rect 6634 3238 6686 3290
rect 11806 3238 11858 3290
rect 11870 3238 11922 3290
rect 11934 3238 11986 3290
rect 11998 3238 12050 3290
rect 12062 3238 12114 3290
rect 17234 3238 17286 3290
rect 17298 3238 17350 3290
rect 17362 3238 17414 3290
rect 17426 3238 17478 3290
rect 17490 3238 17542 3290
rect 22662 3238 22714 3290
rect 22726 3238 22778 3290
rect 22790 3238 22842 3290
rect 22854 3238 22906 3290
rect 22918 3238 22970 3290
rect 3664 2694 3716 2746
rect 3728 2694 3780 2746
rect 3792 2694 3844 2746
rect 3856 2694 3908 2746
rect 3920 2694 3972 2746
rect 9092 2694 9144 2746
rect 9156 2694 9208 2746
rect 9220 2694 9272 2746
rect 9284 2694 9336 2746
rect 9348 2694 9400 2746
rect 14520 2694 14572 2746
rect 14584 2694 14636 2746
rect 14648 2694 14700 2746
rect 14712 2694 14764 2746
rect 14776 2694 14828 2746
rect 19948 2694 20000 2746
rect 20012 2694 20064 2746
rect 20076 2694 20128 2746
rect 20140 2694 20192 2746
rect 20204 2694 20256 2746
rect 10876 2592 10928 2644
rect 6092 2524 6144 2576
rect 8852 2456 8904 2508
rect 4988 2388 5040 2440
rect 5908 2388 5960 2440
rect 8392 2388 8444 2440
rect 8576 2388 8628 2440
rect 20996 2431 21048 2440
rect 20996 2397 21005 2431
rect 21005 2397 21039 2431
rect 21039 2397 21048 2431
rect 20996 2388 21048 2397
rect 1676 2320 1728 2372
rect 4620 2320 4672 2372
rect 7564 2320 7616 2372
rect 10508 2320 10560 2372
rect 13820 2320 13872 2372
rect 16580 2320 16632 2372
rect 19340 2320 19392 2372
rect 22284 2320 22336 2372
rect 6378 2150 6430 2202
rect 6442 2150 6494 2202
rect 6506 2150 6558 2202
rect 6570 2150 6622 2202
rect 6634 2150 6686 2202
rect 11806 2150 11858 2202
rect 11870 2150 11922 2202
rect 11934 2150 11986 2202
rect 11998 2150 12050 2202
rect 12062 2150 12114 2202
rect 17234 2150 17286 2202
rect 17298 2150 17350 2202
rect 17362 2150 17414 2202
rect 17426 2150 17478 2202
rect 17490 2150 17542 2202
rect 22662 2150 22714 2202
rect 22726 2150 22778 2202
rect 22790 2150 22842 2202
rect 22854 2150 22906 2202
rect 22918 2150 22970 2202
<< metal2 >>
rect 3974 23338 4030 24000
rect 11978 23338 12034 24000
rect 3974 23310 4108 23338
rect 3974 23200 4030 23310
rect 1860 21344 1912 21350
rect 1860 21286 1912 21292
rect 1872 20602 1900 21286
rect 3664 21244 3972 21253
rect 3664 21242 3670 21244
rect 3726 21242 3750 21244
rect 3806 21242 3830 21244
rect 3886 21242 3910 21244
rect 3966 21242 3972 21244
rect 3726 21190 3728 21242
rect 3908 21190 3910 21242
rect 3664 21188 3670 21190
rect 3726 21188 3750 21190
rect 3806 21188 3830 21190
rect 3886 21188 3910 21190
rect 3966 21188 3972 21190
rect 3664 21179 3972 21188
rect 2964 21004 3016 21010
rect 2964 20946 3016 20952
rect 2976 20874 3004 20946
rect 2688 20868 2740 20874
rect 2688 20810 2740 20816
rect 2964 20868 3016 20874
rect 2964 20810 3016 20816
rect 1860 20596 1912 20602
rect 1860 20538 1912 20544
rect 1768 20460 1820 20466
rect 1768 20402 1820 20408
rect 1780 19990 1808 20402
rect 1768 19984 1820 19990
rect 1768 19926 1820 19932
rect 1872 19922 1900 20538
rect 2700 20330 2728 20810
rect 2976 20602 3004 20810
rect 3976 20800 4028 20806
rect 3976 20742 4028 20748
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 2688 20324 2740 20330
rect 2688 20266 2740 20272
rect 2228 20256 2280 20262
rect 2228 20198 2280 20204
rect 1860 19916 1912 19922
rect 1860 19858 1912 19864
rect 1872 19378 1900 19858
rect 2240 19854 2268 20198
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 2504 19780 2556 19786
rect 2504 19722 2556 19728
rect 2412 19712 2464 19718
rect 2412 19654 2464 19660
rect 2424 19446 2452 19654
rect 2412 19440 2464 19446
rect 2412 19382 2464 19388
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 2516 19258 2544 19722
rect 2700 19378 2728 20266
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 2884 19854 2912 20198
rect 2872 19848 2924 19854
rect 2872 19790 2924 19796
rect 2976 19786 3004 20538
rect 3056 20460 3108 20466
rect 3056 20402 3108 20408
rect 3068 20058 3096 20402
rect 3988 20262 4016 20742
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3664 20156 3972 20165
rect 3664 20154 3670 20156
rect 3726 20154 3750 20156
rect 3806 20154 3830 20156
rect 3886 20154 3910 20156
rect 3966 20154 3972 20156
rect 3726 20102 3728 20154
rect 3908 20102 3910 20154
rect 3664 20100 3670 20102
rect 3726 20100 3750 20102
rect 3806 20100 3830 20102
rect 3886 20100 3910 20102
rect 3966 20100 3972 20102
rect 3664 20091 3972 20100
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 2964 19780 3016 19786
rect 2964 19722 3016 19728
rect 4080 19718 4108 23310
rect 11978 23310 12204 23338
rect 11978 23200 12034 23310
rect 6378 21788 6686 21797
rect 6378 21786 6384 21788
rect 6440 21786 6464 21788
rect 6520 21786 6544 21788
rect 6600 21786 6624 21788
rect 6680 21786 6686 21788
rect 6440 21734 6442 21786
rect 6622 21734 6624 21786
rect 6378 21732 6384 21734
rect 6440 21732 6464 21734
rect 6520 21732 6544 21734
rect 6600 21732 6624 21734
rect 6680 21732 6686 21734
rect 6378 21723 6686 21732
rect 11806 21788 12114 21797
rect 11806 21786 11812 21788
rect 11868 21786 11892 21788
rect 11948 21786 11972 21788
rect 12028 21786 12052 21788
rect 12108 21786 12114 21788
rect 11868 21734 11870 21786
rect 12050 21734 12052 21786
rect 11806 21732 11812 21734
rect 11868 21732 11892 21734
rect 11948 21732 11972 21734
rect 12028 21732 12052 21734
rect 12108 21732 12114 21734
rect 11806 21723 12114 21732
rect 12176 21622 12204 23310
rect 19982 23200 20038 24000
rect 17234 21788 17542 21797
rect 17234 21786 17240 21788
rect 17296 21786 17320 21788
rect 17376 21786 17400 21788
rect 17456 21786 17480 21788
rect 17536 21786 17542 21788
rect 17296 21734 17298 21786
rect 17478 21734 17480 21786
rect 17234 21732 17240 21734
rect 17296 21732 17320 21734
rect 17376 21732 17400 21734
rect 17456 21732 17480 21734
rect 17536 21732 17542 21734
rect 17234 21723 17542 21732
rect 19996 21622 20024 23200
rect 22662 21788 22970 21797
rect 22662 21786 22668 21788
rect 22724 21786 22748 21788
rect 22804 21786 22828 21788
rect 22884 21786 22908 21788
rect 22964 21786 22970 21788
rect 22724 21734 22726 21786
rect 22906 21734 22908 21786
rect 22662 21732 22668 21734
rect 22724 21732 22748 21734
rect 22804 21732 22828 21734
rect 22884 21732 22908 21734
rect 22964 21732 22970 21734
rect 22662 21723 22970 21732
rect 12164 21616 12216 21622
rect 12164 21558 12216 21564
rect 16488 21616 16540 21622
rect 16488 21558 16540 21564
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 16396 21548 16448 21554
rect 16396 21490 16448 21496
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 15384 21412 15436 21418
rect 15384 21354 15436 21360
rect 10232 21344 10284 21350
rect 10232 21286 10284 21292
rect 9092 21244 9400 21253
rect 9092 21242 9098 21244
rect 9154 21242 9178 21244
rect 9234 21242 9258 21244
rect 9314 21242 9338 21244
rect 9394 21242 9400 21244
rect 9154 21190 9156 21242
rect 9336 21190 9338 21242
rect 9092 21188 9098 21190
rect 9154 21188 9178 21190
rect 9234 21188 9258 21190
rect 9314 21188 9338 21190
rect 9394 21188 9400 21190
rect 9092 21179 9400 21188
rect 10244 21078 10272 21286
rect 14520 21244 14828 21253
rect 14520 21242 14526 21244
rect 14582 21242 14606 21244
rect 14662 21242 14686 21244
rect 14742 21242 14766 21244
rect 14822 21242 14828 21244
rect 14582 21190 14584 21242
rect 14764 21190 14766 21242
rect 14520 21188 14526 21190
rect 14582 21188 14606 21190
rect 14662 21188 14686 21190
rect 14742 21188 14766 21190
rect 14822 21188 14828 21190
rect 14520 21179 14828 21188
rect 10232 21072 10284 21078
rect 10232 21014 10284 21020
rect 13820 21072 13872 21078
rect 13820 21014 13872 21020
rect 6000 20936 6052 20942
rect 6000 20878 6052 20884
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 4252 20868 4304 20874
rect 4252 20810 4304 20816
rect 4264 20602 4292 20810
rect 4252 20596 4304 20602
rect 4252 20538 4304 20544
rect 6012 20398 6040 20878
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6378 20700 6686 20709
rect 6378 20698 6384 20700
rect 6440 20698 6464 20700
rect 6520 20698 6544 20700
rect 6600 20698 6624 20700
rect 6680 20698 6686 20700
rect 6440 20646 6442 20698
rect 6622 20646 6624 20698
rect 6378 20644 6384 20646
rect 6440 20644 6464 20646
rect 6520 20644 6544 20646
rect 6600 20644 6624 20646
rect 6680 20644 6686 20646
rect 6378 20635 6686 20644
rect 6932 20534 6960 20742
rect 6920 20528 6972 20534
rect 6920 20470 6972 20476
rect 7024 20466 7052 20878
rect 9128 20868 9180 20874
rect 9128 20810 9180 20816
rect 9312 20868 9364 20874
rect 9312 20810 9364 20816
rect 9140 20602 9168 20810
rect 9128 20596 9180 20602
rect 9128 20538 9180 20544
rect 9324 20466 9352 20810
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 9968 20534 9996 20742
rect 11806 20700 12114 20709
rect 11806 20698 11812 20700
rect 11868 20698 11892 20700
rect 11948 20698 11972 20700
rect 12028 20698 12052 20700
rect 12108 20698 12114 20700
rect 11868 20646 11870 20698
rect 12050 20646 12052 20698
rect 11806 20644 11812 20646
rect 11868 20644 11892 20646
rect 11948 20644 11972 20646
rect 12028 20644 12052 20646
rect 12108 20644 12114 20646
rect 11806 20635 12114 20644
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 7012 20460 7064 20466
rect 7012 20402 7064 20408
rect 9312 20460 9364 20466
rect 9312 20402 9364 20408
rect 6000 20392 6052 20398
rect 6000 20334 6052 20340
rect 6012 19854 6040 20334
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 4528 19780 4580 19786
rect 4528 19722 4580 19728
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 2424 19230 2544 19258
rect 1860 18216 1912 18222
rect 1860 18158 1912 18164
rect 1872 17678 1900 18158
rect 1860 17672 1912 17678
rect 1860 17614 1912 17620
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17338 1992 17478
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 1964 16658 1992 17274
rect 2332 17202 2360 17614
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 2424 16574 2452 19230
rect 2700 18766 2728 19314
rect 3664 19068 3972 19077
rect 3664 19066 3670 19068
rect 3726 19066 3750 19068
rect 3806 19066 3830 19068
rect 3886 19066 3910 19068
rect 3966 19066 3972 19068
rect 3726 19014 3728 19066
rect 3908 19014 3910 19066
rect 3664 19012 3670 19014
rect 3726 19012 3750 19014
rect 3806 19012 3830 19014
rect 3886 19012 3910 19014
rect 3966 19012 3972 19014
rect 3664 19003 3972 19012
rect 4540 18970 4568 19722
rect 6012 19378 6040 19790
rect 6378 19612 6686 19621
rect 6378 19610 6384 19612
rect 6440 19610 6464 19612
rect 6520 19610 6544 19612
rect 6600 19610 6624 19612
rect 6680 19610 6686 19612
rect 6440 19558 6442 19610
rect 6622 19558 6624 19610
rect 6378 19556 6384 19558
rect 6440 19556 6464 19558
rect 6520 19556 6544 19558
rect 6600 19556 6624 19558
rect 6680 19556 6686 19558
rect 6378 19547 6686 19556
rect 7024 19378 7052 20402
rect 12176 20398 12204 20878
rect 13832 20602 13860 21014
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 15396 20466 15424 21354
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 9496 20392 9548 20398
rect 9496 20334 9548 20340
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 9092 20156 9400 20165
rect 9092 20154 9098 20156
rect 9154 20154 9178 20156
rect 9234 20154 9258 20156
rect 9314 20154 9338 20156
rect 9394 20154 9400 20156
rect 9154 20102 9156 20154
rect 9336 20102 9338 20154
rect 9092 20100 9098 20102
rect 9154 20100 9178 20102
rect 9234 20100 9258 20102
rect 9314 20100 9338 20102
rect 9394 20100 9400 20102
rect 9092 20091 9400 20100
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4528 18964 4580 18970
rect 4528 18906 4580 18912
rect 4632 18766 4660 19110
rect 6012 18834 6040 19314
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 2688 18760 2740 18766
rect 2688 18702 2740 18708
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 2700 18358 2728 18702
rect 4068 18692 4120 18698
rect 4068 18634 4120 18640
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 3436 18358 3464 18566
rect 4080 18426 4108 18634
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 2688 18352 2740 18358
rect 2688 18294 2740 18300
rect 3424 18352 3476 18358
rect 3424 18294 3476 18300
rect 2596 18148 2648 18154
rect 2596 18090 2648 18096
rect 2504 17604 2556 17610
rect 2504 17546 2556 17552
rect 2516 17134 2544 17546
rect 2608 17542 2636 18090
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2504 17128 2556 17134
rect 2504 17070 2556 17076
rect 2056 16546 2452 16574
rect 1768 16516 1820 16522
rect 1768 16458 1820 16464
rect 1780 16250 1808 16458
rect 1768 16244 1820 16250
rect 1768 16186 1820 16192
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 1964 12238 1992 15438
rect 2056 13938 2084 16546
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2424 16250 2452 16390
rect 2412 16244 2464 16250
rect 2412 16186 2464 16192
rect 2320 16176 2372 16182
rect 2320 16118 2372 16124
rect 2136 16040 2188 16046
rect 2136 15982 2188 15988
rect 2148 15706 2176 15982
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2148 14550 2176 15642
rect 2332 15570 2360 16118
rect 2516 16114 2544 17070
rect 2608 16182 2636 17478
rect 2596 16176 2648 16182
rect 2596 16118 2648 16124
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2516 15638 2544 16050
rect 2700 15978 2728 18294
rect 6012 18290 6040 18770
rect 8116 18760 8168 18766
rect 8116 18702 8168 18708
rect 6378 18524 6686 18533
rect 6378 18522 6384 18524
rect 6440 18522 6464 18524
rect 6520 18522 6544 18524
rect 6600 18522 6624 18524
rect 6680 18522 6686 18524
rect 6440 18470 6442 18522
rect 6622 18470 6624 18522
rect 6378 18468 6384 18470
rect 6440 18468 6464 18470
rect 6520 18468 6544 18470
rect 6600 18468 6624 18470
rect 6680 18468 6686 18470
rect 6378 18459 6686 18468
rect 8128 18290 8156 18702
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 6000 18284 6052 18290
rect 6000 18226 6052 18232
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2884 17338 2912 17478
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 3068 17202 3096 17614
rect 3252 17202 3280 18022
rect 3664 17980 3972 17989
rect 3664 17978 3670 17980
rect 3726 17978 3750 17980
rect 3806 17978 3830 17980
rect 3886 17978 3910 17980
rect 3966 17978 3972 17980
rect 3726 17926 3728 17978
rect 3908 17926 3910 17978
rect 3664 17924 3670 17926
rect 3726 17924 3750 17926
rect 3806 17924 3830 17926
rect 3886 17924 3910 17926
rect 3966 17924 3972 17926
rect 3664 17915 3972 17924
rect 4632 17882 4660 18226
rect 6012 17882 6040 18226
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 6012 17202 6040 17818
rect 6378 17436 6686 17445
rect 6378 17434 6384 17436
rect 6440 17434 6464 17436
rect 6520 17434 6544 17436
rect 6600 17434 6624 17436
rect 6680 17434 6686 17436
rect 6440 17382 6442 17434
rect 6622 17382 6624 17434
rect 6378 17380 6384 17382
rect 6440 17380 6464 17382
rect 6520 17380 6544 17382
rect 6600 17380 6624 17382
rect 6680 17380 6686 17382
rect 6378 17371 6686 17380
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 2504 15632 2556 15638
rect 2504 15574 2556 15580
rect 2320 15564 2372 15570
rect 2320 15506 2372 15512
rect 2332 15042 2360 15506
rect 2516 15162 2544 15574
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2504 15156 2556 15162
rect 2504 15098 2556 15104
rect 2240 15026 2452 15042
rect 2240 15020 2464 15026
rect 2240 15014 2412 15020
rect 2240 14618 2268 15014
rect 2412 14962 2464 14968
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 2516 14414 2544 15098
rect 2608 15094 2636 15506
rect 2700 15502 2728 15914
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2884 15162 2912 16050
rect 2976 15978 3004 16186
rect 2964 15972 3016 15978
rect 2964 15914 3016 15920
rect 3068 15570 3096 17138
rect 3148 16992 3200 16998
rect 3148 16934 3200 16940
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 3160 16590 3188 16934
rect 3664 16892 3972 16901
rect 3664 16890 3670 16892
rect 3726 16890 3750 16892
rect 3806 16890 3830 16892
rect 3886 16890 3910 16892
rect 3966 16890 3972 16892
rect 3726 16838 3728 16890
rect 3908 16838 3910 16890
rect 3664 16836 3670 16838
rect 3726 16836 3750 16838
rect 3806 16836 3830 16838
rect 3886 16836 3910 16838
rect 3966 16836 3972 16838
rect 3664 16827 3972 16836
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3160 16182 3188 16526
rect 3252 16250 3280 16526
rect 3896 16454 3924 16526
rect 3884 16448 3936 16454
rect 3884 16390 3936 16396
rect 3240 16244 3292 16250
rect 3240 16186 3292 16192
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 3148 16176 3200 16182
rect 3148 16118 3200 16124
rect 3664 15804 3972 15813
rect 3664 15802 3670 15804
rect 3726 15802 3750 15804
rect 3806 15802 3830 15804
rect 3886 15802 3910 15804
rect 3966 15802 3972 15804
rect 3726 15750 3728 15802
rect 3908 15750 3910 15802
rect 3664 15748 3670 15750
rect 3726 15748 3750 15750
rect 3806 15748 3830 15750
rect 3886 15748 3910 15750
rect 3966 15748 3972 15750
rect 3664 15739 3972 15748
rect 4080 15570 4108 16186
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 2596 15088 2648 15094
rect 2596 15030 2648 15036
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 3528 14074 3556 14962
rect 3664 14716 3972 14725
rect 3664 14714 3670 14716
rect 3726 14714 3750 14716
rect 3806 14714 3830 14716
rect 3886 14714 3910 14716
rect 3966 14714 3972 14716
rect 3726 14662 3728 14714
rect 3908 14662 3910 14714
rect 3664 14660 3670 14662
rect 3726 14660 3750 14662
rect 3806 14660 3830 14662
rect 3886 14660 3910 14662
rect 3966 14660 3972 14662
rect 3664 14651 3972 14660
rect 4080 14618 4108 14962
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4620 14340 4672 14346
rect 4620 14282 4672 14288
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 2056 10742 2084 13874
rect 3664 13628 3972 13637
rect 3664 13626 3670 13628
rect 3726 13626 3750 13628
rect 3806 13626 3830 13628
rect 3886 13626 3910 13628
rect 3966 13626 3972 13628
rect 3726 13574 3728 13626
rect 3908 13574 3910 13626
rect 3664 13572 3670 13574
rect 3726 13572 3750 13574
rect 3806 13572 3830 13574
rect 3886 13572 3910 13574
rect 3966 13572 3972 13574
rect 3664 13563 3972 13572
rect 3664 12540 3972 12549
rect 3664 12538 3670 12540
rect 3726 12538 3750 12540
rect 3806 12538 3830 12540
rect 3886 12538 3910 12540
rect 3966 12538 3972 12540
rect 3726 12486 3728 12538
rect 3908 12486 3910 12538
rect 3664 12484 3670 12486
rect 3726 12484 3750 12486
rect 3806 12484 3830 12486
rect 3886 12484 3910 12486
rect 3966 12484 3972 12486
rect 3664 12475 3972 12484
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2044 10736 2096 10742
rect 2044 10678 2096 10684
rect 2044 10532 2096 10538
rect 2044 10474 2096 10480
rect 1860 9988 1912 9994
rect 1860 9930 1912 9936
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1780 9586 1808 9862
rect 1872 9722 1900 9930
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 2056 9450 2084 10474
rect 2240 9722 2268 12174
rect 2608 11898 2636 12174
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2792 11898 2820 12106
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 3160 11762 3188 12242
rect 4172 12186 4200 14214
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4264 12434 4292 12786
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4264 12406 4384 12434
rect 4172 12158 4292 12186
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4172 11830 4200 12038
rect 4160 11824 4212 11830
rect 4160 11766 4212 11772
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2608 10810 2636 11630
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2332 10266 2360 10610
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2412 10192 2464 10198
rect 2412 10134 2464 10140
rect 2228 9716 2280 9722
rect 2228 9658 2280 9664
rect 2424 9654 2452 10134
rect 2412 9648 2464 9654
rect 2412 9590 2464 9596
rect 2044 9444 2096 9450
rect 2044 9386 2096 9392
rect 2424 9178 2452 9590
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2608 9042 2636 10746
rect 2700 10266 2728 11698
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2700 10130 2728 10202
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 3160 9926 3188 11698
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 3664 11452 3972 11461
rect 3664 11450 3670 11452
rect 3726 11450 3750 11452
rect 3806 11450 3830 11452
rect 3886 11450 3910 11452
rect 3966 11450 3972 11452
rect 3726 11398 3728 11450
rect 3908 11398 3910 11450
rect 3664 11396 3670 11398
rect 3726 11396 3750 11398
rect 3806 11396 3830 11398
rect 3886 11396 3910 11398
rect 3966 11396 3972 11398
rect 3664 11387 3972 11396
rect 4172 10742 4200 11630
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3528 10198 3556 10610
rect 3664 10364 3972 10373
rect 3664 10362 3670 10364
rect 3726 10362 3750 10364
rect 3806 10362 3830 10364
rect 3886 10362 3910 10364
rect 3966 10362 3972 10364
rect 3726 10310 3728 10362
rect 3908 10310 3910 10362
rect 3664 10308 3670 10310
rect 3726 10308 3750 10310
rect 3806 10308 3830 10310
rect 3886 10308 3910 10310
rect 3966 10308 3972 10310
rect 3664 10299 3972 10308
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 4160 10124 4212 10130
rect 4264 10112 4292 12158
rect 4356 10810 4384 12406
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4448 10674 4476 12582
rect 4436 10668 4488 10674
rect 4436 10610 4488 10616
rect 4212 10084 4292 10112
rect 4160 10066 4212 10072
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 3160 8498 3188 9862
rect 3664 9276 3972 9285
rect 3664 9274 3670 9276
rect 3726 9274 3750 9276
rect 3806 9274 3830 9276
rect 3886 9274 3910 9276
rect 3966 9274 3972 9276
rect 3726 9222 3728 9274
rect 3908 9222 3910 9274
rect 3664 9220 3670 9222
rect 3726 9220 3750 9222
rect 3806 9220 3830 9222
rect 3886 9220 3910 9222
rect 3966 9220 3972 9222
rect 3664 9211 3972 9220
rect 4264 8974 4292 10084
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4356 9042 4384 9998
rect 4448 9926 4476 10610
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4172 8498 4200 8774
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3424 8356 3476 8362
rect 3424 8298 3476 8304
rect 3436 8090 3464 8298
rect 3528 8090 3556 8434
rect 3664 8188 3972 8197
rect 3664 8186 3670 8188
rect 3726 8186 3750 8188
rect 3806 8186 3830 8188
rect 3886 8186 3910 8188
rect 3966 8186 3972 8188
rect 3726 8134 3728 8186
rect 3908 8134 3910 8186
rect 3664 8132 3670 8134
rect 3726 8132 3750 8134
rect 3806 8132 3830 8134
rect 3886 8132 3910 8134
rect 3966 8132 3972 8134
rect 3664 8123 3972 8132
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3436 7410 3464 8026
rect 4172 7886 4200 8434
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4264 7818 4292 8026
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 4356 7478 4384 8502
rect 4540 7546 4568 13874
rect 4632 8634 4660 14282
rect 4710 10024 4766 10033
rect 4710 9959 4712 9968
rect 4764 9959 4766 9968
rect 4712 9930 4764 9936
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4724 7886 4752 8366
rect 4908 8090 4936 8434
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4908 7546 4936 8026
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3664 7100 3972 7109
rect 3664 7098 3670 7100
rect 3726 7098 3750 7100
rect 3806 7098 3830 7100
rect 3886 7098 3910 7100
rect 3966 7098 3972 7100
rect 3726 7046 3728 7098
rect 3908 7046 3910 7098
rect 3664 7044 3670 7046
rect 3726 7044 3750 7046
rect 3806 7044 3830 7046
rect 3886 7044 3910 7046
rect 3966 7044 3972 7046
rect 3664 7035 3972 7044
rect 3664 6012 3972 6021
rect 3664 6010 3670 6012
rect 3726 6010 3750 6012
rect 3806 6010 3830 6012
rect 3886 6010 3910 6012
rect 3966 6010 3972 6012
rect 3726 5958 3728 6010
rect 3908 5958 3910 6010
rect 3664 5956 3670 5958
rect 3726 5956 3750 5958
rect 3806 5956 3830 5958
rect 3886 5956 3910 5958
rect 3966 5956 3972 5958
rect 3664 5947 3972 5956
rect 3664 4924 3972 4933
rect 3664 4922 3670 4924
rect 3726 4922 3750 4924
rect 3806 4922 3830 4924
rect 3886 4922 3910 4924
rect 3966 4922 3972 4924
rect 3726 4870 3728 4922
rect 3908 4870 3910 4922
rect 3664 4868 3670 4870
rect 3726 4868 3750 4870
rect 3806 4868 3830 4870
rect 3886 4868 3910 4870
rect 3966 4868 3972 4870
rect 3664 4859 3972 4868
rect 3664 3836 3972 3845
rect 3664 3834 3670 3836
rect 3726 3834 3750 3836
rect 3806 3834 3830 3836
rect 3886 3834 3910 3836
rect 3966 3834 3972 3836
rect 3726 3782 3728 3834
rect 3908 3782 3910 3834
rect 3664 3780 3670 3782
rect 3726 3780 3750 3782
rect 3806 3780 3830 3782
rect 3886 3780 3910 3782
rect 3966 3780 3972 3782
rect 3664 3771 3972 3780
rect 3664 2748 3972 2757
rect 3664 2746 3670 2748
rect 3726 2746 3750 2748
rect 3806 2746 3830 2748
rect 3886 2746 3910 2748
rect 3966 2746 3972 2748
rect 3726 2694 3728 2746
rect 3908 2694 3910 2746
rect 3664 2692 3670 2694
rect 3726 2692 3750 2694
rect 3806 2692 3830 2694
rect 3886 2692 3910 2694
rect 3966 2692 3972 2694
rect 3664 2683 3972 2692
rect 5000 2446 5028 16934
rect 6012 16794 6040 17138
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 7024 16658 7052 17138
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 5816 16448 5868 16454
rect 5816 16390 5868 16396
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5644 14414 5672 14758
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5644 14006 5672 14350
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 5644 13530 5672 13942
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5644 12850 5672 13466
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5644 12730 5672 12786
rect 5552 12702 5672 12730
rect 5552 12220 5580 12702
rect 5736 12594 5764 13670
rect 5644 12566 5764 12594
rect 5644 12322 5672 12566
rect 5722 12472 5778 12481
rect 5722 12407 5724 12416
rect 5776 12407 5778 12416
rect 5724 12378 5776 12384
rect 5644 12294 5764 12322
rect 5632 12232 5684 12238
rect 5552 12192 5632 12220
rect 5632 12174 5684 12180
rect 5644 11830 5672 12174
rect 5632 11824 5684 11830
rect 5632 11766 5684 11772
rect 5644 11218 5672 11766
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5736 11098 5764 12294
rect 5552 11070 5764 11098
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 7954 5120 8230
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 5460 7886 5488 8978
rect 5552 7886 5580 11070
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5644 10266 5672 10746
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5644 9994 5672 10202
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5644 9654 5672 9930
rect 5736 9722 5764 9998
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5552 7750 5580 7822
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5092 7274 5120 7686
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 5552 7002 5580 7686
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5828 2774 5856 16390
rect 6378 16348 6686 16357
rect 6378 16346 6384 16348
rect 6440 16346 6464 16348
rect 6520 16346 6544 16348
rect 6600 16346 6624 16348
rect 6680 16346 6686 16348
rect 6440 16294 6442 16346
rect 6622 16294 6624 16346
rect 6378 16292 6384 16294
rect 6440 16292 6464 16294
rect 6520 16292 6544 16294
rect 6600 16292 6624 16294
rect 6680 16292 6686 16294
rect 6378 16283 6686 16292
rect 7484 15978 7512 17138
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 6378 15260 6686 15269
rect 6378 15258 6384 15260
rect 6440 15258 6464 15260
rect 6520 15258 6544 15260
rect 6600 15258 6624 15260
rect 6680 15258 6686 15260
rect 6440 15206 6442 15258
rect 6622 15206 6624 15258
rect 6378 15204 6384 15206
rect 6440 15204 6464 15206
rect 6520 15204 6544 15206
rect 6600 15204 6624 15206
rect 6680 15204 6686 15206
rect 6378 15195 6686 15204
rect 8128 15162 8156 18226
rect 8312 16182 8340 19654
rect 9508 19310 9536 20334
rect 12176 19854 12204 20334
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 9772 19372 9824 19378
rect 9692 19332 9772 19360
rect 9496 19304 9548 19310
rect 9496 19246 9548 19252
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8404 18766 8432 19110
rect 9092 19068 9400 19077
rect 9092 19066 9098 19068
rect 9154 19066 9178 19068
rect 9234 19066 9258 19068
rect 9314 19066 9338 19068
rect 9394 19066 9400 19068
rect 9154 19014 9156 19066
rect 9336 19014 9338 19066
rect 9092 19012 9098 19014
rect 9154 19012 9178 19014
rect 9234 19012 9258 19014
rect 9314 19012 9338 19014
rect 9394 19012 9400 19014
rect 9092 19003 9400 19012
rect 9508 18850 9536 19246
rect 9692 18970 9720 19332
rect 9772 19314 9824 19320
rect 11716 19310 11744 19790
rect 11806 19612 12114 19621
rect 11806 19610 11812 19612
rect 11868 19610 11892 19612
rect 11948 19610 11972 19612
rect 12028 19610 12052 19612
rect 12108 19610 12114 19612
rect 11868 19558 11870 19610
rect 12050 19558 12052 19610
rect 11806 19556 11812 19558
rect 11868 19556 11892 19558
rect 11948 19556 11972 19558
rect 12028 19556 12052 19558
rect 12108 19556 12114 19558
rect 11806 19547 12114 19556
rect 13372 19446 13400 19790
rect 14384 19786 14412 20402
rect 15200 20324 15252 20330
rect 15200 20266 15252 20272
rect 14520 20156 14828 20165
rect 14520 20154 14526 20156
rect 14582 20154 14606 20156
rect 14662 20154 14686 20156
rect 14742 20154 14766 20156
rect 14822 20154 14828 20156
rect 14582 20102 14584 20154
rect 14764 20102 14766 20154
rect 14520 20100 14526 20102
rect 14582 20100 14606 20102
rect 14662 20100 14686 20102
rect 14742 20100 14766 20102
rect 14822 20100 14828 20102
rect 14520 20091 14828 20100
rect 15212 19786 15240 20266
rect 14280 19780 14332 19786
rect 14280 19722 14332 19728
rect 14372 19780 14424 19786
rect 14372 19722 14424 19728
rect 15200 19780 15252 19786
rect 15200 19722 15252 19728
rect 13360 19440 13412 19446
rect 13360 19382 13412 19388
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9508 18822 9628 18850
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 9600 18630 9628 18822
rect 11716 18766 11744 19246
rect 13556 18834 13584 19382
rect 14292 19242 14320 19722
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14520 19068 14828 19077
rect 14520 19066 14526 19068
rect 14582 19066 14606 19068
rect 14662 19066 14686 19068
rect 14742 19066 14766 19068
rect 14822 19066 14828 19068
rect 14582 19014 14584 19066
rect 14764 19014 14766 19066
rect 14520 19012 14526 19014
rect 14582 19012 14606 19014
rect 14662 19012 14686 19014
rect 14742 19012 14766 19014
rect 14822 19012 14828 19014
rect 14520 19003 14828 19012
rect 15120 18970 15148 19654
rect 15108 18964 15160 18970
rect 15108 18906 15160 18912
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 9092 17980 9400 17989
rect 9092 17978 9098 17980
rect 9154 17978 9178 17980
rect 9234 17978 9258 17980
rect 9314 17978 9338 17980
rect 9394 17978 9400 17980
rect 9154 17926 9156 17978
rect 9336 17926 9338 17978
rect 9092 17924 9098 17926
rect 9154 17924 9178 17926
rect 9234 17924 9258 17926
rect 9314 17924 9338 17926
rect 9394 17924 9400 17926
rect 9092 17915 9400 17924
rect 9600 17898 9628 18566
rect 9600 17882 9720 17898
rect 11716 17882 11744 18702
rect 11806 18524 12114 18533
rect 11806 18522 11812 18524
rect 11868 18522 11892 18524
rect 11948 18522 11972 18524
rect 12028 18522 12052 18524
rect 12108 18522 12114 18524
rect 11868 18470 11870 18522
rect 12050 18470 12052 18522
rect 11806 18468 11812 18470
rect 11868 18468 11892 18470
rect 11948 18468 11972 18470
rect 12028 18468 12052 18470
rect 12108 18468 12114 18470
rect 11806 18459 12114 18468
rect 15304 18426 15332 18702
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 9600 17876 9732 17882
rect 9600 17870 9680 17876
rect 9680 17818 9732 17824
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 9692 17134 9720 17818
rect 10600 17604 10652 17610
rect 10600 17546 10652 17552
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8300 16176 8352 16182
rect 8300 16118 8352 16124
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5920 12481 5948 14214
rect 5906 12472 5962 12481
rect 5906 12407 5962 12416
rect 6012 12434 6040 14758
rect 7564 14340 7616 14346
rect 7564 14282 7616 14288
rect 6378 14172 6686 14181
rect 6378 14170 6384 14172
rect 6440 14170 6464 14172
rect 6520 14170 6544 14172
rect 6600 14170 6624 14172
rect 6680 14170 6686 14172
rect 6440 14118 6442 14170
rect 6622 14118 6624 14170
rect 6378 14116 6384 14118
rect 6440 14116 6464 14118
rect 6520 14116 6544 14118
rect 6600 14116 6624 14118
rect 6680 14116 6686 14118
rect 6378 14107 6686 14116
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6378 13084 6686 13093
rect 6378 13082 6384 13084
rect 6440 13082 6464 13084
rect 6520 13082 6544 13084
rect 6600 13082 6624 13084
rect 6680 13082 6686 13084
rect 6440 13030 6442 13082
rect 6622 13030 6624 13082
rect 6378 13028 6384 13030
rect 6440 13028 6464 13030
rect 6520 13028 6544 13030
rect 6600 13028 6624 13030
rect 6680 13028 6686 13030
rect 6378 13019 6686 13028
rect 6184 12436 6236 12442
rect 6012 12406 6132 12434
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 5908 11076 5960 11082
rect 5908 11018 5960 11024
rect 5920 10577 5948 11018
rect 5906 10568 5962 10577
rect 5906 10503 5962 10512
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5920 10062 5948 10406
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 6012 8906 6040 11494
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5920 7886 5948 8434
rect 6012 8430 6040 8842
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5828 2746 5948 2774
rect 5920 2446 5948 2746
rect 6104 2582 6132 12406
rect 6184 12378 6236 12384
rect 6196 10656 6224 12378
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6378 11996 6686 12005
rect 6378 11994 6384 11996
rect 6440 11994 6464 11996
rect 6520 11994 6544 11996
rect 6600 11994 6624 11996
rect 6680 11994 6686 11996
rect 6440 11942 6442 11994
rect 6622 11942 6624 11994
rect 6378 11940 6384 11942
rect 6440 11940 6464 11942
rect 6520 11940 6544 11942
rect 6600 11940 6624 11942
rect 6680 11940 6686 11942
rect 6378 11931 6686 11940
rect 6378 10908 6686 10917
rect 6378 10906 6384 10908
rect 6440 10906 6464 10908
rect 6520 10906 6544 10908
rect 6600 10906 6624 10908
rect 6680 10906 6686 10908
rect 6440 10854 6442 10906
rect 6622 10854 6624 10906
rect 6378 10852 6384 10854
rect 6440 10852 6464 10854
rect 6520 10852 6544 10854
rect 6600 10852 6624 10854
rect 6680 10852 6686 10854
rect 6378 10843 6686 10852
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6656 10674 6684 10746
rect 6644 10668 6696 10674
rect 6196 10628 6408 10656
rect 6274 10568 6330 10577
rect 6184 10532 6236 10538
rect 6274 10503 6330 10512
rect 6184 10474 6236 10480
rect 6196 10062 6224 10474
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6196 8548 6224 9862
rect 6288 9382 6316 10503
rect 6380 9926 6408 10628
rect 6644 10610 6696 10616
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6656 10146 6684 10406
rect 6748 10266 6776 12106
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6656 10130 6776 10146
rect 6644 10124 6776 10130
rect 6696 10118 6776 10124
rect 6644 10066 6696 10072
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6378 9820 6686 9829
rect 6378 9818 6384 9820
rect 6440 9818 6464 9820
rect 6520 9818 6544 9820
rect 6600 9818 6624 9820
rect 6680 9818 6686 9820
rect 6440 9766 6442 9818
rect 6622 9766 6624 9818
rect 6378 9764 6384 9766
rect 6440 9764 6464 9766
rect 6520 9764 6544 9766
rect 6600 9764 6624 9766
rect 6680 9764 6686 9766
rect 6378 9755 6686 9764
rect 6748 9722 6776 10118
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6378 8732 6686 8741
rect 6378 8730 6384 8732
rect 6440 8730 6464 8732
rect 6520 8730 6544 8732
rect 6600 8730 6624 8732
rect 6680 8730 6686 8732
rect 6440 8678 6442 8730
rect 6622 8678 6624 8730
rect 6378 8676 6384 8678
rect 6440 8676 6464 8678
rect 6520 8676 6544 8678
rect 6600 8676 6624 8678
rect 6680 8676 6686 8678
rect 6378 8667 6686 8676
rect 6840 8634 6868 13806
rect 7300 13530 7328 13874
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7392 10606 7420 12038
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7300 9654 7328 10542
rect 7392 10130 7420 10542
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7300 9042 7328 9386
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6196 8520 6408 8548
rect 6380 7886 6408 8520
rect 7300 8498 7328 8978
rect 7484 8974 7512 11222
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7380 8560 7432 8566
rect 7380 8502 7432 8508
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6748 7818 6776 8434
rect 6736 7812 6788 7818
rect 6736 7754 6788 7760
rect 6378 7644 6686 7653
rect 6378 7642 6384 7644
rect 6440 7642 6464 7644
rect 6520 7642 6544 7644
rect 6600 7642 6624 7644
rect 6680 7642 6686 7644
rect 6440 7590 6442 7642
rect 6622 7590 6624 7642
rect 6378 7588 6384 7590
rect 6440 7588 6464 7590
rect 6520 7588 6544 7590
rect 6600 7588 6624 7590
rect 6680 7588 6686 7590
rect 6378 7579 6686 7588
rect 6748 7410 6776 7754
rect 6932 7546 6960 8434
rect 7392 8242 7420 8502
rect 7484 8362 7512 8910
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7392 8214 7512 8242
rect 7010 7984 7066 7993
rect 7010 7919 7066 7928
rect 7380 7948 7432 7954
rect 7024 7818 7052 7919
rect 7380 7890 7432 7896
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 7024 7342 7052 7754
rect 7288 7472 7340 7478
rect 7392 7426 7420 7890
rect 7340 7420 7420 7426
rect 7288 7414 7420 7420
rect 7300 7398 7420 7414
rect 7392 7342 7420 7398
rect 7484 7342 7512 8214
rect 7576 8090 7604 14282
rect 7668 14006 7696 14894
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8220 14006 8248 14350
rect 7656 14000 7708 14006
rect 7656 13942 7708 13948
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8220 12646 8248 13942
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8220 12238 8248 12582
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8220 11762 8248 12174
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8312 10810 8340 12854
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7668 10062 7696 10610
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7760 9926 7788 10678
rect 8300 10532 8352 10538
rect 8300 10474 8352 10480
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7760 9586 7788 9862
rect 7932 9648 7984 9654
rect 7932 9590 7984 9596
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7760 9178 7788 9522
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7944 7886 7972 9590
rect 8128 9518 8156 10406
rect 8312 10248 8340 10474
rect 8220 10220 8340 10248
rect 8220 9586 8248 10220
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8312 9654 8340 10066
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7944 7410 7972 7822
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 6378 6556 6686 6565
rect 6378 6554 6384 6556
rect 6440 6554 6464 6556
rect 6520 6554 6544 6556
rect 6600 6554 6624 6556
rect 6680 6554 6686 6556
rect 6440 6502 6442 6554
rect 6622 6502 6624 6554
rect 6378 6500 6384 6502
rect 6440 6500 6464 6502
rect 6520 6500 6544 6502
rect 6600 6500 6624 6502
rect 6680 6500 6686 6502
rect 6378 6491 6686 6500
rect 6378 5468 6686 5477
rect 6378 5466 6384 5468
rect 6440 5466 6464 5468
rect 6520 5466 6544 5468
rect 6600 5466 6624 5468
rect 6680 5466 6686 5468
rect 6440 5414 6442 5466
rect 6622 5414 6624 5466
rect 6378 5412 6384 5414
rect 6440 5412 6464 5414
rect 6520 5412 6544 5414
rect 6600 5412 6624 5414
rect 6680 5412 6686 5414
rect 6378 5403 6686 5412
rect 6378 4380 6686 4389
rect 6378 4378 6384 4380
rect 6440 4378 6464 4380
rect 6520 4378 6544 4380
rect 6600 4378 6624 4380
rect 6680 4378 6686 4380
rect 6440 4326 6442 4378
rect 6622 4326 6624 4378
rect 6378 4324 6384 4326
rect 6440 4324 6464 4326
rect 6520 4324 6544 4326
rect 6600 4324 6624 4326
rect 6680 4324 6686 4326
rect 6378 4315 6686 4324
rect 6378 3292 6686 3301
rect 6378 3290 6384 3292
rect 6440 3290 6464 3292
rect 6520 3290 6544 3292
rect 6600 3290 6624 3292
rect 6680 3290 6686 3292
rect 6440 3238 6442 3290
rect 6622 3238 6624 3290
rect 6378 3236 6384 3238
rect 6440 3236 6464 3238
rect 6520 3236 6544 3238
rect 6600 3236 6624 3238
rect 6680 3236 6686 3238
rect 6378 3227 6686 3236
rect 6092 2576 6144 2582
rect 6092 2518 6144 2524
rect 8404 2446 8432 16390
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8496 10266 8524 10610
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8588 9722 8616 11698
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8496 8090 8524 8366
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8496 7478 8524 8026
rect 8680 8022 8708 13670
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8680 7206 8708 7958
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8772 2774 8800 16934
rect 9092 16892 9400 16901
rect 9092 16890 9098 16892
rect 9154 16890 9178 16892
rect 9234 16890 9258 16892
rect 9314 16890 9338 16892
rect 9394 16890 9400 16892
rect 9154 16838 9156 16890
rect 9336 16838 9338 16890
rect 9092 16836 9098 16838
rect 9154 16836 9178 16838
rect 9234 16836 9258 16838
rect 9314 16836 9338 16838
rect 9394 16836 9400 16838
rect 9092 16827 9400 16836
rect 9692 16658 9720 17070
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 10612 15910 10640 17546
rect 11716 17202 11744 17818
rect 11806 17436 12114 17445
rect 11806 17434 11812 17436
rect 11868 17434 11892 17436
rect 11948 17434 11972 17436
rect 12028 17434 12052 17436
rect 12108 17434 12114 17436
rect 11868 17382 11870 17434
rect 12050 17382 12052 17434
rect 11806 17380 11812 17382
rect 11868 17380 11892 17382
rect 11948 17380 11972 17382
rect 12028 17380 12052 17382
rect 12108 17380 12114 17382
rect 11806 17371 12114 17380
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11716 16658 11744 17138
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 12164 16516 12216 16522
rect 12164 16458 12216 16464
rect 11806 16348 12114 16357
rect 11806 16346 11812 16348
rect 11868 16346 11892 16348
rect 11948 16346 11972 16348
rect 12028 16346 12052 16348
rect 12108 16346 12114 16348
rect 11868 16294 11870 16346
rect 12050 16294 12052 16346
rect 11806 16292 11812 16294
rect 11868 16292 11892 16294
rect 11948 16292 11972 16294
rect 12028 16292 12052 16294
rect 12108 16292 12114 16294
rect 11806 16283 12114 16292
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 9092 15804 9400 15813
rect 9092 15802 9098 15804
rect 9154 15802 9178 15804
rect 9234 15802 9258 15804
rect 9314 15802 9338 15804
rect 9394 15802 9400 15804
rect 9154 15750 9156 15802
rect 9336 15750 9338 15802
rect 9092 15748 9098 15750
rect 9154 15748 9178 15750
rect 9234 15748 9258 15750
rect 9314 15748 9338 15750
rect 9394 15748 9400 15750
rect 9092 15739 9400 15748
rect 9692 15502 9720 15846
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8588 2746 8800 2774
rect 8588 2446 8616 2746
rect 8864 2514 8892 14758
rect 9092 14716 9400 14725
rect 9092 14714 9098 14716
rect 9154 14714 9178 14716
rect 9234 14714 9258 14716
rect 9314 14714 9338 14716
rect 9394 14714 9400 14716
rect 9154 14662 9156 14714
rect 9336 14662 9338 14714
rect 9092 14660 9098 14662
rect 9154 14660 9178 14662
rect 9234 14660 9258 14662
rect 9314 14660 9338 14662
rect 9394 14660 9400 14662
rect 9092 14651 9400 14660
rect 9600 14414 9628 15438
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9784 13870 9812 14214
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9092 13628 9400 13637
rect 9092 13626 9098 13628
rect 9154 13626 9178 13628
rect 9234 13626 9258 13628
rect 9314 13626 9338 13628
rect 9394 13626 9400 13628
rect 9154 13574 9156 13626
rect 9336 13574 9338 13626
rect 9092 13572 9098 13574
rect 9154 13572 9178 13574
rect 9234 13572 9258 13574
rect 9314 13572 9338 13574
rect 9394 13572 9400 13574
rect 9092 13563 9400 13572
rect 9784 12782 9812 13806
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9092 12540 9400 12549
rect 9092 12538 9098 12540
rect 9154 12538 9178 12540
rect 9234 12538 9258 12540
rect 9314 12538 9338 12540
rect 9394 12538 9400 12540
rect 9154 12486 9156 12538
rect 9336 12486 9338 12538
rect 9092 12484 9098 12486
rect 9154 12484 9178 12486
rect 9234 12484 9258 12486
rect 9314 12484 9338 12486
rect 9394 12484 9400 12486
rect 9092 12475 9400 12484
rect 9092 11452 9400 11461
rect 9092 11450 9098 11452
rect 9154 11450 9178 11452
rect 9234 11450 9258 11452
rect 9314 11450 9338 11452
rect 9394 11450 9400 11452
rect 9154 11398 9156 11450
rect 9336 11398 9338 11450
rect 9092 11396 9098 11398
rect 9154 11396 9178 11398
rect 9234 11396 9258 11398
rect 9314 11396 9338 11398
rect 9394 11396 9400 11398
rect 9092 11387 9400 11396
rect 9600 10674 9628 12582
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9692 10742 9720 11494
rect 9680 10736 9732 10742
rect 9678 10704 9680 10713
rect 9732 10704 9734 10713
rect 9588 10668 9640 10674
rect 9678 10639 9734 10648
rect 9588 10610 9640 10616
rect 9496 10532 9548 10538
rect 9496 10474 9548 10480
rect 9092 10364 9400 10373
rect 9092 10362 9098 10364
rect 9154 10362 9178 10364
rect 9234 10362 9258 10364
rect 9314 10362 9338 10364
rect 9394 10362 9400 10364
rect 9154 10310 9156 10362
rect 9336 10310 9338 10362
rect 9092 10308 9098 10310
rect 9154 10308 9178 10310
rect 9234 10308 9258 10310
rect 9314 10308 9338 10310
rect 9394 10308 9400 10310
rect 9092 10299 9400 10308
rect 9508 10010 9536 10474
rect 9600 10062 9628 10610
rect 9416 9982 9536 10010
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9416 9432 9444 9982
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9508 9722 9536 9862
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9600 9586 9628 9998
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9416 9404 9536 9432
rect 9092 9276 9400 9285
rect 9092 9274 9098 9276
rect 9154 9274 9178 9276
rect 9234 9274 9258 9276
rect 9314 9274 9338 9276
rect 9394 9274 9400 9276
rect 9154 9222 9156 9274
rect 9336 9222 9338 9274
rect 9092 9220 9098 9222
rect 9154 9220 9178 9222
rect 9234 9220 9258 9222
rect 9314 9220 9338 9222
rect 9394 9220 9400 9222
rect 9092 9211 9400 9220
rect 9508 8548 9536 9404
rect 9416 8520 9536 8548
rect 9416 8430 9444 8520
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9416 8294 9444 8366
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 8956 7970 8984 8230
rect 9092 8188 9400 8197
rect 9092 8186 9098 8188
rect 9154 8186 9178 8188
rect 9234 8186 9258 8188
rect 9314 8186 9338 8188
rect 9394 8186 9400 8188
rect 9154 8134 9156 8186
rect 9336 8134 9338 8186
rect 9092 8132 9098 8134
rect 9154 8132 9178 8134
rect 9234 8132 9258 8134
rect 9314 8132 9338 8134
rect 9394 8132 9400 8134
rect 9092 8123 9400 8132
rect 8956 7942 9260 7970
rect 9232 7206 9260 7942
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9416 7546 9444 7822
rect 9508 7818 9536 8298
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9600 7750 9628 8434
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9600 7274 9628 7686
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9092 7100 9400 7109
rect 9092 7098 9098 7100
rect 9154 7098 9178 7100
rect 9234 7098 9258 7100
rect 9314 7098 9338 7100
rect 9394 7098 9400 7100
rect 9154 7046 9156 7098
rect 9336 7046 9338 7098
rect 9092 7044 9098 7046
rect 9154 7044 9178 7046
rect 9234 7044 9258 7046
rect 9314 7044 9338 7046
rect 9394 7044 9400 7046
rect 9092 7035 9400 7044
rect 9784 7002 9812 8366
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9968 8090 9996 8230
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10060 7546 10088 13874
rect 10612 13326 10640 15846
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10336 10266 10364 12174
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10520 9926 10548 12038
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10612 9450 10640 9998
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10704 8430 10732 14214
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10796 9722 10824 9930
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10612 7546 10640 7686
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10704 7410 10732 7686
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9092 6012 9400 6021
rect 9092 6010 9098 6012
rect 9154 6010 9178 6012
rect 9234 6010 9258 6012
rect 9314 6010 9338 6012
rect 9394 6010 9400 6012
rect 9154 5958 9156 6010
rect 9336 5958 9338 6010
rect 9092 5956 9098 5958
rect 9154 5956 9178 5958
rect 9234 5956 9258 5958
rect 9314 5956 9338 5958
rect 9394 5956 9400 5958
rect 9092 5947 9400 5956
rect 9092 4924 9400 4933
rect 9092 4922 9098 4924
rect 9154 4922 9178 4924
rect 9234 4922 9258 4924
rect 9314 4922 9338 4924
rect 9394 4922 9400 4924
rect 9154 4870 9156 4922
rect 9336 4870 9338 4922
rect 9092 4868 9098 4870
rect 9154 4868 9178 4870
rect 9234 4868 9258 4870
rect 9314 4868 9338 4870
rect 9394 4868 9400 4870
rect 9092 4859 9400 4868
rect 9092 3836 9400 3845
rect 9092 3834 9098 3836
rect 9154 3834 9178 3836
rect 9234 3834 9258 3836
rect 9314 3834 9338 3836
rect 9394 3834 9400 3836
rect 9154 3782 9156 3834
rect 9336 3782 9338 3834
rect 9092 3780 9098 3782
rect 9154 3780 9178 3782
rect 9234 3780 9258 3782
rect 9314 3780 9338 3782
rect 9394 3780 9400 3782
rect 9092 3771 9400 3780
rect 9092 2748 9400 2757
rect 9092 2746 9098 2748
rect 9154 2746 9178 2748
rect 9234 2746 9258 2748
rect 9314 2746 9338 2748
rect 9394 2746 9400 2748
rect 9154 2694 9156 2746
rect 9336 2694 9338 2746
rect 9092 2692 9098 2694
rect 9154 2692 9178 2694
rect 9234 2692 9258 2694
rect 9314 2692 9338 2694
rect 9394 2692 9400 2694
rect 9092 2683 9400 2692
rect 10888 2650 10916 15302
rect 11806 15260 12114 15269
rect 11806 15258 11812 15260
rect 11868 15258 11892 15260
rect 11948 15258 11972 15260
rect 12028 15258 12052 15260
rect 12108 15258 12114 15260
rect 11868 15206 11870 15258
rect 12050 15206 12052 15258
rect 11806 15204 11812 15206
rect 11868 15204 11892 15206
rect 11948 15204 11972 15206
rect 12028 15204 12052 15206
rect 12108 15204 12114 15206
rect 11806 15195 12114 15204
rect 12176 15094 12204 16458
rect 12164 15088 12216 15094
rect 12164 15030 12216 15036
rect 12268 14618 12296 18158
rect 14520 17980 14828 17989
rect 14520 17978 14526 17980
rect 14582 17978 14606 17980
rect 14662 17978 14686 17980
rect 14742 17978 14766 17980
rect 14822 17978 14828 17980
rect 14582 17926 14584 17978
rect 14764 17926 14766 17978
rect 14520 17924 14526 17926
rect 14582 17924 14606 17926
rect 14662 17924 14686 17926
rect 14742 17924 14766 17926
rect 14822 17924 14828 17926
rect 14520 17915 14828 17924
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 12912 17202 12940 17478
rect 15212 17270 15240 17614
rect 15200 17264 15252 17270
rect 15200 17206 15252 17212
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 14924 17060 14976 17066
rect 14924 17002 14976 17008
rect 14520 16892 14828 16901
rect 14520 16890 14526 16892
rect 14582 16890 14606 16892
rect 14662 16890 14686 16892
rect 14742 16890 14766 16892
rect 14822 16890 14828 16892
rect 14582 16838 14584 16890
rect 14764 16838 14766 16890
rect 14520 16836 14526 16838
rect 14582 16836 14606 16838
rect 14662 16836 14686 16838
rect 14742 16836 14766 16838
rect 14822 16836 14828 16838
rect 14520 16827 14828 16836
rect 14936 16522 14964 17002
rect 14924 16516 14976 16522
rect 14924 16458 14976 16464
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12360 15502 12388 15982
rect 14520 15804 14828 15813
rect 14520 15802 14526 15804
rect 14582 15802 14606 15804
rect 14662 15802 14686 15804
rect 14742 15802 14766 15804
rect 14822 15802 14828 15804
rect 14582 15750 14584 15802
rect 14764 15750 14766 15802
rect 14520 15748 14526 15750
rect 14582 15748 14606 15750
rect 14662 15748 14686 15750
rect 14742 15748 14766 15750
rect 14822 15748 14828 15750
rect 14520 15739 14828 15748
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12360 14958 12388 15438
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12360 14414 12388 14894
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 11072 14074 11100 14350
rect 11806 14172 12114 14181
rect 11806 14170 11812 14172
rect 11868 14170 11892 14172
rect 11948 14170 11972 14172
rect 12028 14170 12052 14172
rect 12108 14170 12114 14172
rect 11868 14118 11870 14170
rect 12050 14118 12052 14170
rect 11806 14116 11812 14118
rect 11868 14116 11892 14118
rect 11948 14116 11972 14118
rect 12028 14116 12052 14118
rect 12108 14116 12114 14118
rect 11806 14107 12114 14116
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 12360 13870 12388 14350
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11072 12306 11100 12582
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10980 9586 11008 9862
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 11164 8566 11192 13670
rect 12360 13258 12388 13806
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 11806 13084 12114 13093
rect 11806 13082 11812 13084
rect 11868 13082 11892 13084
rect 11948 13082 11972 13084
rect 12028 13082 12052 13084
rect 12108 13082 12114 13084
rect 11868 13030 11870 13082
rect 12050 13030 12052 13082
rect 11806 13028 11812 13030
rect 11868 13028 11892 13030
rect 11948 13028 11972 13030
rect 12028 13028 12052 13030
rect 12108 13028 12114 13030
rect 11806 13019 12114 13028
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11256 10266 11284 12106
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10980 7970 11008 8230
rect 10980 7942 11100 7970
rect 11072 7886 11100 7942
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10980 6934 11008 7822
rect 11164 7410 11192 8502
rect 11440 8498 11468 9522
rect 11624 8634 11652 12786
rect 12360 12782 12388 13194
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12360 12238 12388 12718
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 11806 11996 12114 12005
rect 11806 11994 11812 11996
rect 11868 11994 11892 11996
rect 11948 11994 11972 11996
rect 12028 11994 12052 11996
rect 12108 11994 12114 11996
rect 11868 11942 11870 11994
rect 12050 11942 12052 11994
rect 11806 11940 11812 11942
rect 11868 11940 11892 11942
rect 11948 11940 11972 11942
rect 12028 11940 12052 11942
rect 12108 11940 12114 11942
rect 11806 11931 12114 11940
rect 12360 11762 12388 12174
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 11806 10908 12114 10917
rect 11806 10906 11812 10908
rect 11868 10906 11892 10908
rect 11948 10906 11972 10908
rect 12028 10906 12052 10908
rect 12108 10906 12114 10908
rect 11868 10854 11870 10906
rect 12050 10854 12052 10906
rect 11806 10852 11812 10854
rect 11868 10852 11892 10854
rect 11948 10852 11972 10854
rect 12028 10852 12052 10854
rect 12108 10852 12114 10854
rect 11806 10843 12114 10852
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 13096 10266 13124 10610
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11716 9450 11744 9998
rect 11806 9820 12114 9829
rect 11806 9818 11812 9820
rect 11868 9818 11892 9820
rect 11948 9818 11972 9820
rect 12028 9818 12052 9820
rect 12108 9818 12114 9820
rect 11868 9766 11870 9818
rect 12050 9766 12052 9818
rect 11806 9764 11812 9766
rect 11868 9764 11892 9766
rect 11948 9764 11972 9766
rect 12028 9764 12052 9766
rect 12108 9764 12114 9766
rect 11806 9755 12114 9764
rect 12268 9518 12296 10202
rect 12360 9994 12388 10202
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 12440 9988 12492 9994
rect 12440 9930 12492 9936
rect 12360 9586 12388 9930
rect 12452 9722 12480 9930
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 11806 8732 12114 8741
rect 11806 8730 11812 8732
rect 11868 8730 11892 8732
rect 11948 8730 11972 8732
rect 12028 8730 12052 8732
rect 12108 8730 12114 8732
rect 11868 8678 11870 8730
rect 12050 8678 12052 8730
rect 11806 8676 11812 8678
rect 11868 8676 11892 8678
rect 11948 8676 11972 8678
rect 12028 8676 12052 8678
rect 12108 8676 12114 8678
rect 11806 8667 12114 8676
rect 12176 8634 12204 8842
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 12176 8022 12204 8570
rect 12268 8362 12296 8774
rect 12256 8356 12308 8362
rect 12256 8298 12308 8304
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 11806 7644 12114 7653
rect 11806 7642 11812 7644
rect 11868 7642 11892 7644
rect 11948 7642 11972 7644
rect 12028 7642 12052 7644
rect 12108 7642 12114 7644
rect 11868 7590 11870 7642
rect 12050 7590 12052 7642
rect 11806 7588 11812 7590
rect 11868 7588 11892 7590
rect 11948 7588 11972 7590
rect 12028 7588 12052 7590
rect 12108 7588 12114 7590
rect 11806 7579 12114 7588
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 12176 7206 12204 7958
rect 12268 7342 12296 8298
rect 12544 7954 12572 9386
rect 13188 9178 13216 11698
rect 13280 9586 13308 12582
rect 13372 10606 13400 14554
rect 13648 13938 13676 14894
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 13648 12434 13676 13874
rect 13556 12406 13676 12434
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13372 9874 13400 10066
rect 13464 10062 13492 10610
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13556 9874 13584 12406
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13372 9846 13584 9874
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13372 9450 13400 9846
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13372 9042 13400 9114
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12636 8566 12664 8910
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 13372 8430 13400 8978
rect 13464 8906 13492 9318
rect 13452 8900 13504 8906
rect 13452 8842 13504 8848
rect 13648 8634 13676 12038
rect 13636 8628 13688 8634
rect 13464 8588 13636 8616
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13464 8090 13492 8588
rect 13636 8570 13688 8576
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 12544 7750 12572 7890
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12360 7478 12388 7686
rect 12348 7472 12400 7478
rect 12348 7414 12400 7420
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 13464 7206 13492 7890
rect 13740 7460 13768 14962
rect 14520 14716 14828 14725
rect 14520 14714 14526 14716
rect 14582 14714 14606 14716
rect 14662 14714 14686 14716
rect 14742 14714 14766 14716
rect 14822 14714 14828 14716
rect 14582 14662 14584 14714
rect 14764 14662 14766 14714
rect 14520 14660 14526 14662
rect 14582 14660 14606 14662
rect 14662 14660 14686 14662
rect 14742 14660 14766 14662
rect 14822 14660 14828 14662
rect 14520 14651 14828 14660
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 13924 13802 13952 13942
rect 14660 13938 14688 14282
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 13912 13796 13964 13802
rect 13912 13738 13964 13744
rect 14520 13628 14828 13637
rect 14520 13626 14526 13628
rect 14582 13626 14606 13628
rect 14662 13626 14686 13628
rect 14742 13626 14766 13628
rect 14822 13626 14828 13628
rect 14582 13574 14584 13626
rect 14764 13574 14766 13626
rect 14520 13572 14526 13574
rect 14582 13572 14606 13574
rect 14662 13572 14686 13574
rect 14742 13572 14766 13574
rect 14822 13572 14828 13574
rect 14520 13563 14828 13572
rect 14520 12540 14828 12549
rect 14520 12538 14526 12540
rect 14582 12538 14606 12540
rect 14662 12538 14686 12540
rect 14742 12538 14766 12540
rect 14822 12538 14828 12540
rect 14582 12486 14584 12538
rect 14764 12486 14766 12538
rect 14520 12484 14526 12486
rect 14582 12484 14606 12486
rect 14662 12484 14686 12486
rect 14742 12484 14766 12486
rect 14822 12484 14828 12486
rect 14520 12475 14828 12484
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 13924 10810 13952 12106
rect 14520 11452 14828 11461
rect 14520 11450 14526 11452
rect 14582 11450 14606 11452
rect 14662 11450 14686 11452
rect 14742 11450 14766 11452
rect 14822 11450 14828 11452
rect 14582 11398 14584 11450
rect 14764 11398 14766 11450
rect 14520 11396 14526 11398
rect 14582 11396 14606 11398
rect 14662 11396 14686 11398
rect 14742 11396 14766 11398
rect 14822 11396 14828 11398
rect 14520 11387 14828 11396
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 14924 10532 14976 10538
rect 14924 10474 14976 10480
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13832 10266 13860 10406
rect 14520 10364 14828 10373
rect 14520 10362 14526 10364
rect 14582 10362 14606 10364
rect 14662 10362 14686 10364
rect 14742 10362 14766 10364
rect 14822 10362 14828 10364
rect 14582 10310 14584 10362
rect 14764 10310 14766 10362
rect 14520 10308 14526 10310
rect 14582 10308 14606 10310
rect 14662 10308 14686 10310
rect 14742 10308 14766 10310
rect 14822 10308 14828 10310
rect 14520 10299 14828 10308
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 14936 10130 14964 10474
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 14844 9586 14872 9998
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 14016 8362 14044 9522
rect 14520 9276 14828 9285
rect 14520 9274 14526 9276
rect 14582 9274 14606 9276
rect 14662 9274 14686 9276
rect 14742 9274 14766 9276
rect 14822 9274 14828 9276
rect 14582 9222 14584 9274
rect 14764 9222 14766 9274
rect 14520 9220 14526 9222
rect 14582 9220 14606 9222
rect 14662 9220 14686 9222
rect 14742 9220 14766 9222
rect 14822 9220 14828 9222
rect 14520 9211 14828 9220
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13924 7886 13952 8230
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13912 7472 13964 7478
rect 13740 7432 13912 7460
rect 13912 7414 13964 7420
rect 14016 7342 14044 8298
rect 14384 7818 14412 8434
rect 14520 8188 14828 8197
rect 14520 8186 14526 8188
rect 14582 8186 14606 8188
rect 14662 8186 14686 8188
rect 14742 8186 14766 8188
rect 14822 8186 14828 8188
rect 14582 8134 14584 8186
rect 14764 8134 14766 8186
rect 14520 8132 14526 8134
rect 14582 8132 14606 8134
rect 14662 8132 14686 8134
rect 14742 8132 14766 8134
rect 14822 8132 14828 8134
rect 14520 8123 14828 8132
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 14292 7410 14320 7754
rect 14936 7750 14964 8434
rect 15028 8294 15056 16390
rect 15396 15502 15424 20402
rect 15488 19310 15516 20878
rect 15948 20466 15976 21286
rect 16028 20868 16080 20874
rect 16028 20810 16080 20816
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 16040 20058 16068 20810
rect 16132 20262 16160 21422
rect 16408 21146 16436 21490
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 16302 21040 16358 21049
rect 16302 20975 16358 20984
rect 16316 20942 16344 20975
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 16132 19514 16160 20198
rect 16408 19922 16436 21082
rect 16500 20942 16528 21558
rect 19708 21480 19760 21486
rect 19708 21422 19760 21428
rect 17132 21412 17184 21418
rect 17132 21354 17184 21360
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16500 20806 16528 20878
rect 16488 20800 16540 20806
rect 16488 20742 16540 20748
rect 16500 20466 16528 20742
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 17052 19990 17080 20402
rect 17040 19984 17092 19990
rect 17040 19926 17092 19932
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16408 19786 16436 19858
rect 16396 19780 16448 19786
rect 16396 19722 16448 19728
rect 16120 19508 16172 19514
rect 16120 19450 16172 19456
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15488 17882 15516 18226
rect 15672 18086 15700 18702
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15764 18290 15792 18566
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15672 17678 15700 18022
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15764 17542 15792 18226
rect 16040 18222 16068 19246
rect 16408 19174 16436 19722
rect 17052 19446 17080 19926
rect 17040 19440 17092 19446
rect 17040 19382 17092 19388
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 16040 16590 16068 18158
rect 16212 18148 16264 18154
rect 16212 18090 16264 18096
rect 16224 17678 16252 18090
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16408 17610 16436 19110
rect 16500 18766 16528 19246
rect 16592 18970 16620 19314
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 17052 18698 17080 19382
rect 17144 19310 17172 21354
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 17236 20874 17264 21082
rect 17316 21072 17368 21078
rect 17314 21040 17316 21049
rect 17368 21040 17370 21049
rect 17314 20975 17370 20984
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 17224 20868 17276 20874
rect 17224 20810 17276 20816
rect 17234 20700 17542 20709
rect 17234 20698 17240 20700
rect 17296 20698 17320 20700
rect 17376 20698 17400 20700
rect 17456 20698 17480 20700
rect 17536 20698 17542 20700
rect 17296 20646 17298 20698
rect 17478 20646 17480 20698
rect 17234 20644 17240 20646
rect 17296 20644 17320 20646
rect 17376 20644 17400 20646
rect 17456 20644 17480 20646
rect 17536 20644 17542 20646
rect 17234 20635 17542 20644
rect 17972 20602 18000 20946
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 18248 20602 18276 20878
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18788 20800 18840 20806
rect 18788 20742 18840 20748
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 18236 20596 18288 20602
rect 18236 20538 18288 20544
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17236 19854 17264 20402
rect 18708 20330 18736 20742
rect 18696 20324 18748 20330
rect 18696 20266 18748 20272
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 17234 19612 17542 19621
rect 17234 19610 17240 19612
rect 17296 19610 17320 19612
rect 17376 19610 17400 19612
rect 17456 19610 17480 19612
rect 17536 19610 17542 19612
rect 17296 19558 17298 19610
rect 17478 19558 17480 19610
rect 17234 19556 17240 19558
rect 17296 19556 17320 19558
rect 17376 19556 17400 19558
rect 17456 19556 17480 19558
rect 17536 19556 17542 19558
rect 17234 19547 17542 19556
rect 18708 19446 18736 20266
rect 18696 19440 18748 19446
rect 18696 19382 18748 19388
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 17040 18692 17092 18698
rect 17040 18634 17092 18640
rect 17144 18630 17172 19246
rect 18616 18766 18644 19314
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18708 18766 18736 19110
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 17234 18524 17542 18533
rect 17234 18522 17240 18524
rect 17296 18522 17320 18524
rect 17376 18522 17400 18524
rect 17456 18522 17480 18524
rect 17536 18522 17542 18524
rect 17296 18470 17298 18522
rect 17478 18470 17480 18522
rect 17234 18468 17240 18470
rect 17296 18468 17320 18470
rect 17376 18468 17400 18470
rect 17456 18468 17480 18470
rect 17536 18468 17542 18470
rect 17234 18459 17542 18468
rect 18524 18358 18552 18566
rect 18512 18352 18564 18358
rect 18512 18294 18564 18300
rect 18800 18222 18828 20742
rect 19444 20466 19472 21286
rect 19720 20942 19748 21422
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 19812 21026 19840 21286
rect 19948 21244 20256 21253
rect 19948 21242 19954 21244
rect 20010 21242 20034 21244
rect 20090 21242 20114 21244
rect 20170 21242 20194 21244
rect 20250 21242 20256 21244
rect 20010 21190 20012 21242
rect 20192 21190 20194 21242
rect 19948 21188 19954 21190
rect 20010 21188 20034 21190
rect 20090 21188 20114 21190
rect 20170 21188 20194 21190
rect 20250 21188 20256 21190
rect 19948 21179 20256 21188
rect 19812 20998 19932 21026
rect 19904 20942 19932 20998
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18984 19378 19012 20334
rect 19948 20156 20256 20165
rect 19948 20154 19954 20156
rect 20010 20154 20034 20156
rect 20090 20154 20114 20156
rect 20170 20154 20194 20156
rect 20250 20154 20256 20156
rect 20010 20102 20012 20154
rect 20192 20102 20194 20154
rect 19948 20100 19954 20102
rect 20010 20100 20034 20102
rect 20090 20100 20114 20102
rect 20170 20100 20194 20102
rect 20250 20100 20256 20102
rect 19948 20091 20256 20100
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 18788 18216 18840 18222
rect 18788 18158 18840 18164
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 16396 17604 16448 17610
rect 16396 17546 16448 17552
rect 16948 17536 17000 17542
rect 16948 17478 17000 17484
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16500 16794 16528 17138
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 16040 15502 16068 16526
rect 16132 15978 16160 16594
rect 16960 16114 16988 17478
rect 17234 17436 17542 17445
rect 17234 17434 17240 17436
rect 17296 17434 17320 17436
rect 17376 17434 17400 17436
rect 17456 17434 17480 17436
rect 17536 17434 17542 17436
rect 17296 17382 17298 17434
rect 17478 17382 17480 17434
rect 17234 17380 17240 17382
rect 17296 17380 17320 17382
rect 17376 17380 17400 17382
rect 17456 17380 17480 17382
rect 17536 17380 17542 17382
rect 17234 17371 17542 17380
rect 18248 17202 18276 18022
rect 18800 17610 18828 18158
rect 18788 17604 18840 17610
rect 18788 17546 18840 17552
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19260 17338 19288 17546
rect 19352 17490 19380 19246
rect 19616 19168 19668 19174
rect 19616 19110 19668 19116
rect 19628 18766 19656 19110
rect 19948 19068 20256 19077
rect 19948 19066 19954 19068
rect 20010 19066 20034 19068
rect 20090 19066 20114 19068
rect 20170 19066 20194 19068
rect 20250 19066 20256 19068
rect 20010 19014 20012 19066
rect 20192 19014 20194 19066
rect 19948 19012 19954 19014
rect 20010 19012 20034 19014
rect 20090 19012 20114 19014
rect 20170 19012 20194 19014
rect 20250 19012 20256 19014
rect 19948 19003 20256 19012
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19616 18624 19668 18630
rect 19616 18566 19668 18572
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19444 17678 19472 18294
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19352 17462 19472 17490
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 17684 17128 17736 17134
rect 17684 17070 17736 17076
rect 17696 16658 17724 17070
rect 18236 17060 18288 17066
rect 18236 17002 18288 17008
rect 17684 16652 17736 16658
rect 17684 16594 17736 16600
rect 18248 16590 18276 17002
rect 18708 16794 18736 17138
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 17224 16584 17276 16590
rect 17144 16532 17224 16538
rect 17144 16526 17276 16532
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 17144 16510 17264 16526
rect 17144 16114 17172 16510
rect 17234 16348 17542 16357
rect 17234 16346 17240 16348
rect 17296 16346 17320 16348
rect 17376 16346 17400 16348
rect 17456 16346 17480 16348
rect 17536 16346 17542 16348
rect 17296 16294 17298 16346
rect 17478 16294 17480 16346
rect 17234 16292 17240 16294
rect 17296 16292 17320 16294
rect 17376 16292 17400 16294
rect 17456 16292 17480 16294
rect 17536 16292 17542 16294
rect 17234 16283 17542 16292
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 17132 16108 17184 16114
rect 17132 16050 17184 16056
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 16120 15972 16172 15978
rect 16120 15914 16172 15920
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 15120 15162 15148 15370
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15108 15156 15160 15162
rect 15108 15098 15160 15104
rect 15580 15026 15608 15302
rect 16132 15026 16160 15914
rect 16776 15706 16804 15982
rect 18340 15978 18368 16526
rect 18524 16182 18552 16526
rect 18512 16176 18564 16182
rect 18512 16118 18564 16124
rect 18328 15972 18380 15978
rect 18328 15914 18380 15920
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 16488 15428 16540 15434
rect 16488 15370 16540 15376
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15212 12850 15240 13874
rect 15396 13870 15424 14826
rect 15580 14074 15608 14962
rect 16500 14958 16528 15370
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16500 14618 16528 14894
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 15752 14340 15804 14346
rect 15752 14282 15804 14288
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15212 12434 15240 12786
rect 15396 12782 15424 13806
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15120 12406 15240 12434
rect 15292 12436 15344 12442
rect 15120 9926 15148 12406
rect 15292 12378 15344 12384
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15212 10062 15240 11630
rect 15304 10674 15332 12378
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15396 10198 15424 12718
rect 15672 12306 15700 14214
rect 15764 14090 15792 14282
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 15764 14062 15884 14090
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15672 11762 15700 12242
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15488 11098 15516 11562
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15580 11286 15608 11494
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15672 11218 15700 11698
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15488 11070 15608 11098
rect 15384 10192 15436 10198
rect 15384 10134 15436 10140
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15212 8566 15240 9590
rect 15304 8974 15332 9930
rect 15488 9518 15516 9998
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15200 8560 15252 8566
rect 15200 8502 15252 8508
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 15028 7970 15056 8230
rect 15028 7942 15148 7970
rect 15120 7818 15148 7942
rect 15016 7812 15068 7818
rect 15016 7754 15068 7760
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 15028 7274 15056 7754
rect 15016 7268 15068 7274
rect 15016 7210 15068 7216
rect 15304 7206 15332 8910
rect 15488 8430 15516 9454
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15580 8090 15608 11070
rect 15672 10606 15700 11154
rect 15764 10674 15792 13942
rect 15856 13938 15884 14062
rect 16040 13938 16068 14214
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 15856 12374 15884 13874
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16224 13190 16252 13806
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16224 12850 16252 13126
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 15844 12368 15896 12374
rect 15844 12310 15896 12316
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15672 10130 15700 10406
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15764 9178 15792 9998
rect 15856 9994 15884 12310
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16028 10124 16080 10130
rect 16028 10066 16080 10072
rect 15844 9988 15896 9994
rect 15844 9930 15896 9936
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 15948 9586 15976 9862
rect 16040 9654 16068 10066
rect 16132 9722 16160 12174
rect 16500 11626 16528 13874
rect 16684 13870 16712 14418
rect 16776 14414 16804 14962
rect 16868 14822 16896 15846
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 17144 15162 17172 15642
rect 18340 15502 18368 15914
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17234 15260 17542 15269
rect 17234 15258 17240 15260
rect 17296 15258 17320 15260
rect 17376 15258 17400 15260
rect 17456 15258 17480 15260
rect 17536 15258 17542 15260
rect 17296 15206 17298 15258
rect 17478 15206 17480 15258
rect 17234 15204 17240 15206
rect 17296 15204 17320 15206
rect 17376 15204 17400 15206
rect 17456 15204 17480 15206
rect 17536 15204 17542 15206
rect 17234 15195 17542 15204
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16776 13394 16804 14350
rect 16868 14346 16896 14758
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 17052 14414 17080 14554
rect 17604 14550 17632 15302
rect 18524 15026 18552 16118
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 17592 14544 17644 14550
rect 17592 14486 17644 14492
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 16868 13258 16896 14282
rect 17604 14278 17632 14486
rect 17972 14414 18000 14962
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17234 14172 17542 14181
rect 17234 14170 17240 14172
rect 17296 14170 17320 14172
rect 17376 14170 17400 14172
rect 17456 14170 17480 14172
rect 17536 14170 17542 14172
rect 17296 14118 17298 14170
rect 17478 14118 17480 14170
rect 17234 14116 17240 14118
rect 17296 14116 17320 14118
rect 17376 14116 17400 14118
rect 17456 14116 17480 14118
rect 17536 14116 17542 14118
rect 17234 14107 17542 14116
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 16960 13326 16988 13806
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16856 13252 16908 13258
rect 16856 13194 16908 13200
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16592 12646 16620 13126
rect 16868 12832 16896 13194
rect 17234 13084 17542 13093
rect 17234 13082 17240 13084
rect 17296 13082 17320 13084
rect 17376 13082 17400 13084
rect 17456 13082 17480 13084
rect 17536 13082 17542 13084
rect 17296 13030 17298 13082
rect 17478 13030 17480 13082
rect 17234 13028 17240 13030
rect 17296 13028 17320 13030
rect 17376 13028 17400 13030
rect 17456 13028 17480 13030
rect 17536 13028 17542 13030
rect 17234 13019 17542 13028
rect 16868 12804 16988 12832
rect 16856 12708 16908 12714
rect 16856 12650 16908 12656
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16592 12306 16620 12582
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16212 10532 16264 10538
rect 16212 10474 16264 10480
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 16132 9178 16160 9658
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 16132 8022 16160 9114
rect 16224 8974 16252 10474
rect 16316 9654 16344 11222
rect 16592 10674 16620 12242
rect 16868 11898 16896 12650
rect 16960 12374 16988 12804
rect 16948 12368 17000 12374
rect 16948 12310 17000 12316
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16592 9994 16620 10610
rect 16960 10470 16988 12310
rect 17234 11996 17542 12005
rect 17234 11994 17240 11996
rect 17296 11994 17320 11996
rect 17376 11994 17400 11996
rect 17456 11994 17480 11996
rect 17536 11994 17542 11996
rect 17296 11942 17298 11994
rect 17478 11942 17480 11994
rect 17234 11940 17240 11942
rect 17296 11940 17320 11942
rect 17376 11940 17400 11942
rect 17456 11940 17480 11942
rect 17536 11940 17542 11942
rect 17234 11931 17542 11940
rect 17604 11762 17632 14214
rect 18064 13326 18092 14962
rect 18616 14618 18644 15982
rect 18788 15360 18840 15366
rect 18788 15302 18840 15308
rect 18800 14890 18828 15302
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18616 14414 18644 14554
rect 18800 14550 18828 14826
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18708 13938 18736 14214
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 17052 11082 17080 11698
rect 17880 11150 17908 12242
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 17052 10130 17080 11018
rect 17234 10908 17542 10917
rect 17234 10906 17240 10908
rect 17296 10906 17320 10908
rect 17376 10906 17400 10908
rect 17456 10906 17480 10908
rect 17536 10906 17542 10908
rect 17296 10854 17298 10906
rect 17478 10854 17480 10906
rect 17234 10852 17240 10854
rect 17296 10852 17320 10854
rect 17376 10852 17400 10854
rect 17456 10852 17480 10854
rect 17536 10852 17542 10854
rect 17234 10843 17542 10852
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 18064 10062 18092 13262
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 16580 9988 16632 9994
rect 16580 9930 16632 9936
rect 17960 9988 18012 9994
rect 17960 9930 18012 9936
rect 17234 9820 17542 9829
rect 17234 9818 17240 9820
rect 17296 9818 17320 9820
rect 17376 9818 17400 9820
rect 17456 9818 17480 9820
rect 17536 9818 17542 9820
rect 17296 9766 17298 9818
rect 17478 9766 17480 9818
rect 17234 9764 17240 9766
rect 17296 9764 17320 9766
rect 17376 9764 17400 9766
rect 17456 9764 17480 9766
rect 17536 9764 17542 9766
rect 17234 9755 17542 9764
rect 17972 9654 18000 9930
rect 16304 9648 16356 9654
rect 16304 9590 16356 9596
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 16316 8090 16344 9590
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16408 8906 16436 9454
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16120 8016 16172 8022
rect 16120 7958 16172 7964
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 15844 7472 15896 7478
rect 15844 7414 15896 7420
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 14520 7100 14828 7109
rect 14520 7098 14526 7100
rect 14582 7098 14606 7100
rect 14662 7098 14686 7100
rect 14742 7098 14766 7100
rect 14822 7098 14828 7100
rect 14582 7046 14584 7098
rect 14764 7046 14766 7098
rect 14520 7044 14526 7046
rect 14582 7044 14606 7046
rect 14662 7044 14686 7046
rect 14742 7044 14766 7046
rect 14822 7044 14828 7046
rect 14520 7035 14828 7044
rect 15856 7002 15884 7414
rect 16040 7206 16068 7686
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 16132 6798 16160 7822
rect 16408 7478 16436 8842
rect 17234 8732 17542 8741
rect 17234 8730 17240 8732
rect 17296 8730 17320 8732
rect 17376 8730 17400 8732
rect 17456 8730 17480 8732
rect 17536 8730 17542 8732
rect 17296 8678 17298 8730
rect 17478 8678 17480 8730
rect 17234 8676 17240 8678
rect 17296 8676 17320 8678
rect 17376 8676 17400 8678
rect 17456 8676 17480 8678
rect 17536 8676 17542 8678
rect 17234 8667 17542 8676
rect 17972 8634 18000 9590
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 16488 8560 16540 8566
rect 16540 8508 16620 8514
rect 16488 8502 16620 8508
rect 16500 8486 16620 8502
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16500 7886 16528 8366
rect 16592 8362 16620 8486
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16488 7880 16540 7886
rect 16488 7822 16540 7828
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 16500 6798 16528 7822
rect 16592 7818 16620 8298
rect 17040 8016 17092 8022
rect 16946 7984 17002 7993
rect 17040 7958 17092 7964
rect 16946 7919 17002 7928
rect 16960 7886 16988 7919
rect 17052 7886 17080 7958
rect 18156 7954 18184 12582
rect 18328 12300 18380 12306
rect 18328 12242 18380 12248
rect 18236 12164 18288 12170
rect 18236 12106 18288 12112
rect 18248 11762 18276 12106
rect 18340 11898 18368 12242
rect 18524 12102 18552 12650
rect 18616 12170 18644 12718
rect 18708 12646 18736 13126
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18340 11150 18368 11834
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18234 10704 18290 10713
rect 18616 10674 18644 11154
rect 18234 10639 18236 10648
rect 18288 10639 18290 10648
rect 18604 10668 18656 10674
rect 18236 10610 18288 10616
rect 18604 10610 18656 10616
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18420 10192 18472 10198
rect 18420 10134 18472 10140
rect 18432 10033 18460 10134
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18418 10024 18474 10033
rect 18418 9959 18474 9968
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18340 8566 18368 8910
rect 18328 8560 18380 8566
rect 18328 8502 18380 8508
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 16580 7812 16632 7818
rect 16580 7754 16632 7760
rect 16592 7410 16620 7754
rect 16960 7478 16988 7822
rect 16948 7472 17000 7478
rect 16948 7414 17000 7420
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 17052 7342 17080 7822
rect 17234 7644 17542 7653
rect 17234 7642 17240 7644
rect 17296 7642 17320 7644
rect 17376 7642 17400 7644
rect 17456 7642 17480 7644
rect 17536 7642 17542 7644
rect 17296 7590 17298 7642
rect 17478 7590 17480 7642
rect 17234 7588 17240 7590
rect 17296 7588 17320 7590
rect 17376 7588 17400 7590
rect 17456 7588 17480 7590
rect 17536 7588 17542 7590
rect 17234 7579 17542 7588
rect 18064 7546 18092 7822
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 18248 6934 18276 8434
rect 18340 8022 18368 8502
rect 18524 8090 18552 10066
rect 18708 9586 18736 10610
rect 18800 9722 18828 14350
rect 18892 13870 18920 15098
rect 19260 14958 19288 16594
rect 19352 16114 19380 17206
rect 19444 16590 19472 17462
rect 19628 17202 19656 18566
rect 19948 17980 20256 17989
rect 19948 17978 19954 17980
rect 20010 17978 20034 17980
rect 20090 17978 20114 17980
rect 20170 17978 20194 17980
rect 20250 17978 20256 17980
rect 20010 17926 20012 17978
rect 20192 17926 20194 17978
rect 19948 17924 19954 17926
rect 20010 17924 20034 17926
rect 20090 17924 20114 17926
rect 20170 17924 20194 17926
rect 20250 17924 20256 17926
rect 19948 17915 20256 17924
rect 19800 17604 19852 17610
rect 19800 17546 19852 17552
rect 19812 17270 19840 17546
rect 19800 17264 19852 17270
rect 19800 17206 19852 17212
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19536 16114 19564 17138
rect 19628 16658 19656 17138
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19720 16590 19748 16934
rect 19948 16892 20256 16901
rect 19948 16890 19954 16892
rect 20010 16890 20034 16892
rect 20090 16890 20114 16892
rect 20170 16890 20194 16892
rect 20250 16890 20256 16892
rect 20010 16838 20012 16890
rect 20192 16838 20194 16890
rect 19948 16836 19954 16838
rect 20010 16836 20034 16838
rect 20090 16836 20114 16838
rect 20170 16836 20194 16838
rect 20250 16836 20256 16838
rect 19948 16827 20256 16836
rect 19708 16584 19760 16590
rect 19708 16526 19760 16532
rect 19616 16516 19668 16522
rect 19616 16458 19668 16464
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19352 15026 19380 15438
rect 19536 15162 19564 16050
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 18892 9586 18920 13806
rect 18984 13326 19012 13806
rect 18972 13320 19024 13326
rect 18972 13262 19024 13268
rect 18984 13190 19012 13262
rect 19260 13258 19288 14894
rect 19248 13252 19300 13258
rect 19248 13194 19300 13200
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 18984 12646 19012 13126
rect 19064 12912 19116 12918
rect 19064 12854 19116 12860
rect 18972 12640 19024 12646
rect 18972 12582 19024 12588
rect 18984 11762 19012 12582
rect 18972 11756 19024 11762
rect 18972 11698 19024 11704
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18984 10266 19012 10406
rect 18972 10260 19024 10266
rect 18972 10202 19024 10208
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 18708 8974 18736 9522
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 19076 8498 19104 12854
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 19168 11762 19196 12038
rect 19156 11756 19208 11762
rect 19156 11698 19208 11704
rect 19260 10198 19288 13194
rect 19352 12764 19380 14962
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19432 14884 19484 14890
rect 19432 14826 19484 14832
rect 19444 13394 19472 14826
rect 19536 14414 19564 14894
rect 19628 14618 19656 16458
rect 19948 15804 20256 15813
rect 19948 15802 19954 15804
rect 20010 15802 20034 15804
rect 20090 15802 20114 15804
rect 20170 15802 20194 15804
rect 20250 15802 20256 15804
rect 20010 15750 20012 15802
rect 20192 15750 20194 15802
rect 19948 15748 19954 15750
rect 20010 15748 20034 15750
rect 20090 15748 20114 15750
rect 20170 15748 20194 15750
rect 20250 15748 20256 15750
rect 19948 15739 20256 15748
rect 20076 15632 20128 15638
rect 20076 15574 20128 15580
rect 19708 15428 19760 15434
rect 19708 15370 19760 15376
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 19720 14362 19748 15370
rect 20088 15026 20116 15574
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 19800 14884 19852 14890
rect 19800 14826 19852 14832
rect 19812 14618 19840 14826
rect 19948 14716 20256 14725
rect 19948 14714 19954 14716
rect 20010 14714 20034 14716
rect 20090 14714 20114 14716
rect 20170 14714 20194 14716
rect 20250 14714 20256 14716
rect 20010 14662 20012 14714
rect 20192 14662 20194 14714
rect 19948 14660 19954 14662
rect 20010 14660 20034 14662
rect 20090 14660 20114 14662
rect 20170 14660 20194 14662
rect 20250 14660 20256 14662
rect 19948 14651 20256 14660
rect 19800 14612 19852 14618
rect 19800 14554 19852 14560
rect 20260 14544 20312 14550
rect 20260 14486 20312 14492
rect 19720 14334 19840 14362
rect 19812 14278 19840 14334
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19536 12918 19564 13806
rect 19708 13456 19760 13462
rect 19708 13398 19760 13404
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 19352 12736 19564 12764
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19352 12102 19380 12582
rect 19432 12164 19484 12170
rect 19432 12106 19484 12112
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19352 11898 19380 12038
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19248 10192 19300 10198
rect 19248 10134 19300 10140
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18328 8016 18380 8022
rect 18328 7958 18380 7964
rect 18340 7410 18368 7958
rect 18800 7886 18828 8298
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18432 7546 18460 7822
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18800 7410 18828 7822
rect 19260 7546 19288 10134
rect 19352 9042 19380 10610
rect 19444 10146 19472 12106
rect 19536 11898 19564 12736
rect 19628 12306 19656 12786
rect 19616 12300 19668 12306
rect 19616 12242 19668 12248
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19628 11762 19656 12242
rect 19616 11756 19668 11762
rect 19616 11698 19668 11704
rect 19720 10606 19748 13398
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19812 10266 19840 14214
rect 20272 13818 20300 14486
rect 20364 13938 20392 21286
rect 20444 20868 20496 20874
rect 20444 20810 20496 20816
rect 20456 20534 20484 20810
rect 22662 20700 22970 20709
rect 22662 20698 22668 20700
rect 22724 20698 22748 20700
rect 22804 20698 22828 20700
rect 22884 20698 22908 20700
rect 22964 20698 22970 20700
rect 22724 20646 22726 20698
rect 22906 20646 22908 20698
rect 22662 20644 22668 20646
rect 22724 20644 22748 20646
rect 22804 20644 22828 20646
rect 22884 20644 22908 20646
rect 22964 20644 22970 20646
rect 22662 20635 22970 20644
rect 20444 20528 20496 20534
rect 20444 20470 20496 20476
rect 20456 18834 20484 20470
rect 22662 19612 22970 19621
rect 22662 19610 22668 19612
rect 22724 19610 22748 19612
rect 22804 19610 22828 19612
rect 22884 19610 22908 19612
rect 22964 19610 22970 19612
rect 22724 19558 22726 19610
rect 22906 19558 22908 19610
rect 22662 19556 22668 19558
rect 22724 19556 22748 19558
rect 22804 19556 22828 19558
rect 22884 19556 22908 19558
rect 22964 19556 22970 19558
rect 22662 19547 22970 19556
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20456 18290 20484 18770
rect 20996 18692 21048 18698
rect 20996 18634 21048 18640
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 21008 17202 21036 18634
rect 22662 18524 22970 18533
rect 22662 18522 22668 18524
rect 22724 18522 22748 18524
rect 22804 18522 22828 18524
rect 22884 18522 22908 18524
rect 22964 18522 22970 18524
rect 22724 18470 22726 18522
rect 22906 18470 22908 18522
rect 22662 18468 22668 18470
rect 22724 18468 22748 18470
rect 22804 18468 22828 18470
rect 22884 18468 22908 18470
rect 22964 18468 22970 18470
rect 22662 18459 22970 18468
rect 22662 17436 22970 17445
rect 22662 17434 22668 17436
rect 22724 17434 22748 17436
rect 22804 17434 22828 17436
rect 22884 17434 22908 17436
rect 22964 17434 22970 17436
rect 22724 17382 22726 17434
rect 22906 17382 22908 17434
rect 22662 17380 22668 17382
rect 22724 17380 22748 17382
rect 22804 17380 22828 17382
rect 22884 17380 22908 17382
rect 22964 17380 22970 17382
rect 22662 17371 22970 17380
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20916 16114 20944 16934
rect 22662 16348 22970 16357
rect 22662 16346 22668 16348
rect 22724 16346 22748 16348
rect 22804 16346 22828 16348
rect 22884 16346 22908 16348
rect 22964 16346 22970 16348
rect 22724 16294 22726 16346
rect 22906 16294 22908 16346
rect 22662 16292 22668 16294
rect 22724 16292 22748 16294
rect 22804 16292 22828 16294
rect 22884 16292 22908 16294
rect 22964 16292 22970 16294
rect 22662 16283 22970 16292
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 22662 15260 22970 15269
rect 22662 15258 22668 15260
rect 22724 15258 22748 15260
rect 22804 15258 22828 15260
rect 22884 15258 22908 15260
rect 22964 15258 22970 15260
rect 22724 15206 22726 15258
rect 22906 15206 22908 15258
rect 22662 15204 22668 15206
rect 22724 15204 22748 15206
rect 22804 15204 22828 15206
rect 22884 15204 22908 15206
rect 22964 15204 22970 15206
rect 22662 15195 22970 15204
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20272 13790 20392 13818
rect 19948 13628 20256 13637
rect 19948 13626 19954 13628
rect 20010 13626 20034 13628
rect 20090 13626 20114 13628
rect 20170 13626 20194 13628
rect 20250 13626 20256 13628
rect 20010 13574 20012 13626
rect 20192 13574 20194 13626
rect 19948 13572 19954 13574
rect 20010 13572 20034 13574
rect 20090 13572 20114 13574
rect 20170 13572 20194 13574
rect 20250 13572 20256 13574
rect 19948 13563 20256 13572
rect 19892 13388 19944 13394
rect 19892 13330 19944 13336
rect 19904 12986 19932 13330
rect 19892 12980 19944 12986
rect 19892 12922 19944 12928
rect 19904 12646 19932 12922
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 19948 12540 20256 12549
rect 19948 12538 19954 12540
rect 20010 12538 20034 12540
rect 20090 12538 20114 12540
rect 20170 12538 20194 12540
rect 20250 12538 20256 12540
rect 20010 12486 20012 12538
rect 20192 12486 20194 12538
rect 19948 12484 19954 12486
rect 20010 12484 20034 12486
rect 20090 12484 20114 12486
rect 20170 12484 20194 12486
rect 20250 12484 20256 12486
rect 19948 12475 20256 12484
rect 19892 12300 19944 12306
rect 19892 12242 19944 12248
rect 19904 12102 19932 12242
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 19948 11452 20256 11461
rect 19948 11450 19954 11452
rect 20010 11450 20034 11452
rect 20090 11450 20114 11452
rect 20170 11450 20194 11452
rect 20250 11450 20256 11452
rect 20010 11398 20012 11450
rect 20192 11398 20194 11450
rect 19948 11396 19954 11398
rect 20010 11396 20034 11398
rect 20090 11396 20114 11398
rect 20170 11396 20194 11398
rect 20250 11396 20256 11398
rect 19948 11387 20256 11396
rect 19948 10364 20256 10373
rect 19948 10362 19954 10364
rect 20010 10362 20034 10364
rect 20090 10362 20114 10364
rect 20170 10362 20194 10364
rect 20250 10362 20256 10364
rect 20010 10310 20012 10362
rect 20192 10310 20194 10362
rect 19948 10308 19954 10310
rect 20010 10308 20034 10310
rect 20090 10308 20114 10310
rect 20170 10308 20194 10310
rect 20250 10308 20256 10310
rect 19948 10299 20256 10308
rect 19800 10260 19852 10266
rect 19800 10202 19852 10208
rect 19444 10118 19564 10146
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19444 9178 19472 9998
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19352 8362 19380 8978
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19536 7954 19564 10118
rect 20364 9926 20392 13790
rect 20456 10674 20484 14282
rect 22662 14172 22970 14181
rect 22662 14170 22668 14172
rect 22724 14170 22748 14172
rect 22804 14170 22828 14172
rect 22884 14170 22908 14172
rect 22964 14170 22970 14172
rect 22724 14118 22726 14170
rect 22906 14118 22908 14170
rect 22662 14116 22668 14118
rect 22724 14116 22748 14118
rect 22804 14116 22828 14118
rect 22884 14116 22908 14118
rect 22964 14116 22970 14118
rect 22662 14107 22970 14116
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 20352 9920 20404 9926
rect 20352 9862 20404 9868
rect 19948 9276 20256 9285
rect 19948 9274 19954 9276
rect 20010 9274 20034 9276
rect 20090 9274 20114 9276
rect 20170 9274 20194 9276
rect 20250 9274 20256 9276
rect 20010 9222 20012 9274
rect 20192 9222 20194 9274
rect 19948 9220 19954 9222
rect 20010 9220 20034 9222
rect 20090 9220 20114 9222
rect 20170 9220 20194 9222
rect 20250 9220 20256 9222
rect 19948 9211 20256 9220
rect 19948 8188 20256 8197
rect 19948 8186 19954 8188
rect 20010 8186 20034 8188
rect 20090 8186 20114 8188
rect 20170 8186 20194 8188
rect 20250 8186 20256 8188
rect 20010 8134 20012 8186
rect 20192 8134 20194 8186
rect 19948 8132 19954 8134
rect 20010 8132 20034 8134
rect 20090 8132 20114 8134
rect 20170 8132 20194 8134
rect 20250 8132 20256 8134
rect 19948 8123 20256 8132
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19536 7478 19564 7890
rect 19524 7472 19576 7478
rect 19524 7414 19576 7420
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 19948 7100 20256 7109
rect 19948 7098 19954 7100
rect 20010 7098 20034 7100
rect 20090 7098 20114 7100
rect 20170 7098 20194 7100
rect 20250 7098 20256 7100
rect 20010 7046 20012 7098
rect 20192 7046 20194 7098
rect 19948 7044 19954 7046
rect 20010 7044 20034 7046
rect 20090 7044 20114 7046
rect 20170 7044 20194 7046
rect 20250 7044 20256 7046
rect 19948 7035 20256 7044
rect 18236 6928 18288 6934
rect 18236 6870 18288 6876
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 11806 6556 12114 6565
rect 11806 6554 11812 6556
rect 11868 6554 11892 6556
rect 11948 6554 11972 6556
rect 12028 6554 12052 6556
rect 12108 6554 12114 6556
rect 11868 6502 11870 6554
rect 12050 6502 12052 6554
rect 11806 6500 11812 6502
rect 11868 6500 11892 6502
rect 11948 6500 11972 6502
rect 12028 6500 12052 6502
rect 12108 6500 12114 6502
rect 11806 6491 12114 6500
rect 17234 6556 17542 6565
rect 17234 6554 17240 6556
rect 17296 6554 17320 6556
rect 17376 6554 17400 6556
rect 17456 6554 17480 6556
rect 17536 6554 17542 6556
rect 17296 6502 17298 6554
rect 17478 6502 17480 6554
rect 17234 6500 17240 6502
rect 17296 6500 17320 6502
rect 17376 6500 17400 6502
rect 17456 6500 17480 6502
rect 17536 6500 17542 6502
rect 17234 6491 17542 6500
rect 14520 6012 14828 6021
rect 14520 6010 14526 6012
rect 14582 6010 14606 6012
rect 14662 6010 14686 6012
rect 14742 6010 14766 6012
rect 14822 6010 14828 6012
rect 14582 5958 14584 6010
rect 14764 5958 14766 6010
rect 14520 5956 14526 5958
rect 14582 5956 14606 5958
rect 14662 5956 14686 5958
rect 14742 5956 14766 5958
rect 14822 5956 14828 5958
rect 14520 5947 14828 5956
rect 19948 6012 20256 6021
rect 19948 6010 19954 6012
rect 20010 6010 20034 6012
rect 20090 6010 20114 6012
rect 20170 6010 20194 6012
rect 20250 6010 20256 6012
rect 20010 5958 20012 6010
rect 20192 5958 20194 6010
rect 19948 5956 19954 5958
rect 20010 5956 20034 5958
rect 20090 5956 20114 5958
rect 20170 5956 20194 5958
rect 20250 5956 20256 5958
rect 19948 5947 20256 5956
rect 11806 5468 12114 5477
rect 11806 5466 11812 5468
rect 11868 5466 11892 5468
rect 11948 5466 11972 5468
rect 12028 5466 12052 5468
rect 12108 5466 12114 5468
rect 11868 5414 11870 5466
rect 12050 5414 12052 5466
rect 11806 5412 11812 5414
rect 11868 5412 11892 5414
rect 11948 5412 11972 5414
rect 12028 5412 12052 5414
rect 12108 5412 12114 5414
rect 11806 5403 12114 5412
rect 17234 5468 17542 5477
rect 17234 5466 17240 5468
rect 17296 5466 17320 5468
rect 17376 5466 17400 5468
rect 17456 5466 17480 5468
rect 17536 5466 17542 5468
rect 17296 5414 17298 5466
rect 17478 5414 17480 5466
rect 17234 5412 17240 5414
rect 17296 5412 17320 5414
rect 17376 5412 17400 5414
rect 17456 5412 17480 5414
rect 17536 5412 17542 5414
rect 17234 5403 17542 5412
rect 14520 4924 14828 4933
rect 14520 4922 14526 4924
rect 14582 4922 14606 4924
rect 14662 4922 14686 4924
rect 14742 4922 14766 4924
rect 14822 4922 14828 4924
rect 14582 4870 14584 4922
rect 14764 4870 14766 4922
rect 14520 4868 14526 4870
rect 14582 4868 14606 4870
rect 14662 4868 14686 4870
rect 14742 4868 14766 4870
rect 14822 4868 14828 4870
rect 14520 4859 14828 4868
rect 19948 4924 20256 4933
rect 19948 4922 19954 4924
rect 20010 4922 20034 4924
rect 20090 4922 20114 4924
rect 20170 4922 20194 4924
rect 20250 4922 20256 4924
rect 20010 4870 20012 4922
rect 20192 4870 20194 4922
rect 19948 4868 19954 4870
rect 20010 4868 20034 4870
rect 20090 4868 20114 4870
rect 20170 4868 20194 4870
rect 20250 4868 20256 4870
rect 19948 4859 20256 4868
rect 11806 4380 12114 4389
rect 11806 4378 11812 4380
rect 11868 4378 11892 4380
rect 11948 4378 11972 4380
rect 12028 4378 12052 4380
rect 12108 4378 12114 4380
rect 11868 4326 11870 4378
rect 12050 4326 12052 4378
rect 11806 4324 11812 4326
rect 11868 4324 11892 4326
rect 11948 4324 11972 4326
rect 12028 4324 12052 4326
rect 12108 4324 12114 4326
rect 11806 4315 12114 4324
rect 17234 4380 17542 4389
rect 17234 4378 17240 4380
rect 17296 4378 17320 4380
rect 17376 4378 17400 4380
rect 17456 4378 17480 4380
rect 17536 4378 17542 4380
rect 17296 4326 17298 4378
rect 17478 4326 17480 4378
rect 17234 4324 17240 4326
rect 17296 4324 17320 4326
rect 17376 4324 17400 4326
rect 17456 4324 17480 4326
rect 17536 4324 17542 4326
rect 17234 4315 17542 4324
rect 14520 3836 14828 3845
rect 14520 3834 14526 3836
rect 14582 3834 14606 3836
rect 14662 3834 14686 3836
rect 14742 3834 14766 3836
rect 14822 3834 14828 3836
rect 14582 3782 14584 3834
rect 14764 3782 14766 3834
rect 14520 3780 14526 3782
rect 14582 3780 14606 3782
rect 14662 3780 14686 3782
rect 14742 3780 14766 3782
rect 14822 3780 14828 3782
rect 14520 3771 14828 3780
rect 19948 3836 20256 3845
rect 19948 3834 19954 3836
rect 20010 3834 20034 3836
rect 20090 3834 20114 3836
rect 20170 3834 20194 3836
rect 20250 3834 20256 3836
rect 20010 3782 20012 3834
rect 20192 3782 20194 3834
rect 19948 3780 19954 3782
rect 20010 3780 20034 3782
rect 20090 3780 20114 3782
rect 20170 3780 20194 3782
rect 20250 3780 20256 3782
rect 19948 3771 20256 3780
rect 11806 3292 12114 3301
rect 11806 3290 11812 3292
rect 11868 3290 11892 3292
rect 11948 3290 11972 3292
rect 12028 3290 12052 3292
rect 12108 3290 12114 3292
rect 11868 3238 11870 3290
rect 12050 3238 12052 3290
rect 11806 3236 11812 3238
rect 11868 3236 11892 3238
rect 11948 3236 11972 3238
rect 12028 3236 12052 3238
rect 12108 3236 12114 3238
rect 11806 3227 12114 3236
rect 17234 3292 17542 3301
rect 17234 3290 17240 3292
rect 17296 3290 17320 3292
rect 17376 3290 17400 3292
rect 17456 3290 17480 3292
rect 17536 3290 17542 3292
rect 17296 3238 17298 3290
rect 17478 3238 17480 3290
rect 17234 3236 17240 3238
rect 17296 3236 17320 3238
rect 17376 3236 17400 3238
rect 17456 3236 17480 3238
rect 17536 3236 17542 3238
rect 17234 3227 17542 3236
rect 14520 2748 14828 2757
rect 14520 2746 14526 2748
rect 14582 2746 14606 2748
rect 14662 2746 14686 2748
rect 14742 2746 14766 2748
rect 14822 2746 14828 2748
rect 14582 2694 14584 2746
rect 14764 2694 14766 2746
rect 14520 2692 14526 2694
rect 14582 2692 14606 2694
rect 14662 2692 14686 2694
rect 14742 2692 14766 2694
rect 14822 2692 14828 2694
rect 14520 2683 14828 2692
rect 19948 2748 20256 2757
rect 19948 2746 19954 2748
rect 20010 2746 20034 2748
rect 20090 2746 20114 2748
rect 20170 2746 20194 2748
rect 20250 2746 20256 2748
rect 20010 2694 20012 2746
rect 20192 2694 20194 2746
rect 19948 2692 19954 2694
rect 20010 2692 20034 2694
rect 20090 2692 20114 2694
rect 20170 2692 20194 2694
rect 20250 2692 20256 2694
rect 19948 2683 20256 2692
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 8852 2508 8904 2514
rect 8852 2450 8904 2456
rect 21008 2446 21036 14010
rect 22662 13084 22970 13093
rect 22662 13082 22668 13084
rect 22724 13082 22748 13084
rect 22804 13082 22828 13084
rect 22884 13082 22908 13084
rect 22964 13082 22970 13084
rect 22724 13030 22726 13082
rect 22906 13030 22908 13082
rect 22662 13028 22668 13030
rect 22724 13028 22748 13030
rect 22804 13028 22828 13030
rect 22884 13028 22908 13030
rect 22964 13028 22970 13030
rect 22662 13019 22970 13028
rect 22662 11996 22970 12005
rect 22662 11994 22668 11996
rect 22724 11994 22748 11996
rect 22804 11994 22828 11996
rect 22884 11994 22908 11996
rect 22964 11994 22970 11996
rect 22724 11942 22726 11994
rect 22906 11942 22908 11994
rect 22662 11940 22668 11942
rect 22724 11940 22748 11942
rect 22804 11940 22828 11942
rect 22884 11940 22908 11942
rect 22964 11940 22970 11942
rect 22662 11931 22970 11940
rect 22662 10908 22970 10917
rect 22662 10906 22668 10908
rect 22724 10906 22748 10908
rect 22804 10906 22828 10908
rect 22884 10906 22908 10908
rect 22964 10906 22970 10908
rect 22724 10854 22726 10906
rect 22906 10854 22908 10906
rect 22662 10852 22668 10854
rect 22724 10852 22748 10854
rect 22804 10852 22828 10854
rect 22884 10852 22908 10854
rect 22964 10852 22970 10854
rect 22662 10843 22970 10852
rect 22662 9820 22970 9829
rect 22662 9818 22668 9820
rect 22724 9818 22748 9820
rect 22804 9818 22828 9820
rect 22884 9818 22908 9820
rect 22964 9818 22970 9820
rect 22724 9766 22726 9818
rect 22906 9766 22908 9818
rect 22662 9764 22668 9766
rect 22724 9764 22748 9766
rect 22804 9764 22828 9766
rect 22884 9764 22908 9766
rect 22964 9764 22970 9766
rect 22662 9755 22970 9764
rect 22662 8732 22970 8741
rect 22662 8730 22668 8732
rect 22724 8730 22748 8732
rect 22804 8730 22828 8732
rect 22884 8730 22908 8732
rect 22964 8730 22970 8732
rect 22724 8678 22726 8730
rect 22906 8678 22908 8730
rect 22662 8676 22668 8678
rect 22724 8676 22748 8678
rect 22804 8676 22828 8678
rect 22884 8676 22908 8678
rect 22964 8676 22970 8678
rect 22662 8667 22970 8676
rect 22662 7644 22970 7653
rect 22662 7642 22668 7644
rect 22724 7642 22748 7644
rect 22804 7642 22828 7644
rect 22884 7642 22908 7644
rect 22964 7642 22970 7644
rect 22724 7590 22726 7642
rect 22906 7590 22908 7642
rect 22662 7588 22668 7590
rect 22724 7588 22748 7590
rect 22804 7588 22828 7590
rect 22884 7588 22908 7590
rect 22964 7588 22970 7590
rect 22662 7579 22970 7588
rect 22662 6556 22970 6565
rect 22662 6554 22668 6556
rect 22724 6554 22748 6556
rect 22804 6554 22828 6556
rect 22884 6554 22908 6556
rect 22964 6554 22970 6556
rect 22724 6502 22726 6554
rect 22906 6502 22908 6554
rect 22662 6500 22668 6502
rect 22724 6500 22748 6502
rect 22804 6500 22828 6502
rect 22884 6500 22908 6502
rect 22964 6500 22970 6502
rect 22662 6491 22970 6500
rect 22662 5468 22970 5477
rect 22662 5466 22668 5468
rect 22724 5466 22748 5468
rect 22804 5466 22828 5468
rect 22884 5466 22908 5468
rect 22964 5466 22970 5468
rect 22724 5414 22726 5466
rect 22906 5414 22908 5466
rect 22662 5412 22668 5414
rect 22724 5412 22748 5414
rect 22804 5412 22828 5414
rect 22884 5412 22908 5414
rect 22964 5412 22970 5414
rect 22662 5403 22970 5412
rect 22662 4380 22970 4389
rect 22662 4378 22668 4380
rect 22724 4378 22748 4380
rect 22804 4378 22828 4380
rect 22884 4378 22908 4380
rect 22964 4378 22970 4380
rect 22724 4326 22726 4378
rect 22906 4326 22908 4378
rect 22662 4324 22668 4326
rect 22724 4324 22748 4326
rect 22804 4324 22828 4326
rect 22884 4324 22908 4326
rect 22964 4324 22970 4326
rect 22662 4315 22970 4324
rect 22662 3292 22970 3301
rect 22662 3290 22668 3292
rect 22724 3290 22748 3292
rect 22804 3290 22828 3292
rect 22884 3290 22908 3292
rect 22964 3290 22970 3292
rect 22724 3238 22726 3290
rect 22906 3238 22908 3290
rect 22662 3236 22668 3238
rect 22724 3236 22748 3238
rect 22804 3236 22828 3238
rect 22884 3236 22908 3238
rect 22964 3236 22970 3238
rect 22662 3227 22970 3236
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 1676 2372 1728 2378
rect 1676 2314 1728 2320
rect 4620 2372 4672 2378
rect 4620 2314 4672 2320
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 10508 2372 10560 2378
rect 10508 2314 10560 2320
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 16580 2372 16632 2378
rect 16580 2314 16632 2320
rect 19340 2372 19392 2378
rect 19340 2314 19392 2320
rect 22284 2372 22336 2378
rect 22284 2314 22336 2320
rect 1688 800 1716 2314
rect 4632 800 4660 2314
rect 6378 2204 6686 2213
rect 6378 2202 6384 2204
rect 6440 2202 6464 2204
rect 6520 2202 6544 2204
rect 6600 2202 6624 2204
rect 6680 2202 6686 2204
rect 6440 2150 6442 2202
rect 6622 2150 6624 2202
rect 6378 2148 6384 2150
rect 6440 2148 6464 2150
rect 6520 2148 6544 2150
rect 6600 2148 6624 2150
rect 6680 2148 6686 2150
rect 6378 2139 6686 2148
rect 7576 800 7604 2314
rect 10520 800 10548 2314
rect 11806 2204 12114 2213
rect 11806 2202 11812 2204
rect 11868 2202 11892 2204
rect 11948 2202 11972 2204
rect 12028 2202 12052 2204
rect 12108 2202 12114 2204
rect 11868 2150 11870 2202
rect 12050 2150 12052 2202
rect 11806 2148 11812 2150
rect 11868 2148 11892 2150
rect 11948 2148 11972 2150
rect 12028 2148 12052 2150
rect 12108 2148 12114 2150
rect 11806 2139 12114 2148
rect 13832 898 13860 2314
rect 16592 898 16620 2314
rect 17234 2204 17542 2213
rect 17234 2202 17240 2204
rect 17296 2202 17320 2204
rect 17376 2202 17400 2204
rect 17456 2202 17480 2204
rect 17536 2202 17542 2204
rect 17296 2150 17298 2202
rect 17478 2150 17480 2202
rect 17234 2148 17240 2150
rect 17296 2148 17320 2150
rect 17376 2148 17400 2150
rect 17456 2148 17480 2150
rect 17536 2148 17542 2150
rect 17234 2139 17542 2148
rect 13464 870 13860 898
rect 16408 870 16620 898
rect 13464 800 13492 870
rect 16408 800 16436 870
rect 19352 800 19380 2314
rect 22296 800 22324 2314
rect 22662 2204 22970 2213
rect 22662 2202 22668 2204
rect 22724 2202 22748 2204
rect 22804 2202 22828 2204
rect 22884 2202 22908 2204
rect 22964 2202 22970 2204
rect 22724 2150 22726 2202
rect 22906 2150 22908 2202
rect 22662 2148 22668 2150
rect 22724 2148 22748 2150
rect 22804 2148 22828 2150
rect 22884 2148 22908 2150
rect 22964 2148 22970 2150
rect 22662 2139 22970 2148
rect 1674 0 1730 800
rect 4618 0 4674 800
rect 7562 0 7618 800
rect 10506 0 10562 800
rect 13450 0 13506 800
rect 16394 0 16450 800
rect 19338 0 19394 800
rect 22282 0 22338 800
<< via2 >>
rect 3670 21242 3726 21244
rect 3750 21242 3806 21244
rect 3830 21242 3886 21244
rect 3910 21242 3966 21244
rect 3670 21190 3716 21242
rect 3716 21190 3726 21242
rect 3750 21190 3780 21242
rect 3780 21190 3792 21242
rect 3792 21190 3806 21242
rect 3830 21190 3844 21242
rect 3844 21190 3856 21242
rect 3856 21190 3886 21242
rect 3910 21190 3920 21242
rect 3920 21190 3966 21242
rect 3670 21188 3726 21190
rect 3750 21188 3806 21190
rect 3830 21188 3886 21190
rect 3910 21188 3966 21190
rect 3670 20154 3726 20156
rect 3750 20154 3806 20156
rect 3830 20154 3886 20156
rect 3910 20154 3966 20156
rect 3670 20102 3716 20154
rect 3716 20102 3726 20154
rect 3750 20102 3780 20154
rect 3780 20102 3792 20154
rect 3792 20102 3806 20154
rect 3830 20102 3844 20154
rect 3844 20102 3856 20154
rect 3856 20102 3886 20154
rect 3910 20102 3920 20154
rect 3920 20102 3966 20154
rect 3670 20100 3726 20102
rect 3750 20100 3806 20102
rect 3830 20100 3886 20102
rect 3910 20100 3966 20102
rect 6384 21786 6440 21788
rect 6464 21786 6520 21788
rect 6544 21786 6600 21788
rect 6624 21786 6680 21788
rect 6384 21734 6430 21786
rect 6430 21734 6440 21786
rect 6464 21734 6494 21786
rect 6494 21734 6506 21786
rect 6506 21734 6520 21786
rect 6544 21734 6558 21786
rect 6558 21734 6570 21786
rect 6570 21734 6600 21786
rect 6624 21734 6634 21786
rect 6634 21734 6680 21786
rect 6384 21732 6440 21734
rect 6464 21732 6520 21734
rect 6544 21732 6600 21734
rect 6624 21732 6680 21734
rect 11812 21786 11868 21788
rect 11892 21786 11948 21788
rect 11972 21786 12028 21788
rect 12052 21786 12108 21788
rect 11812 21734 11858 21786
rect 11858 21734 11868 21786
rect 11892 21734 11922 21786
rect 11922 21734 11934 21786
rect 11934 21734 11948 21786
rect 11972 21734 11986 21786
rect 11986 21734 11998 21786
rect 11998 21734 12028 21786
rect 12052 21734 12062 21786
rect 12062 21734 12108 21786
rect 11812 21732 11868 21734
rect 11892 21732 11948 21734
rect 11972 21732 12028 21734
rect 12052 21732 12108 21734
rect 17240 21786 17296 21788
rect 17320 21786 17376 21788
rect 17400 21786 17456 21788
rect 17480 21786 17536 21788
rect 17240 21734 17286 21786
rect 17286 21734 17296 21786
rect 17320 21734 17350 21786
rect 17350 21734 17362 21786
rect 17362 21734 17376 21786
rect 17400 21734 17414 21786
rect 17414 21734 17426 21786
rect 17426 21734 17456 21786
rect 17480 21734 17490 21786
rect 17490 21734 17536 21786
rect 17240 21732 17296 21734
rect 17320 21732 17376 21734
rect 17400 21732 17456 21734
rect 17480 21732 17536 21734
rect 22668 21786 22724 21788
rect 22748 21786 22804 21788
rect 22828 21786 22884 21788
rect 22908 21786 22964 21788
rect 22668 21734 22714 21786
rect 22714 21734 22724 21786
rect 22748 21734 22778 21786
rect 22778 21734 22790 21786
rect 22790 21734 22804 21786
rect 22828 21734 22842 21786
rect 22842 21734 22854 21786
rect 22854 21734 22884 21786
rect 22908 21734 22918 21786
rect 22918 21734 22964 21786
rect 22668 21732 22724 21734
rect 22748 21732 22804 21734
rect 22828 21732 22884 21734
rect 22908 21732 22964 21734
rect 9098 21242 9154 21244
rect 9178 21242 9234 21244
rect 9258 21242 9314 21244
rect 9338 21242 9394 21244
rect 9098 21190 9144 21242
rect 9144 21190 9154 21242
rect 9178 21190 9208 21242
rect 9208 21190 9220 21242
rect 9220 21190 9234 21242
rect 9258 21190 9272 21242
rect 9272 21190 9284 21242
rect 9284 21190 9314 21242
rect 9338 21190 9348 21242
rect 9348 21190 9394 21242
rect 9098 21188 9154 21190
rect 9178 21188 9234 21190
rect 9258 21188 9314 21190
rect 9338 21188 9394 21190
rect 14526 21242 14582 21244
rect 14606 21242 14662 21244
rect 14686 21242 14742 21244
rect 14766 21242 14822 21244
rect 14526 21190 14572 21242
rect 14572 21190 14582 21242
rect 14606 21190 14636 21242
rect 14636 21190 14648 21242
rect 14648 21190 14662 21242
rect 14686 21190 14700 21242
rect 14700 21190 14712 21242
rect 14712 21190 14742 21242
rect 14766 21190 14776 21242
rect 14776 21190 14822 21242
rect 14526 21188 14582 21190
rect 14606 21188 14662 21190
rect 14686 21188 14742 21190
rect 14766 21188 14822 21190
rect 6384 20698 6440 20700
rect 6464 20698 6520 20700
rect 6544 20698 6600 20700
rect 6624 20698 6680 20700
rect 6384 20646 6430 20698
rect 6430 20646 6440 20698
rect 6464 20646 6494 20698
rect 6494 20646 6506 20698
rect 6506 20646 6520 20698
rect 6544 20646 6558 20698
rect 6558 20646 6570 20698
rect 6570 20646 6600 20698
rect 6624 20646 6634 20698
rect 6634 20646 6680 20698
rect 6384 20644 6440 20646
rect 6464 20644 6520 20646
rect 6544 20644 6600 20646
rect 6624 20644 6680 20646
rect 11812 20698 11868 20700
rect 11892 20698 11948 20700
rect 11972 20698 12028 20700
rect 12052 20698 12108 20700
rect 11812 20646 11858 20698
rect 11858 20646 11868 20698
rect 11892 20646 11922 20698
rect 11922 20646 11934 20698
rect 11934 20646 11948 20698
rect 11972 20646 11986 20698
rect 11986 20646 11998 20698
rect 11998 20646 12028 20698
rect 12052 20646 12062 20698
rect 12062 20646 12108 20698
rect 11812 20644 11868 20646
rect 11892 20644 11948 20646
rect 11972 20644 12028 20646
rect 12052 20644 12108 20646
rect 3670 19066 3726 19068
rect 3750 19066 3806 19068
rect 3830 19066 3886 19068
rect 3910 19066 3966 19068
rect 3670 19014 3716 19066
rect 3716 19014 3726 19066
rect 3750 19014 3780 19066
rect 3780 19014 3792 19066
rect 3792 19014 3806 19066
rect 3830 19014 3844 19066
rect 3844 19014 3856 19066
rect 3856 19014 3886 19066
rect 3910 19014 3920 19066
rect 3920 19014 3966 19066
rect 3670 19012 3726 19014
rect 3750 19012 3806 19014
rect 3830 19012 3886 19014
rect 3910 19012 3966 19014
rect 6384 19610 6440 19612
rect 6464 19610 6520 19612
rect 6544 19610 6600 19612
rect 6624 19610 6680 19612
rect 6384 19558 6430 19610
rect 6430 19558 6440 19610
rect 6464 19558 6494 19610
rect 6494 19558 6506 19610
rect 6506 19558 6520 19610
rect 6544 19558 6558 19610
rect 6558 19558 6570 19610
rect 6570 19558 6600 19610
rect 6624 19558 6634 19610
rect 6634 19558 6680 19610
rect 6384 19556 6440 19558
rect 6464 19556 6520 19558
rect 6544 19556 6600 19558
rect 6624 19556 6680 19558
rect 9098 20154 9154 20156
rect 9178 20154 9234 20156
rect 9258 20154 9314 20156
rect 9338 20154 9394 20156
rect 9098 20102 9144 20154
rect 9144 20102 9154 20154
rect 9178 20102 9208 20154
rect 9208 20102 9220 20154
rect 9220 20102 9234 20154
rect 9258 20102 9272 20154
rect 9272 20102 9284 20154
rect 9284 20102 9314 20154
rect 9338 20102 9348 20154
rect 9348 20102 9394 20154
rect 9098 20100 9154 20102
rect 9178 20100 9234 20102
rect 9258 20100 9314 20102
rect 9338 20100 9394 20102
rect 6384 18522 6440 18524
rect 6464 18522 6520 18524
rect 6544 18522 6600 18524
rect 6624 18522 6680 18524
rect 6384 18470 6430 18522
rect 6430 18470 6440 18522
rect 6464 18470 6494 18522
rect 6494 18470 6506 18522
rect 6506 18470 6520 18522
rect 6544 18470 6558 18522
rect 6558 18470 6570 18522
rect 6570 18470 6600 18522
rect 6624 18470 6634 18522
rect 6634 18470 6680 18522
rect 6384 18468 6440 18470
rect 6464 18468 6520 18470
rect 6544 18468 6600 18470
rect 6624 18468 6680 18470
rect 3670 17978 3726 17980
rect 3750 17978 3806 17980
rect 3830 17978 3886 17980
rect 3910 17978 3966 17980
rect 3670 17926 3716 17978
rect 3716 17926 3726 17978
rect 3750 17926 3780 17978
rect 3780 17926 3792 17978
rect 3792 17926 3806 17978
rect 3830 17926 3844 17978
rect 3844 17926 3856 17978
rect 3856 17926 3886 17978
rect 3910 17926 3920 17978
rect 3920 17926 3966 17978
rect 3670 17924 3726 17926
rect 3750 17924 3806 17926
rect 3830 17924 3886 17926
rect 3910 17924 3966 17926
rect 6384 17434 6440 17436
rect 6464 17434 6520 17436
rect 6544 17434 6600 17436
rect 6624 17434 6680 17436
rect 6384 17382 6430 17434
rect 6430 17382 6440 17434
rect 6464 17382 6494 17434
rect 6494 17382 6506 17434
rect 6506 17382 6520 17434
rect 6544 17382 6558 17434
rect 6558 17382 6570 17434
rect 6570 17382 6600 17434
rect 6624 17382 6634 17434
rect 6634 17382 6680 17434
rect 6384 17380 6440 17382
rect 6464 17380 6520 17382
rect 6544 17380 6600 17382
rect 6624 17380 6680 17382
rect 3670 16890 3726 16892
rect 3750 16890 3806 16892
rect 3830 16890 3886 16892
rect 3910 16890 3966 16892
rect 3670 16838 3716 16890
rect 3716 16838 3726 16890
rect 3750 16838 3780 16890
rect 3780 16838 3792 16890
rect 3792 16838 3806 16890
rect 3830 16838 3844 16890
rect 3844 16838 3856 16890
rect 3856 16838 3886 16890
rect 3910 16838 3920 16890
rect 3920 16838 3966 16890
rect 3670 16836 3726 16838
rect 3750 16836 3806 16838
rect 3830 16836 3886 16838
rect 3910 16836 3966 16838
rect 3670 15802 3726 15804
rect 3750 15802 3806 15804
rect 3830 15802 3886 15804
rect 3910 15802 3966 15804
rect 3670 15750 3716 15802
rect 3716 15750 3726 15802
rect 3750 15750 3780 15802
rect 3780 15750 3792 15802
rect 3792 15750 3806 15802
rect 3830 15750 3844 15802
rect 3844 15750 3856 15802
rect 3856 15750 3886 15802
rect 3910 15750 3920 15802
rect 3920 15750 3966 15802
rect 3670 15748 3726 15750
rect 3750 15748 3806 15750
rect 3830 15748 3886 15750
rect 3910 15748 3966 15750
rect 3670 14714 3726 14716
rect 3750 14714 3806 14716
rect 3830 14714 3886 14716
rect 3910 14714 3966 14716
rect 3670 14662 3716 14714
rect 3716 14662 3726 14714
rect 3750 14662 3780 14714
rect 3780 14662 3792 14714
rect 3792 14662 3806 14714
rect 3830 14662 3844 14714
rect 3844 14662 3856 14714
rect 3856 14662 3886 14714
rect 3910 14662 3920 14714
rect 3920 14662 3966 14714
rect 3670 14660 3726 14662
rect 3750 14660 3806 14662
rect 3830 14660 3886 14662
rect 3910 14660 3966 14662
rect 3670 13626 3726 13628
rect 3750 13626 3806 13628
rect 3830 13626 3886 13628
rect 3910 13626 3966 13628
rect 3670 13574 3716 13626
rect 3716 13574 3726 13626
rect 3750 13574 3780 13626
rect 3780 13574 3792 13626
rect 3792 13574 3806 13626
rect 3830 13574 3844 13626
rect 3844 13574 3856 13626
rect 3856 13574 3886 13626
rect 3910 13574 3920 13626
rect 3920 13574 3966 13626
rect 3670 13572 3726 13574
rect 3750 13572 3806 13574
rect 3830 13572 3886 13574
rect 3910 13572 3966 13574
rect 3670 12538 3726 12540
rect 3750 12538 3806 12540
rect 3830 12538 3886 12540
rect 3910 12538 3966 12540
rect 3670 12486 3716 12538
rect 3716 12486 3726 12538
rect 3750 12486 3780 12538
rect 3780 12486 3792 12538
rect 3792 12486 3806 12538
rect 3830 12486 3844 12538
rect 3844 12486 3856 12538
rect 3856 12486 3886 12538
rect 3910 12486 3920 12538
rect 3920 12486 3966 12538
rect 3670 12484 3726 12486
rect 3750 12484 3806 12486
rect 3830 12484 3886 12486
rect 3910 12484 3966 12486
rect 3670 11450 3726 11452
rect 3750 11450 3806 11452
rect 3830 11450 3886 11452
rect 3910 11450 3966 11452
rect 3670 11398 3716 11450
rect 3716 11398 3726 11450
rect 3750 11398 3780 11450
rect 3780 11398 3792 11450
rect 3792 11398 3806 11450
rect 3830 11398 3844 11450
rect 3844 11398 3856 11450
rect 3856 11398 3886 11450
rect 3910 11398 3920 11450
rect 3920 11398 3966 11450
rect 3670 11396 3726 11398
rect 3750 11396 3806 11398
rect 3830 11396 3886 11398
rect 3910 11396 3966 11398
rect 3670 10362 3726 10364
rect 3750 10362 3806 10364
rect 3830 10362 3886 10364
rect 3910 10362 3966 10364
rect 3670 10310 3716 10362
rect 3716 10310 3726 10362
rect 3750 10310 3780 10362
rect 3780 10310 3792 10362
rect 3792 10310 3806 10362
rect 3830 10310 3844 10362
rect 3844 10310 3856 10362
rect 3856 10310 3886 10362
rect 3910 10310 3920 10362
rect 3920 10310 3966 10362
rect 3670 10308 3726 10310
rect 3750 10308 3806 10310
rect 3830 10308 3886 10310
rect 3910 10308 3966 10310
rect 3670 9274 3726 9276
rect 3750 9274 3806 9276
rect 3830 9274 3886 9276
rect 3910 9274 3966 9276
rect 3670 9222 3716 9274
rect 3716 9222 3726 9274
rect 3750 9222 3780 9274
rect 3780 9222 3792 9274
rect 3792 9222 3806 9274
rect 3830 9222 3844 9274
rect 3844 9222 3856 9274
rect 3856 9222 3886 9274
rect 3910 9222 3920 9274
rect 3920 9222 3966 9274
rect 3670 9220 3726 9222
rect 3750 9220 3806 9222
rect 3830 9220 3886 9222
rect 3910 9220 3966 9222
rect 3670 8186 3726 8188
rect 3750 8186 3806 8188
rect 3830 8186 3886 8188
rect 3910 8186 3966 8188
rect 3670 8134 3716 8186
rect 3716 8134 3726 8186
rect 3750 8134 3780 8186
rect 3780 8134 3792 8186
rect 3792 8134 3806 8186
rect 3830 8134 3844 8186
rect 3844 8134 3856 8186
rect 3856 8134 3886 8186
rect 3910 8134 3920 8186
rect 3920 8134 3966 8186
rect 3670 8132 3726 8134
rect 3750 8132 3806 8134
rect 3830 8132 3886 8134
rect 3910 8132 3966 8134
rect 4710 9988 4766 10024
rect 4710 9968 4712 9988
rect 4712 9968 4764 9988
rect 4764 9968 4766 9988
rect 3670 7098 3726 7100
rect 3750 7098 3806 7100
rect 3830 7098 3886 7100
rect 3910 7098 3966 7100
rect 3670 7046 3716 7098
rect 3716 7046 3726 7098
rect 3750 7046 3780 7098
rect 3780 7046 3792 7098
rect 3792 7046 3806 7098
rect 3830 7046 3844 7098
rect 3844 7046 3856 7098
rect 3856 7046 3886 7098
rect 3910 7046 3920 7098
rect 3920 7046 3966 7098
rect 3670 7044 3726 7046
rect 3750 7044 3806 7046
rect 3830 7044 3886 7046
rect 3910 7044 3966 7046
rect 3670 6010 3726 6012
rect 3750 6010 3806 6012
rect 3830 6010 3886 6012
rect 3910 6010 3966 6012
rect 3670 5958 3716 6010
rect 3716 5958 3726 6010
rect 3750 5958 3780 6010
rect 3780 5958 3792 6010
rect 3792 5958 3806 6010
rect 3830 5958 3844 6010
rect 3844 5958 3856 6010
rect 3856 5958 3886 6010
rect 3910 5958 3920 6010
rect 3920 5958 3966 6010
rect 3670 5956 3726 5958
rect 3750 5956 3806 5958
rect 3830 5956 3886 5958
rect 3910 5956 3966 5958
rect 3670 4922 3726 4924
rect 3750 4922 3806 4924
rect 3830 4922 3886 4924
rect 3910 4922 3966 4924
rect 3670 4870 3716 4922
rect 3716 4870 3726 4922
rect 3750 4870 3780 4922
rect 3780 4870 3792 4922
rect 3792 4870 3806 4922
rect 3830 4870 3844 4922
rect 3844 4870 3856 4922
rect 3856 4870 3886 4922
rect 3910 4870 3920 4922
rect 3920 4870 3966 4922
rect 3670 4868 3726 4870
rect 3750 4868 3806 4870
rect 3830 4868 3886 4870
rect 3910 4868 3966 4870
rect 3670 3834 3726 3836
rect 3750 3834 3806 3836
rect 3830 3834 3886 3836
rect 3910 3834 3966 3836
rect 3670 3782 3716 3834
rect 3716 3782 3726 3834
rect 3750 3782 3780 3834
rect 3780 3782 3792 3834
rect 3792 3782 3806 3834
rect 3830 3782 3844 3834
rect 3844 3782 3856 3834
rect 3856 3782 3886 3834
rect 3910 3782 3920 3834
rect 3920 3782 3966 3834
rect 3670 3780 3726 3782
rect 3750 3780 3806 3782
rect 3830 3780 3886 3782
rect 3910 3780 3966 3782
rect 3670 2746 3726 2748
rect 3750 2746 3806 2748
rect 3830 2746 3886 2748
rect 3910 2746 3966 2748
rect 3670 2694 3716 2746
rect 3716 2694 3726 2746
rect 3750 2694 3780 2746
rect 3780 2694 3792 2746
rect 3792 2694 3806 2746
rect 3830 2694 3844 2746
rect 3844 2694 3856 2746
rect 3856 2694 3886 2746
rect 3910 2694 3920 2746
rect 3920 2694 3966 2746
rect 3670 2692 3726 2694
rect 3750 2692 3806 2694
rect 3830 2692 3886 2694
rect 3910 2692 3966 2694
rect 5722 12436 5778 12472
rect 5722 12416 5724 12436
rect 5724 12416 5776 12436
rect 5776 12416 5778 12436
rect 6384 16346 6440 16348
rect 6464 16346 6520 16348
rect 6544 16346 6600 16348
rect 6624 16346 6680 16348
rect 6384 16294 6430 16346
rect 6430 16294 6440 16346
rect 6464 16294 6494 16346
rect 6494 16294 6506 16346
rect 6506 16294 6520 16346
rect 6544 16294 6558 16346
rect 6558 16294 6570 16346
rect 6570 16294 6600 16346
rect 6624 16294 6634 16346
rect 6634 16294 6680 16346
rect 6384 16292 6440 16294
rect 6464 16292 6520 16294
rect 6544 16292 6600 16294
rect 6624 16292 6680 16294
rect 6384 15258 6440 15260
rect 6464 15258 6520 15260
rect 6544 15258 6600 15260
rect 6624 15258 6680 15260
rect 6384 15206 6430 15258
rect 6430 15206 6440 15258
rect 6464 15206 6494 15258
rect 6494 15206 6506 15258
rect 6506 15206 6520 15258
rect 6544 15206 6558 15258
rect 6558 15206 6570 15258
rect 6570 15206 6600 15258
rect 6624 15206 6634 15258
rect 6634 15206 6680 15258
rect 6384 15204 6440 15206
rect 6464 15204 6520 15206
rect 6544 15204 6600 15206
rect 6624 15204 6680 15206
rect 9098 19066 9154 19068
rect 9178 19066 9234 19068
rect 9258 19066 9314 19068
rect 9338 19066 9394 19068
rect 9098 19014 9144 19066
rect 9144 19014 9154 19066
rect 9178 19014 9208 19066
rect 9208 19014 9220 19066
rect 9220 19014 9234 19066
rect 9258 19014 9272 19066
rect 9272 19014 9284 19066
rect 9284 19014 9314 19066
rect 9338 19014 9348 19066
rect 9348 19014 9394 19066
rect 9098 19012 9154 19014
rect 9178 19012 9234 19014
rect 9258 19012 9314 19014
rect 9338 19012 9394 19014
rect 11812 19610 11868 19612
rect 11892 19610 11948 19612
rect 11972 19610 12028 19612
rect 12052 19610 12108 19612
rect 11812 19558 11858 19610
rect 11858 19558 11868 19610
rect 11892 19558 11922 19610
rect 11922 19558 11934 19610
rect 11934 19558 11948 19610
rect 11972 19558 11986 19610
rect 11986 19558 11998 19610
rect 11998 19558 12028 19610
rect 12052 19558 12062 19610
rect 12062 19558 12108 19610
rect 11812 19556 11868 19558
rect 11892 19556 11948 19558
rect 11972 19556 12028 19558
rect 12052 19556 12108 19558
rect 14526 20154 14582 20156
rect 14606 20154 14662 20156
rect 14686 20154 14742 20156
rect 14766 20154 14822 20156
rect 14526 20102 14572 20154
rect 14572 20102 14582 20154
rect 14606 20102 14636 20154
rect 14636 20102 14648 20154
rect 14648 20102 14662 20154
rect 14686 20102 14700 20154
rect 14700 20102 14712 20154
rect 14712 20102 14742 20154
rect 14766 20102 14776 20154
rect 14776 20102 14822 20154
rect 14526 20100 14582 20102
rect 14606 20100 14662 20102
rect 14686 20100 14742 20102
rect 14766 20100 14822 20102
rect 14526 19066 14582 19068
rect 14606 19066 14662 19068
rect 14686 19066 14742 19068
rect 14766 19066 14822 19068
rect 14526 19014 14572 19066
rect 14572 19014 14582 19066
rect 14606 19014 14636 19066
rect 14636 19014 14648 19066
rect 14648 19014 14662 19066
rect 14686 19014 14700 19066
rect 14700 19014 14712 19066
rect 14712 19014 14742 19066
rect 14766 19014 14776 19066
rect 14776 19014 14822 19066
rect 14526 19012 14582 19014
rect 14606 19012 14662 19014
rect 14686 19012 14742 19014
rect 14766 19012 14822 19014
rect 9098 17978 9154 17980
rect 9178 17978 9234 17980
rect 9258 17978 9314 17980
rect 9338 17978 9394 17980
rect 9098 17926 9144 17978
rect 9144 17926 9154 17978
rect 9178 17926 9208 17978
rect 9208 17926 9220 17978
rect 9220 17926 9234 17978
rect 9258 17926 9272 17978
rect 9272 17926 9284 17978
rect 9284 17926 9314 17978
rect 9338 17926 9348 17978
rect 9348 17926 9394 17978
rect 9098 17924 9154 17926
rect 9178 17924 9234 17926
rect 9258 17924 9314 17926
rect 9338 17924 9394 17926
rect 11812 18522 11868 18524
rect 11892 18522 11948 18524
rect 11972 18522 12028 18524
rect 12052 18522 12108 18524
rect 11812 18470 11858 18522
rect 11858 18470 11868 18522
rect 11892 18470 11922 18522
rect 11922 18470 11934 18522
rect 11934 18470 11948 18522
rect 11972 18470 11986 18522
rect 11986 18470 11998 18522
rect 11998 18470 12028 18522
rect 12052 18470 12062 18522
rect 12062 18470 12108 18522
rect 11812 18468 11868 18470
rect 11892 18468 11948 18470
rect 11972 18468 12028 18470
rect 12052 18468 12108 18470
rect 5906 12416 5962 12472
rect 6384 14170 6440 14172
rect 6464 14170 6520 14172
rect 6544 14170 6600 14172
rect 6624 14170 6680 14172
rect 6384 14118 6430 14170
rect 6430 14118 6440 14170
rect 6464 14118 6494 14170
rect 6494 14118 6506 14170
rect 6506 14118 6520 14170
rect 6544 14118 6558 14170
rect 6558 14118 6570 14170
rect 6570 14118 6600 14170
rect 6624 14118 6634 14170
rect 6634 14118 6680 14170
rect 6384 14116 6440 14118
rect 6464 14116 6520 14118
rect 6544 14116 6600 14118
rect 6624 14116 6680 14118
rect 6384 13082 6440 13084
rect 6464 13082 6520 13084
rect 6544 13082 6600 13084
rect 6624 13082 6680 13084
rect 6384 13030 6430 13082
rect 6430 13030 6440 13082
rect 6464 13030 6494 13082
rect 6494 13030 6506 13082
rect 6506 13030 6520 13082
rect 6544 13030 6558 13082
rect 6558 13030 6570 13082
rect 6570 13030 6600 13082
rect 6624 13030 6634 13082
rect 6634 13030 6680 13082
rect 6384 13028 6440 13030
rect 6464 13028 6520 13030
rect 6544 13028 6600 13030
rect 6624 13028 6680 13030
rect 5906 10512 5962 10568
rect 6384 11994 6440 11996
rect 6464 11994 6520 11996
rect 6544 11994 6600 11996
rect 6624 11994 6680 11996
rect 6384 11942 6430 11994
rect 6430 11942 6440 11994
rect 6464 11942 6494 11994
rect 6494 11942 6506 11994
rect 6506 11942 6520 11994
rect 6544 11942 6558 11994
rect 6558 11942 6570 11994
rect 6570 11942 6600 11994
rect 6624 11942 6634 11994
rect 6634 11942 6680 11994
rect 6384 11940 6440 11942
rect 6464 11940 6520 11942
rect 6544 11940 6600 11942
rect 6624 11940 6680 11942
rect 6384 10906 6440 10908
rect 6464 10906 6520 10908
rect 6544 10906 6600 10908
rect 6624 10906 6680 10908
rect 6384 10854 6430 10906
rect 6430 10854 6440 10906
rect 6464 10854 6494 10906
rect 6494 10854 6506 10906
rect 6506 10854 6520 10906
rect 6544 10854 6558 10906
rect 6558 10854 6570 10906
rect 6570 10854 6600 10906
rect 6624 10854 6634 10906
rect 6634 10854 6680 10906
rect 6384 10852 6440 10854
rect 6464 10852 6520 10854
rect 6544 10852 6600 10854
rect 6624 10852 6680 10854
rect 6274 10512 6330 10568
rect 6384 9818 6440 9820
rect 6464 9818 6520 9820
rect 6544 9818 6600 9820
rect 6624 9818 6680 9820
rect 6384 9766 6430 9818
rect 6430 9766 6440 9818
rect 6464 9766 6494 9818
rect 6494 9766 6506 9818
rect 6506 9766 6520 9818
rect 6544 9766 6558 9818
rect 6558 9766 6570 9818
rect 6570 9766 6600 9818
rect 6624 9766 6634 9818
rect 6634 9766 6680 9818
rect 6384 9764 6440 9766
rect 6464 9764 6520 9766
rect 6544 9764 6600 9766
rect 6624 9764 6680 9766
rect 6384 8730 6440 8732
rect 6464 8730 6520 8732
rect 6544 8730 6600 8732
rect 6624 8730 6680 8732
rect 6384 8678 6430 8730
rect 6430 8678 6440 8730
rect 6464 8678 6494 8730
rect 6494 8678 6506 8730
rect 6506 8678 6520 8730
rect 6544 8678 6558 8730
rect 6558 8678 6570 8730
rect 6570 8678 6600 8730
rect 6624 8678 6634 8730
rect 6634 8678 6680 8730
rect 6384 8676 6440 8678
rect 6464 8676 6520 8678
rect 6544 8676 6600 8678
rect 6624 8676 6680 8678
rect 6384 7642 6440 7644
rect 6464 7642 6520 7644
rect 6544 7642 6600 7644
rect 6624 7642 6680 7644
rect 6384 7590 6430 7642
rect 6430 7590 6440 7642
rect 6464 7590 6494 7642
rect 6494 7590 6506 7642
rect 6506 7590 6520 7642
rect 6544 7590 6558 7642
rect 6558 7590 6570 7642
rect 6570 7590 6600 7642
rect 6624 7590 6634 7642
rect 6634 7590 6680 7642
rect 6384 7588 6440 7590
rect 6464 7588 6520 7590
rect 6544 7588 6600 7590
rect 6624 7588 6680 7590
rect 7010 7928 7066 7984
rect 6384 6554 6440 6556
rect 6464 6554 6520 6556
rect 6544 6554 6600 6556
rect 6624 6554 6680 6556
rect 6384 6502 6430 6554
rect 6430 6502 6440 6554
rect 6464 6502 6494 6554
rect 6494 6502 6506 6554
rect 6506 6502 6520 6554
rect 6544 6502 6558 6554
rect 6558 6502 6570 6554
rect 6570 6502 6600 6554
rect 6624 6502 6634 6554
rect 6634 6502 6680 6554
rect 6384 6500 6440 6502
rect 6464 6500 6520 6502
rect 6544 6500 6600 6502
rect 6624 6500 6680 6502
rect 6384 5466 6440 5468
rect 6464 5466 6520 5468
rect 6544 5466 6600 5468
rect 6624 5466 6680 5468
rect 6384 5414 6430 5466
rect 6430 5414 6440 5466
rect 6464 5414 6494 5466
rect 6494 5414 6506 5466
rect 6506 5414 6520 5466
rect 6544 5414 6558 5466
rect 6558 5414 6570 5466
rect 6570 5414 6600 5466
rect 6624 5414 6634 5466
rect 6634 5414 6680 5466
rect 6384 5412 6440 5414
rect 6464 5412 6520 5414
rect 6544 5412 6600 5414
rect 6624 5412 6680 5414
rect 6384 4378 6440 4380
rect 6464 4378 6520 4380
rect 6544 4378 6600 4380
rect 6624 4378 6680 4380
rect 6384 4326 6430 4378
rect 6430 4326 6440 4378
rect 6464 4326 6494 4378
rect 6494 4326 6506 4378
rect 6506 4326 6520 4378
rect 6544 4326 6558 4378
rect 6558 4326 6570 4378
rect 6570 4326 6600 4378
rect 6624 4326 6634 4378
rect 6634 4326 6680 4378
rect 6384 4324 6440 4326
rect 6464 4324 6520 4326
rect 6544 4324 6600 4326
rect 6624 4324 6680 4326
rect 6384 3290 6440 3292
rect 6464 3290 6520 3292
rect 6544 3290 6600 3292
rect 6624 3290 6680 3292
rect 6384 3238 6430 3290
rect 6430 3238 6440 3290
rect 6464 3238 6494 3290
rect 6494 3238 6506 3290
rect 6506 3238 6520 3290
rect 6544 3238 6558 3290
rect 6558 3238 6570 3290
rect 6570 3238 6600 3290
rect 6624 3238 6634 3290
rect 6634 3238 6680 3290
rect 6384 3236 6440 3238
rect 6464 3236 6520 3238
rect 6544 3236 6600 3238
rect 6624 3236 6680 3238
rect 9098 16890 9154 16892
rect 9178 16890 9234 16892
rect 9258 16890 9314 16892
rect 9338 16890 9394 16892
rect 9098 16838 9144 16890
rect 9144 16838 9154 16890
rect 9178 16838 9208 16890
rect 9208 16838 9220 16890
rect 9220 16838 9234 16890
rect 9258 16838 9272 16890
rect 9272 16838 9284 16890
rect 9284 16838 9314 16890
rect 9338 16838 9348 16890
rect 9348 16838 9394 16890
rect 9098 16836 9154 16838
rect 9178 16836 9234 16838
rect 9258 16836 9314 16838
rect 9338 16836 9394 16838
rect 11812 17434 11868 17436
rect 11892 17434 11948 17436
rect 11972 17434 12028 17436
rect 12052 17434 12108 17436
rect 11812 17382 11858 17434
rect 11858 17382 11868 17434
rect 11892 17382 11922 17434
rect 11922 17382 11934 17434
rect 11934 17382 11948 17434
rect 11972 17382 11986 17434
rect 11986 17382 11998 17434
rect 11998 17382 12028 17434
rect 12052 17382 12062 17434
rect 12062 17382 12108 17434
rect 11812 17380 11868 17382
rect 11892 17380 11948 17382
rect 11972 17380 12028 17382
rect 12052 17380 12108 17382
rect 11812 16346 11868 16348
rect 11892 16346 11948 16348
rect 11972 16346 12028 16348
rect 12052 16346 12108 16348
rect 11812 16294 11858 16346
rect 11858 16294 11868 16346
rect 11892 16294 11922 16346
rect 11922 16294 11934 16346
rect 11934 16294 11948 16346
rect 11972 16294 11986 16346
rect 11986 16294 11998 16346
rect 11998 16294 12028 16346
rect 12052 16294 12062 16346
rect 12062 16294 12108 16346
rect 11812 16292 11868 16294
rect 11892 16292 11948 16294
rect 11972 16292 12028 16294
rect 12052 16292 12108 16294
rect 9098 15802 9154 15804
rect 9178 15802 9234 15804
rect 9258 15802 9314 15804
rect 9338 15802 9394 15804
rect 9098 15750 9144 15802
rect 9144 15750 9154 15802
rect 9178 15750 9208 15802
rect 9208 15750 9220 15802
rect 9220 15750 9234 15802
rect 9258 15750 9272 15802
rect 9272 15750 9284 15802
rect 9284 15750 9314 15802
rect 9338 15750 9348 15802
rect 9348 15750 9394 15802
rect 9098 15748 9154 15750
rect 9178 15748 9234 15750
rect 9258 15748 9314 15750
rect 9338 15748 9394 15750
rect 9098 14714 9154 14716
rect 9178 14714 9234 14716
rect 9258 14714 9314 14716
rect 9338 14714 9394 14716
rect 9098 14662 9144 14714
rect 9144 14662 9154 14714
rect 9178 14662 9208 14714
rect 9208 14662 9220 14714
rect 9220 14662 9234 14714
rect 9258 14662 9272 14714
rect 9272 14662 9284 14714
rect 9284 14662 9314 14714
rect 9338 14662 9348 14714
rect 9348 14662 9394 14714
rect 9098 14660 9154 14662
rect 9178 14660 9234 14662
rect 9258 14660 9314 14662
rect 9338 14660 9394 14662
rect 9098 13626 9154 13628
rect 9178 13626 9234 13628
rect 9258 13626 9314 13628
rect 9338 13626 9394 13628
rect 9098 13574 9144 13626
rect 9144 13574 9154 13626
rect 9178 13574 9208 13626
rect 9208 13574 9220 13626
rect 9220 13574 9234 13626
rect 9258 13574 9272 13626
rect 9272 13574 9284 13626
rect 9284 13574 9314 13626
rect 9338 13574 9348 13626
rect 9348 13574 9394 13626
rect 9098 13572 9154 13574
rect 9178 13572 9234 13574
rect 9258 13572 9314 13574
rect 9338 13572 9394 13574
rect 9098 12538 9154 12540
rect 9178 12538 9234 12540
rect 9258 12538 9314 12540
rect 9338 12538 9394 12540
rect 9098 12486 9144 12538
rect 9144 12486 9154 12538
rect 9178 12486 9208 12538
rect 9208 12486 9220 12538
rect 9220 12486 9234 12538
rect 9258 12486 9272 12538
rect 9272 12486 9284 12538
rect 9284 12486 9314 12538
rect 9338 12486 9348 12538
rect 9348 12486 9394 12538
rect 9098 12484 9154 12486
rect 9178 12484 9234 12486
rect 9258 12484 9314 12486
rect 9338 12484 9394 12486
rect 9098 11450 9154 11452
rect 9178 11450 9234 11452
rect 9258 11450 9314 11452
rect 9338 11450 9394 11452
rect 9098 11398 9144 11450
rect 9144 11398 9154 11450
rect 9178 11398 9208 11450
rect 9208 11398 9220 11450
rect 9220 11398 9234 11450
rect 9258 11398 9272 11450
rect 9272 11398 9284 11450
rect 9284 11398 9314 11450
rect 9338 11398 9348 11450
rect 9348 11398 9394 11450
rect 9098 11396 9154 11398
rect 9178 11396 9234 11398
rect 9258 11396 9314 11398
rect 9338 11396 9394 11398
rect 9678 10684 9680 10704
rect 9680 10684 9732 10704
rect 9732 10684 9734 10704
rect 9678 10648 9734 10684
rect 9098 10362 9154 10364
rect 9178 10362 9234 10364
rect 9258 10362 9314 10364
rect 9338 10362 9394 10364
rect 9098 10310 9144 10362
rect 9144 10310 9154 10362
rect 9178 10310 9208 10362
rect 9208 10310 9220 10362
rect 9220 10310 9234 10362
rect 9258 10310 9272 10362
rect 9272 10310 9284 10362
rect 9284 10310 9314 10362
rect 9338 10310 9348 10362
rect 9348 10310 9394 10362
rect 9098 10308 9154 10310
rect 9178 10308 9234 10310
rect 9258 10308 9314 10310
rect 9338 10308 9394 10310
rect 9098 9274 9154 9276
rect 9178 9274 9234 9276
rect 9258 9274 9314 9276
rect 9338 9274 9394 9276
rect 9098 9222 9144 9274
rect 9144 9222 9154 9274
rect 9178 9222 9208 9274
rect 9208 9222 9220 9274
rect 9220 9222 9234 9274
rect 9258 9222 9272 9274
rect 9272 9222 9284 9274
rect 9284 9222 9314 9274
rect 9338 9222 9348 9274
rect 9348 9222 9394 9274
rect 9098 9220 9154 9222
rect 9178 9220 9234 9222
rect 9258 9220 9314 9222
rect 9338 9220 9394 9222
rect 9098 8186 9154 8188
rect 9178 8186 9234 8188
rect 9258 8186 9314 8188
rect 9338 8186 9394 8188
rect 9098 8134 9144 8186
rect 9144 8134 9154 8186
rect 9178 8134 9208 8186
rect 9208 8134 9220 8186
rect 9220 8134 9234 8186
rect 9258 8134 9272 8186
rect 9272 8134 9284 8186
rect 9284 8134 9314 8186
rect 9338 8134 9348 8186
rect 9348 8134 9394 8186
rect 9098 8132 9154 8134
rect 9178 8132 9234 8134
rect 9258 8132 9314 8134
rect 9338 8132 9394 8134
rect 9098 7098 9154 7100
rect 9178 7098 9234 7100
rect 9258 7098 9314 7100
rect 9338 7098 9394 7100
rect 9098 7046 9144 7098
rect 9144 7046 9154 7098
rect 9178 7046 9208 7098
rect 9208 7046 9220 7098
rect 9220 7046 9234 7098
rect 9258 7046 9272 7098
rect 9272 7046 9284 7098
rect 9284 7046 9314 7098
rect 9338 7046 9348 7098
rect 9348 7046 9394 7098
rect 9098 7044 9154 7046
rect 9178 7044 9234 7046
rect 9258 7044 9314 7046
rect 9338 7044 9394 7046
rect 9098 6010 9154 6012
rect 9178 6010 9234 6012
rect 9258 6010 9314 6012
rect 9338 6010 9394 6012
rect 9098 5958 9144 6010
rect 9144 5958 9154 6010
rect 9178 5958 9208 6010
rect 9208 5958 9220 6010
rect 9220 5958 9234 6010
rect 9258 5958 9272 6010
rect 9272 5958 9284 6010
rect 9284 5958 9314 6010
rect 9338 5958 9348 6010
rect 9348 5958 9394 6010
rect 9098 5956 9154 5958
rect 9178 5956 9234 5958
rect 9258 5956 9314 5958
rect 9338 5956 9394 5958
rect 9098 4922 9154 4924
rect 9178 4922 9234 4924
rect 9258 4922 9314 4924
rect 9338 4922 9394 4924
rect 9098 4870 9144 4922
rect 9144 4870 9154 4922
rect 9178 4870 9208 4922
rect 9208 4870 9220 4922
rect 9220 4870 9234 4922
rect 9258 4870 9272 4922
rect 9272 4870 9284 4922
rect 9284 4870 9314 4922
rect 9338 4870 9348 4922
rect 9348 4870 9394 4922
rect 9098 4868 9154 4870
rect 9178 4868 9234 4870
rect 9258 4868 9314 4870
rect 9338 4868 9394 4870
rect 9098 3834 9154 3836
rect 9178 3834 9234 3836
rect 9258 3834 9314 3836
rect 9338 3834 9394 3836
rect 9098 3782 9144 3834
rect 9144 3782 9154 3834
rect 9178 3782 9208 3834
rect 9208 3782 9220 3834
rect 9220 3782 9234 3834
rect 9258 3782 9272 3834
rect 9272 3782 9284 3834
rect 9284 3782 9314 3834
rect 9338 3782 9348 3834
rect 9348 3782 9394 3834
rect 9098 3780 9154 3782
rect 9178 3780 9234 3782
rect 9258 3780 9314 3782
rect 9338 3780 9394 3782
rect 9098 2746 9154 2748
rect 9178 2746 9234 2748
rect 9258 2746 9314 2748
rect 9338 2746 9394 2748
rect 9098 2694 9144 2746
rect 9144 2694 9154 2746
rect 9178 2694 9208 2746
rect 9208 2694 9220 2746
rect 9220 2694 9234 2746
rect 9258 2694 9272 2746
rect 9272 2694 9284 2746
rect 9284 2694 9314 2746
rect 9338 2694 9348 2746
rect 9348 2694 9394 2746
rect 9098 2692 9154 2694
rect 9178 2692 9234 2694
rect 9258 2692 9314 2694
rect 9338 2692 9394 2694
rect 11812 15258 11868 15260
rect 11892 15258 11948 15260
rect 11972 15258 12028 15260
rect 12052 15258 12108 15260
rect 11812 15206 11858 15258
rect 11858 15206 11868 15258
rect 11892 15206 11922 15258
rect 11922 15206 11934 15258
rect 11934 15206 11948 15258
rect 11972 15206 11986 15258
rect 11986 15206 11998 15258
rect 11998 15206 12028 15258
rect 12052 15206 12062 15258
rect 12062 15206 12108 15258
rect 11812 15204 11868 15206
rect 11892 15204 11948 15206
rect 11972 15204 12028 15206
rect 12052 15204 12108 15206
rect 14526 17978 14582 17980
rect 14606 17978 14662 17980
rect 14686 17978 14742 17980
rect 14766 17978 14822 17980
rect 14526 17926 14572 17978
rect 14572 17926 14582 17978
rect 14606 17926 14636 17978
rect 14636 17926 14648 17978
rect 14648 17926 14662 17978
rect 14686 17926 14700 17978
rect 14700 17926 14712 17978
rect 14712 17926 14742 17978
rect 14766 17926 14776 17978
rect 14776 17926 14822 17978
rect 14526 17924 14582 17926
rect 14606 17924 14662 17926
rect 14686 17924 14742 17926
rect 14766 17924 14822 17926
rect 14526 16890 14582 16892
rect 14606 16890 14662 16892
rect 14686 16890 14742 16892
rect 14766 16890 14822 16892
rect 14526 16838 14572 16890
rect 14572 16838 14582 16890
rect 14606 16838 14636 16890
rect 14636 16838 14648 16890
rect 14648 16838 14662 16890
rect 14686 16838 14700 16890
rect 14700 16838 14712 16890
rect 14712 16838 14742 16890
rect 14766 16838 14776 16890
rect 14776 16838 14822 16890
rect 14526 16836 14582 16838
rect 14606 16836 14662 16838
rect 14686 16836 14742 16838
rect 14766 16836 14822 16838
rect 14526 15802 14582 15804
rect 14606 15802 14662 15804
rect 14686 15802 14742 15804
rect 14766 15802 14822 15804
rect 14526 15750 14572 15802
rect 14572 15750 14582 15802
rect 14606 15750 14636 15802
rect 14636 15750 14648 15802
rect 14648 15750 14662 15802
rect 14686 15750 14700 15802
rect 14700 15750 14712 15802
rect 14712 15750 14742 15802
rect 14766 15750 14776 15802
rect 14776 15750 14822 15802
rect 14526 15748 14582 15750
rect 14606 15748 14662 15750
rect 14686 15748 14742 15750
rect 14766 15748 14822 15750
rect 11812 14170 11868 14172
rect 11892 14170 11948 14172
rect 11972 14170 12028 14172
rect 12052 14170 12108 14172
rect 11812 14118 11858 14170
rect 11858 14118 11868 14170
rect 11892 14118 11922 14170
rect 11922 14118 11934 14170
rect 11934 14118 11948 14170
rect 11972 14118 11986 14170
rect 11986 14118 11998 14170
rect 11998 14118 12028 14170
rect 12052 14118 12062 14170
rect 12062 14118 12108 14170
rect 11812 14116 11868 14118
rect 11892 14116 11948 14118
rect 11972 14116 12028 14118
rect 12052 14116 12108 14118
rect 11812 13082 11868 13084
rect 11892 13082 11948 13084
rect 11972 13082 12028 13084
rect 12052 13082 12108 13084
rect 11812 13030 11858 13082
rect 11858 13030 11868 13082
rect 11892 13030 11922 13082
rect 11922 13030 11934 13082
rect 11934 13030 11948 13082
rect 11972 13030 11986 13082
rect 11986 13030 11998 13082
rect 11998 13030 12028 13082
rect 12052 13030 12062 13082
rect 12062 13030 12108 13082
rect 11812 13028 11868 13030
rect 11892 13028 11948 13030
rect 11972 13028 12028 13030
rect 12052 13028 12108 13030
rect 11812 11994 11868 11996
rect 11892 11994 11948 11996
rect 11972 11994 12028 11996
rect 12052 11994 12108 11996
rect 11812 11942 11858 11994
rect 11858 11942 11868 11994
rect 11892 11942 11922 11994
rect 11922 11942 11934 11994
rect 11934 11942 11948 11994
rect 11972 11942 11986 11994
rect 11986 11942 11998 11994
rect 11998 11942 12028 11994
rect 12052 11942 12062 11994
rect 12062 11942 12108 11994
rect 11812 11940 11868 11942
rect 11892 11940 11948 11942
rect 11972 11940 12028 11942
rect 12052 11940 12108 11942
rect 11812 10906 11868 10908
rect 11892 10906 11948 10908
rect 11972 10906 12028 10908
rect 12052 10906 12108 10908
rect 11812 10854 11858 10906
rect 11858 10854 11868 10906
rect 11892 10854 11922 10906
rect 11922 10854 11934 10906
rect 11934 10854 11948 10906
rect 11972 10854 11986 10906
rect 11986 10854 11998 10906
rect 11998 10854 12028 10906
rect 12052 10854 12062 10906
rect 12062 10854 12108 10906
rect 11812 10852 11868 10854
rect 11892 10852 11948 10854
rect 11972 10852 12028 10854
rect 12052 10852 12108 10854
rect 11812 9818 11868 9820
rect 11892 9818 11948 9820
rect 11972 9818 12028 9820
rect 12052 9818 12108 9820
rect 11812 9766 11858 9818
rect 11858 9766 11868 9818
rect 11892 9766 11922 9818
rect 11922 9766 11934 9818
rect 11934 9766 11948 9818
rect 11972 9766 11986 9818
rect 11986 9766 11998 9818
rect 11998 9766 12028 9818
rect 12052 9766 12062 9818
rect 12062 9766 12108 9818
rect 11812 9764 11868 9766
rect 11892 9764 11948 9766
rect 11972 9764 12028 9766
rect 12052 9764 12108 9766
rect 11812 8730 11868 8732
rect 11892 8730 11948 8732
rect 11972 8730 12028 8732
rect 12052 8730 12108 8732
rect 11812 8678 11858 8730
rect 11858 8678 11868 8730
rect 11892 8678 11922 8730
rect 11922 8678 11934 8730
rect 11934 8678 11948 8730
rect 11972 8678 11986 8730
rect 11986 8678 11998 8730
rect 11998 8678 12028 8730
rect 12052 8678 12062 8730
rect 12062 8678 12108 8730
rect 11812 8676 11868 8678
rect 11892 8676 11948 8678
rect 11972 8676 12028 8678
rect 12052 8676 12108 8678
rect 11812 7642 11868 7644
rect 11892 7642 11948 7644
rect 11972 7642 12028 7644
rect 12052 7642 12108 7644
rect 11812 7590 11858 7642
rect 11858 7590 11868 7642
rect 11892 7590 11922 7642
rect 11922 7590 11934 7642
rect 11934 7590 11948 7642
rect 11972 7590 11986 7642
rect 11986 7590 11998 7642
rect 11998 7590 12028 7642
rect 12052 7590 12062 7642
rect 12062 7590 12108 7642
rect 11812 7588 11868 7590
rect 11892 7588 11948 7590
rect 11972 7588 12028 7590
rect 12052 7588 12108 7590
rect 14526 14714 14582 14716
rect 14606 14714 14662 14716
rect 14686 14714 14742 14716
rect 14766 14714 14822 14716
rect 14526 14662 14572 14714
rect 14572 14662 14582 14714
rect 14606 14662 14636 14714
rect 14636 14662 14648 14714
rect 14648 14662 14662 14714
rect 14686 14662 14700 14714
rect 14700 14662 14712 14714
rect 14712 14662 14742 14714
rect 14766 14662 14776 14714
rect 14776 14662 14822 14714
rect 14526 14660 14582 14662
rect 14606 14660 14662 14662
rect 14686 14660 14742 14662
rect 14766 14660 14822 14662
rect 14526 13626 14582 13628
rect 14606 13626 14662 13628
rect 14686 13626 14742 13628
rect 14766 13626 14822 13628
rect 14526 13574 14572 13626
rect 14572 13574 14582 13626
rect 14606 13574 14636 13626
rect 14636 13574 14648 13626
rect 14648 13574 14662 13626
rect 14686 13574 14700 13626
rect 14700 13574 14712 13626
rect 14712 13574 14742 13626
rect 14766 13574 14776 13626
rect 14776 13574 14822 13626
rect 14526 13572 14582 13574
rect 14606 13572 14662 13574
rect 14686 13572 14742 13574
rect 14766 13572 14822 13574
rect 14526 12538 14582 12540
rect 14606 12538 14662 12540
rect 14686 12538 14742 12540
rect 14766 12538 14822 12540
rect 14526 12486 14572 12538
rect 14572 12486 14582 12538
rect 14606 12486 14636 12538
rect 14636 12486 14648 12538
rect 14648 12486 14662 12538
rect 14686 12486 14700 12538
rect 14700 12486 14712 12538
rect 14712 12486 14742 12538
rect 14766 12486 14776 12538
rect 14776 12486 14822 12538
rect 14526 12484 14582 12486
rect 14606 12484 14662 12486
rect 14686 12484 14742 12486
rect 14766 12484 14822 12486
rect 14526 11450 14582 11452
rect 14606 11450 14662 11452
rect 14686 11450 14742 11452
rect 14766 11450 14822 11452
rect 14526 11398 14572 11450
rect 14572 11398 14582 11450
rect 14606 11398 14636 11450
rect 14636 11398 14648 11450
rect 14648 11398 14662 11450
rect 14686 11398 14700 11450
rect 14700 11398 14712 11450
rect 14712 11398 14742 11450
rect 14766 11398 14776 11450
rect 14776 11398 14822 11450
rect 14526 11396 14582 11398
rect 14606 11396 14662 11398
rect 14686 11396 14742 11398
rect 14766 11396 14822 11398
rect 14526 10362 14582 10364
rect 14606 10362 14662 10364
rect 14686 10362 14742 10364
rect 14766 10362 14822 10364
rect 14526 10310 14572 10362
rect 14572 10310 14582 10362
rect 14606 10310 14636 10362
rect 14636 10310 14648 10362
rect 14648 10310 14662 10362
rect 14686 10310 14700 10362
rect 14700 10310 14712 10362
rect 14712 10310 14742 10362
rect 14766 10310 14776 10362
rect 14776 10310 14822 10362
rect 14526 10308 14582 10310
rect 14606 10308 14662 10310
rect 14686 10308 14742 10310
rect 14766 10308 14822 10310
rect 14526 9274 14582 9276
rect 14606 9274 14662 9276
rect 14686 9274 14742 9276
rect 14766 9274 14822 9276
rect 14526 9222 14572 9274
rect 14572 9222 14582 9274
rect 14606 9222 14636 9274
rect 14636 9222 14648 9274
rect 14648 9222 14662 9274
rect 14686 9222 14700 9274
rect 14700 9222 14712 9274
rect 14712 9222 14742 9274
rect 14766 9222 14776 9274
rect 14776 9222 14822 9274
rect 14526 9220 14582 9222
rect 14606 9220 14662 9222
rect 14686 9220 14742 9222
rect 14766 9220 14822 9222
rect 14526 8186 14582 8188
rect 14606 8186 14662 8188
rect 14686 8186 14742 8188
rect 14766 8186 14822 8188
rect 14526 8134 14572 8186
rect 14572 8134 14582 8186
rect 14606 8134 14636 8186
rect 14636 8134 14648 8186
rect 14648 8134 14662 8186
rect 14686 8134 14700 8186
rect 14700 8134 14712 8186
rect 14712 8134 14742 8186
rect 14766 8134 14776 8186
rect 14776 8134 14822 8186
rect 14526 8132 14582 8134
rect 14606 8132 14662 8134
rect 14686 8132 14742 8134
rect 14766 8132 14822 8134
rect 16302 20984 16358 21040
rect 17314 21020 17316 21040
rect 17316 21020 17368 21040
rect 17368 21020 17370 21040
rect 17314 20984 17370 21020
rect 17240 20698 17296 20700
rect 17320 20698 17376 20700
rect 17400 20698 17456 20700
rect 17480 20698 17536 20700
rect 17240 20646 17286 20698
rect 17286 20646 17296 20698
rect 17320 20646 17350 20698
rect 17350 20646 17362 20698
rect 17362 20646 17376 20698
rect 17400 20646 17414 20698
rect 17414 20646 17426 20698
rect 17426 20646 17456 20698
rect 17480 20646 17490 20698
rect 17490 20646 17536 20698
rect 17240 20644 17296 20646
rect 17320 20644 17376 20646
rect 17400 20644 17456 20646
rect 17480 20644 17536 20646
rect 17240 19610 17296 19612
rect 17320 19610 17376 19612
rect 17400 19610 17456 19612
rect 17480 19610 17536 19612
rect 17240 19558 17286 19610
rect 17286 19558 17296 19610
rect 17320 19558 17350 19610
rect 17350 19558 17362 19610
rect 17362 19558 17376 19610
rect 17400 19558 17414 19610
rect 17414 19558 17426 19610
rect 17426 19558 17456 19610
rect 17480 19558 17490 19610
rect 17490 19558 17536 19610
rect 17240 19556 17296 19558
rect 17320 19556 17376 19558
rect 17400 19556 17456 19558
rect 17480 19556 17536 19558
rect 17240 18522 17296 18524
rect 17320 18522 17376 18524
rect 17400 18522 17456 18524
rect 17480 18522 17536 18524
rect 17240 18470 17286 18522
rect 17286 18470 17296 18522
rect 17320 18470 17350 18522
rect 17350 18470 17362 18522
rect 17362 18470 17376 18522
rect 17400 18470 17414 18522
rect 17414 18470 17426 18522
rect 17426 18470 17456 18522
rect 17480 18470 17490 18522
rect 17490 18470 17536 18522
rect 17240 18468 17296 18470
rect 17320 18468 17376 18470
rect 17400 18468 17456 18470
rect 17480 18468 17536 18470
rect 19954 21242 20010 21244
rect 20034 21242 20090 21244
rect 20114 21242 20170 21244
rect 20194 21242 20250 21244
rect 19954 21190 20000 21242
rect 20000 21190 20010 21242
rect 20034 21190 20064 21242
rect 20064 21190 20076 21242
rect 20076 21190 20090 21242
rect 20114 21190 20128 21242
rect 20128 21190 20140 21242
rect 20140 21190 20170 21242
rect 20194 21190 20204 21242
rect 20204 21190 20250 21242
rect 19954 21188 20010 21190
rect 20034 21188 20090 21190
rect 20114 21188 20170 21190
rect 20194 21188 20250 21190
rect 19954 20154 20010 20156
rect 20034 20154 20090 20156
rect 20114 20154 20170 20156
rect 20194 20154 20250 20156
rect 19954 20102 20000 20154
rect 20000 20102 20010 20154
rect 20034 20102 20064 20154
rect 20064 20102 20076 20154
rect 20076 20102 20090 20154
rect 20114 20102 20128 20154
rect 20128 20102 20140 20154
rect 20140 20102 20170 20154
rect 20194 20102 20204 20154
rect 20204 20102 20250 20154
rect 19954 20100 20010 20102
rect 20034 20100 20090 20102
rect 20114 20100 20170 20102
rect 20194 20100 20250 20102
rect 17240 17434 17296 17436
rect 17320 17434 17376 17436
rect 17400 17434 17456 17436
rect 17480 17434 17536 17436
rect 17240 17382 17286 17434
rect 17286 17382 17296 17434
rect 17320 17382 17350 17434
rect 17350 17382 17362 17434
rect 17362 17382 17376 17434
rect 17400 17382 17414 17434
rect 17414 17382 17426 17434
rect 17426 17382 17456 17434
rect 17480 17382 17490 17434
rect 17490 17382 17536 17434
rect 17240 17380 17296 17382
rect 17320 17380 17376 17382
rect 17400 17380 17456 17382
rect 17480 17380 17536 17382
rect 19954 19066 20010 19068
rect 20034 19066 20090 19068
rect 20114 19066 20170 19068
rect 20194 19066 20250 19068
rect 19954 19014 20000 19066
rect 20000 19014 20010 19066
rect 20034 19014 20064 19066
rect 20064 19014 20076 19066
rect 20076 19014 20090 19066
rect 20114 19014 20128 19066
rect 20128 19014 20140 19066
rect 20140 19014 20170 19066
rect 20194 19014 20204 19066
rect 20204 19014 20250 19066
rect 19954 19012 20010 19014
rect 20034 19012 20090 19014
rect 20114 19012 20170 19014
rect 20194 19012 20250 19014
rect 17240 16346 17296 16348
rect 17320 16346 17376 16348
rect 17400 16346 17456 16348
rect 17480 16346 17536 16348
rect 17240 16294 17286 16346
rect 17286 16294 17296 16346
rect 17320 16294 17350 16346
rect 17350 16294 17362 16346
rect 17362 16294 17376 16346
rect 17400 16294 17414 16346
rect 17414 16294 17426 16346
rect 17426 16294 17456 16346
rect 17480 16294 17490 16346
rect 17490 16294 17536 16346
rect 17240 16292 17296 16294
rect 17320 16292 17376 16294
rect 17400 16292 17456 16294
rect 17480 16292 17536 16294
rect 17240 15258 17296 15260
rect 17320 15258 17376 15260
rect 17400 15258 17456 15260
rect 17480 15258 17536 15260
rect 17240 15206 17286 15258
rect 17286 15206 17296 15258
rect 17320 15206 17350 15258
rect 17350 15206 17362 15258
rect 17362 15206 17376 15258
rect 17400 15206 17414 15258
rect 17414 15206 17426 15258
rect 17426 15206 17456 15258
rect 17480 15206 17490 15258
rect 17490 15206 17536 15258
rect 17240 15204 17296 15206
rect 17320 15204 17376 15206
rect 17400 15204 17456 15206
rect 17480 15204 17536 15206
rect 17240 14170 17296 14172
rect 17320 14170 17376 14172
rect 17400 14170 17456 14172
rect 17480 14170 17536 14172
rect 17240 14118 17286 14170
rect 17286 14118 17296 14170
rect 17320 14118 17350 14170
rect 17350 14118 17362 14170
rect 17362 14118 17376 14170
rect 17400 14118 17414 14170
rect 17414 14118 17426 14170
rect 17426 14118 17456 14170
rect 17480 14118 17490 14170
rect 17490 14118 17536 14170
rect 17240 14116 17296 14118
rect 17320 14116 17376 14118
rect 17400 14116 17456 14118
rect 17480 14116 17536 14118
rect 17240 13082 17296 13084
rect 17320 13082 17376 13084
rect 17400 13082 17456 13084
rect 17480 13082 17536 13084
rect 17240 13030 17286 13082
rect 17286 13030 17296 13082
rect 17320 13030 17350 13082
rect 17350 13030 17362 13082
rect 17362 13030 17376 13082
rect 17400 13030 17414 13082
rect 17414 13030 17426 13082
rect 17426 13030 17456 13082
rect 17480 13030 17490 13082
rect 17490 13030 17536 13082
rect 17240 13028 17296 13030
rect 17320 13028 17376 13030
rect 17400 13028 17456 13030
rect 17480 13028 17536 13030
rect 17240 11994 17296 11996
rect 17320 11994 17376 11996
rect 17400 11994 17456 11996
rect 17480 11994 17536 11996
rect 17240 11942 17286 11994
rect 17286 11942 17296 11994
rect 17320 11942 17350 11994
rect 17350 11942 17362 11994
rect 17362 11942 17376 11994
rect 17400 11942 17414 11994
rect 17414 11942 17426 11994
rect 17426 11942 17456 11994
rect 17480 11942 17490 11994
rect 17490 11942 17536 11994
rect 17240 11940 17296 11942
rect 17320 11940 17376 11942
rect 17400 11940 17456 11942
rect 17480 11940 17536 11942
rect 17240 10906 17296 10908
rect 17320 10906 17376 10908
rect 17400 10906 17456 10908
rect 17480 10906 17536 10908
rect 17240 10854 17286 10906
rect 17286 10854 17296 10906
rect 17320 10854 17350 10906
rect 17350 10854 17362 10906
rect 17362 10854 17376 10906
rect 17400 10854 17414 10906
rect 17414 10854 17426 10906
rect 17426 10854 17456 10906
rect 17480 10854 17490 10906
rect 17490 10854 17536 10906
rect 17240 10852 17296 10854
rect 17320 10852 17376 10854
rect 17400 10852 17456 10854
rect 17480 10852 17536 10854
rect 17240 9818 17296 9820
rect 17320 9818 17376 9820
rect 17400 9818 17456 9820
rect 17480 9818 17536 9820
rect 17240 9766 17286 9818
rect 17286 9766 17296 9818
rect 17320 9766 17350 9818
rect 17350 9766 17362 9818
rect 17362 9766 17376 9818
rect 17400 9766 17414 9818
rect 17414 9766 17426 9818
rect 17426 9766 17456 9818
rect 17480 9766 17490 9818
rect 17490 9766 17536 9818
rect 17240 9764 17296 9766
rect 17320 9764 17376 9766
rect 17400 9764 17456 9766
rect 17480 9764 17536 9766
rect 14526 7098 14582 7100
rect 14606 7098 14662 7100
rect 14686 7098 14742 7100
rect 14766 7098 14822 7100
rect 14526 7046 14572 7098
rect 14572 7046 14582 7098
rect 14606 7046 14636 7098
rect 14636 7046 14648 7098
rect 14648 7046 14662 7098
rect 14686 7046 14700 7098
rect 14700 7046 14712 7098
rect 14712 7046 14742 7098
rect 14766 7046 14776 7098
rect 14776 7046 14822 7098
rect 14526 7044 14582 7046
rect 14606 7044 14662 7046
rect 14686 7044 14742 7046
rect 14766 7044 14822 7046
rect 17240 8730 17296 8732
rect 17320 8730 17376 8732
rect 17400 8730 17456 8732
rect 17480 8730 17536 8732
rect 17240 8678 17286 8730
rect 17286 8678 17296 8730
rect 17320 8678 17350 8730
rect 17350 8678 17362 8730
rect 17362 8678 17376 8730
rect 17400 8678 17414 8730
rect 17414 8678 17426 8730
rect 17426 8678 17456 8730
rect 17480 8678 17490 8730
rect 17490 8678 17536 8730
rect 17240 8676 17296 8678
rect 17320 8676 17376 8678
rect 17400 8676 17456 8678
rect 17480 8676 17536 8678
rect 16946 7928 17002 7984
rect 18234 10668 18290 10704
rect 18234 10648 18236 10668
rect 18236 10648 18288 10668
rect 18288 10648 18290 10668
rect 18418 9968 18474 10024
rect 17240 7642 17296 7644
rect 17320 7642 17376 7644
rect 17400 7642 17456 7644
rect 17480 7642 17536 7644
rect 17240 7590 17286 7642
rect 17286 7590 17296 7642
rect 17320 7590 17350 7642
rect 17350 7590 17362 7642
rect 17362 7590 17376 7642
rect 17400 7590 17414 7642
rect 17414 7590 17426 7642
rect 17426 7590 17456 7642
rect 17480 7590 17490 7642
rect 17490 7590 17536 7642
rect 17240 7588 17296 7590
rect 17320 7588 17376 7590
rect 17400 7588 17456 7590
rect 17480 7588 17536 7590
rect 19954 17978 20010 17980
rect 20034 17978 20090 17980
rect 20114 17978 20170 17980
rect 20194 17978 20250 17980
rect 19954 17926 20000 17978
rect 20000 17926 20010 17978
rect 20034 17926 20064 17978
rect 20064 17926 20076 17978
rect 20076 17926 20090 17978
rect 20114 17926 20128 17978
rect 20128 17926 20140 17978
rect 20140 17926 20170 17978
rect 20194 17926 20204 17978
rect 20204 17926 20250 17978
rect 19954 17924 20010 17926
rect 20034 17924 20090 17926
rect 20114 17924 20170 17926
rect 20194 17924 20250 17926
rect 19954 16890 20010 16892
rect 20034 16890 20090 16892
rect 20114 16890 20170 16892
rect 20194 16890 20250 16892
rect 19954 16838 20000 16890
rect 20000 16838 20010 16890
rect 20034 16838 20064 16890
rect 20064 16838 20076 16890
rect 20076 16838 20090 16890
rect 20114 16838 20128 16890
rect 20128 16838 20140 16890
rect 20140 16838 20170 16890
rect 20194 16838 20204 16890
rect 20204 16838 20250 16890
rect 19954 16836 20010 16838
rect 20034 16836 20090 16838
rect 20114 16836 20170 16838
rect 20194 16836 20250 16838
rect 19954 15802 20010 15804
rect 20034 15802 20090 15804
rect 20114 15802 20170 15804
rect 20194 15802 20250 15804
rect 19954 15750 20000 15802
rect 20000 15750 20010 15802
rect 20034 15750 20064 15802
rect 20064 15750 20076 15802
rect 20076 15750 20090 15802
rect 20114 15750 20128 15802
rect 20128 15750 20140 15802
rect 20140 15750 20170 15802
rect 20194 15750 20204 15802
rect 20204 15750 20250 15802
rect 19954 15748 20010 15750
rect 20034 15748 20090 15750
rect 20114 15748 20170 15750
rect 20194 15748 20250 15750
rect 19954 14714 20010 14716
rect 20034 14714 20090 14716
rect 20114 14714 20170 14716
rect 20194 14714 20250 14716
rect 19954 14662 20000 14714
rect 20000 14662 20010 14714
rect 20034 14662 20064 14714
rect 20064 14662 20076 14714
rect 20076 14662 20090 14714
rect 20114 14662 20128 14714
rect 20128 14662 20140 14714
rect 20140 14662 20170 14714
rect 20194 14662 20204 14714
rect 20204 14662 20250 14714
rect 19954 14660 20010 14662
rect 20034 14660 20090 14662
rect 20114 14660 20170 14662
rect 20194 14660 20250 14662
rect 22668 20698 22724 20700
rect 22748 20698 22804 20700
rect 22828 20698 22884 20700
rect 22908 20698 22964 20700
rect 22668 20646 22714 20698
rect 22714 20646 22724 20698
rect 22748 20646 22778 20698
rect 22778 20646 22790 20698
rect 22790 20646 22804 20698
rect 22828 20646 22842 20698
rect 22842 20646 22854 20698
rect 22854 20646 22884 20698
rect 22908 20646 22918 20698
rect 22918 20646 22964 20698
rect 22668 20644 22724 20646
rect 22748 20644 22804 20646
rect 22828 20644 22884 20646
rect 22908 20644 22964 20646
rect 22668 19610 22724 19612
rect 22748 19610 22804 19612
rect 22828 19610 22884 19612
rect 22908 19610 22964 19612
rect 22668 19558 22714 19610
rect 22714 19558 22724 19610
rect 22748 19558 22778 19610
rect 22778 19558 22790 19610
rect 22790 19558 22804 19610
rect 22828 19558 22842 19610
rect 22842 19558 22854 19610
rect 22854 19558 22884 19610
rect 22908 19558 22918 19610
rect 22918 19558 22964 19610
rect 22668 19556 22724 19558
rect 22748 19556 22804 19558
rect 22828 19556 22884 19558
rect 22908 19556 22964 19558
rect 22668 18522 22724 18524
rect 22748 18522 22804 18524
rect 22828 18522 22884 18524
rect 22908 18522 22964 18524
rect 22668 18470 22714 18522
rect 22714 18470 22724 18522
rect 22748 18470 22778 18522
rect 22778 18470 22790 18522
rect 22790 18470 22804 18522
rect 22828 18470 22842 18522
rect 22842 18470 22854 18522
rect 22854 18470 22884 18522
rect 22908 18470 22918 18522
rect 22918 18470 22964 18522
rect 22668 18468 22724 18470
rect 22748 18468 22804 18470
rect 22828 18468 22884 18470
rect 22908 18468 22964 18470
rect 22668 17434 22724 17436
rect 22748 17434 22804 17436
rect 22828 17434 22884 17436
rect 22908 17434 22964 17436
rect 22668 17382 22714 17434
rect 22714 17382 22724 17434
rect 22748 17382 22778 17434
rect 22778 17382 22790 17434
rect 22790 17382 22804 17434
rect 22828 17382 22842 17434
rect 22842 17382 22854 17434
rect 22854 17382 22884 17434
rect 22908 17382 22918 17434
rect 22918 17382 22964 17434
rect 22668 17380 22724 17382
rect 22748 17380 22804 17382
rect 22828 17380 22884 17382
rect 22908 17380 22964 17382
rect 22668 16346 22724 16348
rect 22748 16346 22804 16348
rect 22828 16346 22884 16348
rect 22908 16346 22964 16348
rect 22668 16294 22714 16346
rect 22714 16294 22724 16346
rect 22748 16294 22778 16346
rect 22778 16294 22790 16346
rect 22790 16294 22804 16346
rect 22828 16294 22842 16346
rect 22842 16294 22854 16346
rect 22854 16294 22884 16346
rect 22908 16294 22918 16346
rect 22918 16294 22964 16346
rect 22668 16292 22724 16294
rect 22748 16292 22804 16294
rect 22828 16292 22884 16294
rect 22908 16292 22964 16294
rect 22668 15258 22724 15260
rect 22748 15258 22804 15260
rect 22828 15258 22884 15260
rect 22908 15258 22964 15260
rect 22668 15206 22714 15258
rect 22714 15206 22724 15258
rect 22748 15206 22778 15258
rect 22778 15206 22790 15258
rect 22790 15206 22804 15258
rect 22828 15206 22842 15258
rect 22842 15206 22854 15258
rect 22854 15206 22884 15258
rect 22908 15206 22918 15258
rect 22918 15206 22964 15258
rect 22668 15204 22724 15206
rect 22748 15204 22804 15206
rect 22828 15204 22884 15206
rect 22908 15204 22964 15206
rect 19954 13626 20010 13628
rect 20034 13626 20090 13628
rect 20114 13626 20170 13628
rect 20194 13626 20250 13628
rect 19954 13574 20000 13626
rect 20000 13574 20010 13626
rect 20034 13574 20064 13626
rect 20064 13574 20076 13626
rect 20076 13574 20090 13626
rect 20114 13574 20128 13626
rect 20128 13574 20140 13626
rect 20140 13574 20170 13626
rect 20194 13574 20204 13626
rect 20204 13574 20250 13626
rect 19954 13572 20010 13574
rect 20034 13572 20090 13574
rect 20114 13572 20170 13574
rect 20194 13572 20250 13574
rect 19954 12538 20010 12540
rect 20034 12538 20090 12540
rect 20114 12538 20170 12540
rect 20194 12538 20250 12540
rect 19954 12486 20000 12538
rect 20000 12486 20010 12538
rect 20034 12486 20064 12538
rect 20064 12486 20076 12538
rect 20076 12486 20090 12538
rect 20114 12486 20128 12538
rect 20128 12486 20140 12538
rect 20140 12486 20170 12538
rect 20194 12486 20204 12538
rect 20204 12486 20250 12538
rect 19954 12484 20010 12486
rect 20034 12484 20090 12486
rect 20114 12484 20170 12486
rect 20194 12484 20250 12486
rect 19954 11450 20010 11452
rect 20034 11450 20090 11452
rect 20114 11450 20170 11452
rect 20194 11450 20250 11452
rect 19954 11398 20000 11450
rect 20000 11398 20010 11450
rect 20034 11398 20064 11450
rect 20064 11398 20076 11450
rect 20076 11398 20090 11450
rect 20114 11398 20128 11450
rect 20128 11398 20140 11450
rect 20140 11398 20170 11450
rect 20194 11398 20204 11450
rect 20204 11398 20250 11450
rect 19954 11396 20010 11398
rect 20034 11396 20090 11398
rect 20114 11396 20170 11398
rect 20194 11396 20250 11398
rect 19954 10362 20010 10364
rect 20034 10362 20090 10364
rect 20114 10362 20170 10364
rect 20194 10362 20250 10364
rect 19954 10310 20000 10362
rect 20000 10310 20010 10362
rect 20034 10310 20064 10362
rect 20064 10310 20076 10362
rect 20076 10310 20090 10362
rect 20114 10310 20128 10362
rect 20128 10310 20140 10362
rect 20140 10310 20170 10362
rect 20194 10310 20204 10362
rect 20204 10310 20250 10362
rect 19954 10308 20010 10310
rect 20034 10308 20090 10310
rect 20114 10308 20170 10310
rect 20194 10308 20250 10310
rect 22668 14170 22724 14172
rect 22748 14170 22804 14172
rect 22828 14170 22884 14172
rect 22908 14170 22964 14172
rect 22668 14118 22714 14170
rect 22714 14118 22724 14170
rect 22748 14118 22778 14170
rect 22778 14118 22790 14170
rect 22790 14118 22804 14170
rect 22828 14118 22842 14170
rect 22842 14118 22854 14170
rect 22854 14118 22884 14170
rect 22908 14118 22918 14170
rect 22918 14118 22964 14170
rect 22668 14116 22724 14118
rect 22748 14116 22804 14118
rect 22828 14116 22884 14118
rect 22908 14116 22964 14118
rect 19954 9274 20010 9276
rect 20034 9274 20090 9276
rect 20114 9274 20170 9276
rect 20194 9274 20250 9276
rect 19954 9222 20000 9274
rect 20000 9222 20010 9274
rect 20034 9222 20064 9274
rect 20064 9222 20076 9274
rect 20076 9222 20090 9274
rect 20114 9222 20128 9274
rect 20128 9222 20140 9274
rect 20140 9222 20170 9274
rect 20194 9222 20204 9274
rect 20204 9222 20250 9274
rect 19954 9220 20010 9222
rect 20034 9220 20090 9222
rect 20114 9220 20170 9222
rect 20194 9220 20250 9222
rect 19954 8186 20010 8188
rect 20034 8186 20090 8188
rect 20114 8186 20170 8188
rect 20194 8186 20250 8188
rect 19954 8134 20000 8186
rect 20000 8134 20010 8186
rect 20034 8134 20064 8186
rect 20064 8134 20076 8186
rect 20076 8134 20090 8186
rect 20114 8134 20128 8186
rect 20128 8134 20140 8186
rect 20140 8134 20170 8186
rect 20194 8134 20204 8186
rect 20204 8134 20250 8186
rect 19954 8132 20010 8134
rect 20034 8132 20090 8134
rect 20114 8132 20170 8134
rect 20194 8132 20250 8134
rect 19954 7098 20010 7100
rect 20034 7098 20090 7100
rect 20114 7098 20170 7100
rect 20194 7098 20250 7100
rect 19954 7046 20000 7098
rect 20000 7046 20010 7098
rect 20034 7046 20064 7098
rect 20064 7046 20076 7098
rect 20076 7046 20090 7098
rect 20114 7046 20128 7098
rect 20128 7046 20140 7098
rect 20140 7046 20170 7098
rect 20194 7046 20204 7098
rect 20204 7046 20250 7098
rect 19954 7044 20010 7046
rect 20034 7044 20090 7046
rect 20114 7044 20170 7046
rect 20194 7044 20250 7046
rect 11812 6554 11868 6556
rect 11892 6554 11948 6556
rect 11972 6554 12028 6556
rect 12052 6554 12108 6556
rect 11812 6502 11858 6554
rect 11858 6502 11868 6554
rect 11892 6502 11922 6554
rect 11922 6502 11934 6554
rect 11934 6502 11948 6554
rect 11972 6502 11986 6554
rect 11986 6502 11998 6554
rect 11998 6502 12028 6554
rect 12052 6502 12062 6554
rect 12062 6502 12108 6554
rect 11812 6500 11868 6502
rect 11892 6500 11948 6502
rect 11972 6500 12028 6502
rect 12052 6500 12108 6502
rect 17240 6554 17296 6556
rect 17320 6554 17376 6556
rect 17400 6554 17456 6556
rect 17480 6554 17536 6556
rect 17240 6502 17286 6554
rect 17286 6502 17296 6554
rect 17320 6502 17350 6554
rect 17350 6502 17362 6554
rect 17362 6502 17376 6554
rect 17400 6502 17414 6554
rect 17414 6502 17426 6554
rect 17426 6502 17456 6554
rect 17480 6502 17490 6554
rect 17490 6502 17536 6554
rect 17240 6500 17296 6502
rect 17320 6500 17376 6502
rect 17400 6500 17456 6502
rect 17480 6500 17536 6502
rect 14526 6010 14582 6012
rect 14606 6010 14662 6012
rect 14686 6010 14742 6012
rect 14766 6010 14822 6012
rect 14526 5958 14572 6010
rect 14572 5958 14582 6010
rect 14606 5958 14636 6010
rect 14636 5958 14648 6010
rect 14648 5958 14662 6010
rect 14686 5958 14700 6010
rect 14700 5958 14712 6010
rect 14712 5958 14742 6010
rect 14766 5958 14776 6010
rect 14776 5958 14822 6010
rect 14526 5956 14582 5958
rect 14606 5956 14662 5958
rect 14686 5956 14742 5958
rect 14766 5956 14822 5958
rect 19954 6010 20010 6012
rect 20034 6010 20090 6012
rect 20114 6010 20170 6012
rect 20194 6010 20250 6012
rect 19954 5958 20000 6010
rect 20000 5958 20010 6010
rect 20034 5958 20064 6010
rect 20064 5958 20076 6010
rect 20076 5958 20090 6010
rect 20114 5958 20128 6010
rect 20128 5958 20140 6010
rect 20140 5958 20170 6010
rect 20194 5958 20204 6010
rect 20204 5958 20250 6010
rect 19954 5956 20010 5958
rect 20034 5956 20090 5958
rect 20114 5956 20170 5958
rect 20194 5956 20250 5958
rect 11812 5466 11868 5468
rect 11892 5466 11948 5468
rect 11972 5466 12028 5468
rect 12052 5466 12108 5468
rect 11812 5414 11858 5466
rect 11858 5414 11868 5466
rect 11892 5414 11922 5466
rect 11922 5414 11934 5466
rect 11934 5414 11948 5466
rect 11972 5414 11986 5466
rect 11986 5414 11998 5466
rect 11998 5414 12028 5466
rect 12052 5414 12062 5466
rect 12062 5414 12108 5466
rect 11812 5412 11868 5414
rect 11892 5412 11948 5414
rect 11972 5412 12028 5414
rect 12052 5412 12108 5414
rect 17240 5466 17296 5468
rect 17320 5466 17376 5468
rect 17400 5466 17456 5468
rect 17480 5466 17536 5468
rect 17240 5414 17286 5466
rect 17286 5414 17296 5466
rect 17320 5414 17350 5466
rect 17350 5414 17362 5466
rect 17362 5414 17376 5466
rect 17400 5414 17414 5466
rect 17414 5414 17426 5466
rect 17426 5414 17456 5466
rect 17480 5414 17490 5466
rect 17490 5414 17536 5466
rect 17240 5412 17296 5414
rect 17320 5412 17376 5414
rect 17400 5412 17456 5414
rect 17480 5412 17536 5414
rect 14526 4922 14582 4924
rect 14606 4922 14662 4924
rect 14686 4922 14742 4924
rect 14766 4922 14822 4924
rect 14526 4870 14572 4922
rect 14572 4870 14582 4922
rect 14606 4870 14636 4922
rect 14636 4870 14648 4922
rect 14648 4870 14662 4922
rect 14686 4870 14700 4922
rect 14700 4870 14712 4922
rect 14712 4870 14742 4922
rect 14766 4870 14776 4922
rect 14776 4870 14822 4922
rect 14526 4868 14582 4870
rect 14606 4868 14662 4870
rect 14686 4868 14742 4870
rect 14766 4868 14822 4870
rect 19954 4922 20010 4924
rect 20034 4922 20090 4924
rect 20114 4922 20170 4924
rect 20194 4922 20250 4924
rect 19954 4870 20000 4922
rect 20000 4870 20010 4922
rect 20034 4870 20064 4922
rect 20064 4870 20076 4922
rect 20076 4870 20090 4922
rect 20114 4870 20128 4922
rect 20128 4870 20140 4922
rect 20140 4870 20170 4922
rect 20194 4870 20204 4922
rect 20204 4870 20250 4922
rect 19954 4868 20010 4870
rect 20034 4868 20090 4870
rect 20114 4868 20170 4870
rect 20194 4868 20250 4870
rect 11812 4378 11868 4380
rect 11892 4378 11948 4380
rect 11972 4378 12028 4380
rect 12052 4378 12108 4380
rect 11812 4326 11858 4378
rect 11858 4326 11868 4378
rect 11892 4326 11922 4378
rect 11922 4326 11934 4378
rect 11934 4326 11948 4378
rect 11972 4326 11986 4378
rect 11986 4326 11998 4378
rect 11998 4326 12028 4378
rect 12052 4326 12062 4378
rect 12062 4326 12108 4378
rect 11812 4324 11868 4326
rect 11892 4324 11948 4326
rect 11972 4324 12028 4326
rect 12052 4324 12108 4326
rect 17240 4378 17296 4380
rect 17320 4378 17376 4380
rect 17400 4378 17456 4380
rect 17480 4378 17536 4380
rect 17240 4326 17286 4378
rect 17286 4326 17296 4378
rect 17320 4326 17350 4378
rect 17350 4326 17362 4378
rect 17362 4326 17376 4378
rect 17400 4326 17414 4378
rect 17414 4326 17426 4378
rect 17426 4326 17456 4378
rect 17480 4326 17490 4378
rect 17490 4326 17536 4378
rect 17240 4324 17296 4326
rect 17320 4324 17376 4326
rect 17400 4324 17456 4326
rect 17480 4324 17536 4326
rect 14526 3834 14582 3836
rect 14606 3834 14662 3836
rect 14686 3834 14742 3836
rect 14766 3834 14822 3836
rect 14526 3782 14572 3834
rect 14572 3782 14582 3834
rect 14606 3782 14636 3834
rect 14636 3782 14648 3834
rect 14648 3782 14662 3834
rect 14686 3782 14700 3834
rect 14700 3782 14712 3834
rect 14712 3782 14742 3834
rect 14766 3782 14776 3834
rect 14776 3782 14822 3834
rect 14526 3780 14582 3782
rect 14606 3780 14662 3782
rect 14686 3780 14742 3782
rect 14766 3780 14822 3782
rect 19954 3834 20010 3836
rect 20034 3834 20090 3836
rect 20114 3834 20170 3836
rect 20194 3834 20250 3836
rect 19954 3782 20000 3834
rect 20000 3782 20010 3834
rect 20034 3782 20064 3834
rect 20064 3782 20076 3834
rect 20076 3782 20090 3834
rect 20114 3782 20128 3834
rect 20128 3782 20140 3834
rect 20140 3782 20170 3834
rect 20194 3782 20204 3834
rect 20204 3782 20250 3834
rect 19954 3780 20010 3782
rect 20034 3780 20090 3782
rect 20114 3780 20170 3782
rect 20194 3780 20250 3782
rect 11812 3290 11868 3292
rect 11892 3290 11948 3292
rect 11972 3290 12028 3292
rect 12052 3290 12108 3292
rect 11812 3238 11858 3290
rect 11858 3238 11868 3290
rect 11892 3238 11922 3290
rect 11922 3238 11934 3290
rect 11934 3238 11948 3290
rect 11972 3238 11986 3290
rect 11986 3238 11998 3290
rect 11998 3238 12028 3290
rect 12052 3238 12062 3290
rect 12062 3238 12108 3290
rect 11812 3236 11868 3238
rect 11892 3236 11948 3238
rect 11972 3236 12028 3238
rect 12052 3236 12108 3238
rect 17240 3290 17296 3292
rect 17320 3290 17376 3292
rect 17400 3290 17456 3292
rect 17480 3290 17536 3292
rect 17240 3238 17286 3290
rect 17286 3238 17296 3290
rect 17320 3238 17350 3290
rect 17350 3238 17362 3290
rect 17362 3238 17376 3290
rect 17400 3238 17414 3290
rect 17414 3238 17426 3290
rect 17426 3238 17456 3290
rect 17480 3238 17490 3290
rect 17490 3238 17536 3290
rect 17240 3236 17296 3238
rect 17320 3236 17376 3238
rect 17400 3236 17456 3238
rect 17480 3236 17536 3238
rect 14526 2746 14582 2748
rect 14606 2746 14662 2748
rect 14686 2746 14742 2748
rect 14766 2746 14822 2748
rect 14526 2694 14572 2746
rect 14572 2694 14582 2746
rect 14606 2694 14636 2746
rect 14636 2694 14648 2746
rect 14648 2694 14662 2746
rect 14686 2694 14700 2746
rect 14700 2694 14712 2746
rect 14712 2694 14742 2746
rect 14766 2694 14776 2746
rect 14776 2694 14822 2746
rect 14526 2692 14582 2694
rect 14606 2692 14662 2694
rect 14686 2692 14742 2694
rect 14766 2692 14822 2694
rect 19954 2746 20010 2748
rect 20034 2746 20090 2748
rect 20114 2746 20170 2748
rect 20194 2746 20250 2748
rect 19954 2694 20000 2746
rect 20000 2694 20010 2746
rect 20034 2694 20064 2746
rect 20064 2694 20076 2746
rect 20076 2694 20090 2746
rect 20114 2694 20128 2746
rect 20128 2694 20140 2746
rect 20140 2694 20170 2746
rect 20194 2694 20204 2746
rect 20204 2694 20250 2746
rect 19954 2692 20010 2694
rect 20034 2692 20090 2694
rect 20114 2692 20170 2694
rect 20194 2692 20250 2694
rect 22668 13082 22724 13084
rect 22748 13082 22804 13084
rect 22828 13082 22884 13084
rect 22908 13082 22964 13084
rect 22668 13030 22714 13082
rect 22714 13030 22724 13082
rect 22748 13030 22778 13082
rect 22778 13030 22790 13082
rect 22790 13030 22804 13082
rect 22828 13030 22842 13082
rect 22842 13030 22854 13082
rect 22854 13030 22884 13082
rect 22908 13030 22918 13082
rect 22918 13030 22964 13082
rect 22668 13028 22724 13030
rect 22748 13028 22804 13030
rect 22828 13028 22884 13030
rect 22908 13028 22964 13030
rect 22668 11994 22724 11996
rect 22748 11994 22804 11996
rect 22828 11994 22884 11996
rect 22908 11994 22964 11996
rect 22668 11942 22714 11994
rect 22714 11942 22724 11994
rect 22748 11942 22778 11994
rect 22778 11942 22790 11994
rect 22790 11942 22804 11994
rect 22828 11942 22842 11994
rect 22842 11942 22854 11994
rect 22854 11942 22884 11994
rect 22908 11942 22918 11994
rect 22918 11942 22964 11994
rect 22668 11940 22724 11942
rect 22748 11940 22804 11942
rect 22828 11940 22884 11942
rect 22908 11940 22964 11942
rect 22668 10906 22724 10908
rect 22748 10906 22804 10908
rect 22828 10906 22884 10908
rect 22908 10906 22964 10908
rect 22668 10854 22714 10906
rect 22714 10854 22724 10906
rect 22748 10854 22778 10906
rect 22778 10854 22790 10906
rect 22790 10854 22804 10906
rect 22828 10854 22842 10906
rect 22842 10854 22854 10906
rect 22854 10854 22884 10906
rect 22908 10854 22918 10906
rect 22918 10854 22964 10906
rect 22668 10852 22724 10854
rect 22748 10852 22804 10854
rect 22828 10852 22884 10854
rect 22908 10852 22964 10854
rect 22668 9818 22724 9820
rect 22748 9818 22804 9820
rect 22828 9818 22884 9820
rect 22908 9818 22964 9820
rect 22668 9766 22714 9818
rect 22714 9766 22724 9818
rect 22748 9766 22778 9818
rect 22778 9766 22790 9818
rect 22790 9766 22804 9818
rect 22828 9766 22842 9818
rect 22842 9766 22854 9818
rect 22854 9766 22884 9818
rect 22908 9766 22918 9818
rect 22918 9766 22964 9818
rect 22668 9764 22724 9766
rect 22748 9764 22804 9766
rect 22828 9764 22884 9766
rect 22908 9764 22964 9766
rect 22668 8730 22724 8732
rect 22748 8730 22804 8732
rect 22828 8730 22884 8732
rect 22908 8730 22964 8732
rect 22668 8678 22714 8730
rect 22714 8678 22724 8730
rect 22748 8678 22778 8730
rect 22778 8678 22790 8730
rect 22790 8678 22804 8730
rect 22828 8678 22842 8730
rect 22842 8678 22854 8730
rect 22854 8678 22884 8730
rect 22908 8678 22918 8730
rect 22918 8678 22964 8730
rect 22668 8676 22724 8678
rect 22748 8676 22804 8678
rect 22828 8676 22884 8678
rect 22908 8676 22964 8678
rect 22668 7642 22724 7644
rect 22748 7642 22804 7644
rect 22828 7642 22884 7644
rect 22908 7642 22964 7644
rect 22668 7590 22714 7642
rect 22714 7590 22724 7642
rect 22748 7590 22778 7642
rect 22778 7590 22790 7642
rect 22790 7590 22804 7642
rect 22828 7590 22842 7642
rect 22842 7590 22854 7642
rect 22854 7590 22884 7642
rect 22908 7590 22918 7642
rect 22918 7590 22964 7642
rect 22668 7588 22724 7590
rect 22748 7588 22804 7590
rect 22828 7588 22884 7590
rect 22908 7588 22964 7590
rect 22668 6554 22724 6556
rect 22748 6554 22804 6556
rect 22828 6554 22884 6556
rect 22908 6554 22964 6556
rect 22668 6502 22714 6554
rect 22714 6502 22724 6554
rect 22748 6502 22778 6554
rect 22778 6502 22790 6554
rect 22790 6502 22804 6554
rect 22828 6502 22842 6554
rect 22842 6502 22854 6554
rect 22854 6502 22884 6554
rect 22908 6502 22918 6554
rect 22918 6502 22964 6554
rect 22668 6500 22724 6502
rect 22748 6500 22804 6502
rect 22828 6500 22884 6502
rect 22908 6500 22964 6502
rect 22668 5466 22724 5468
rect 22748 5466 22804 5468
rect 22828 5466 22884 5468
rect 22908 5466 22964 5468
rect 22668 5414 22714 5466
rect 22714 5414 22724 5466
rect 22748 5414 22778 5466
rect 22778 5414 22790 5466
rect 22790 5414 22804 5466
rect 22828 5414 22842 5466
rect 22842 5414 22854 5466
rect 22854 5414 22884 5466
rect 22908 5414 22918 5466
rect 22918 5414 22964 5466
rect 22668 5412 22724 5414
rect 22748 5412 22804 5414
rect 22828 5412 22884 5414
rect 22908 5412 22964 5414
rect 22668 4378 22724 4380
rect 22748 4378 22804 4380
rect 22828 4378 22884 4380
rect 22908 4378 22964 4380
rect 22668 4326 22714 4378
rect 22714 4326 22724 4378
rect 22748 4326 22778 4378
rect 22778 4326 22790 4378
rect 22790 4326 22804 4378
rect 22828 4326 22842 4378
rect 22842 4326 22854 4378
rect 22854 4326 22884 4378
rect 22908 4326 22918 4378
rect 22918 4326 22964 4378
rect 22668 4324 22724 4326
rect 22748 4324 22804 4326
rect 22828 4324 22884 4326
rect 22908 4324 22964 4326
rect 22668 3290 22724 3292
rect 22748 3290 22804 3292
rect 22828 3290 22884 3292
rect 22908 3290 22964 3292
rect 22668 3238 22714 3290
rect 22714 3238 22724 3290
rect 22748 3238 22778 3290
rect 22778 3238 22790 3290
rect 22790 3238 22804 3290
rect 22828 3238 22842 3290
rect 22842 3238 22854 3290
rect 22854 3238 22884 3290
rect 22908 3238 22918 3290
rect 22918 3238 22964 3290
rect 22668 3236 22724 3238
rect 22748 3236 22804 3238
rect 22828 3236 22884 3238
rect 22908 3236 22964 3238
rect 6384 2202 6440 2204
rect 6464 2202 6520 2204
rect 6544 2202 6600 2204
rect 6624 2202 6680 2204
rect 6384 2150 6430 2202
rect 6430 2150 6440 2202
rect 6464 2150 6494 2202
rect 6494 2150 6506 2202
rect 6506 2150 6520 2202
rect 6544 2150 6558 2202
rect 6558 2150 6570 2202
rect 6570 2150 6600 2202
rect 6624 2150 6634 2202
rect 6634 2150 6680 2202
rect 6384 2148 6440 2150
rect 6464 2148 6520 2150
rect 6544 2148 6600 2150
rect 6624 2148 6680 2150
rect 11812 2202 11868 2204
rect 11892 2202 11948 2204
rect 11972 2202 12028 2204
rect 12052 2202 12108 2204
rect 11812 2150 11858 2202
rect 11858 2150 11868 2202
rect 11892 2150 11922 2202
rect 11922 2150 11934 2202
rect 11934 2150 11948 2202
rect 11972 2150 11986 2202
rect 11986 2150 11998 2202
rect 11998 2150 12028 2202
rect 12052 2150 12062 2202
rect 12062 2150 12108 2202
rect 11812 2148 11868 2150
rect 11892 2148 11948 2150
rect 11972 2148 12028 2150
rect 12052 2148 12108 2150
rect 17240 2202 17296 2204
rect 17320 2202 17376 2204
rect 17400 2202 17456 2204
rect 17480 2202 17536 2204
rect 17240 2150 17286 2202
rect 17286 2150 17296 2202
rect 17320 2150 17350 2202
rect 17350 2150 17362 2202
rect 17362 2150 17376 2202
rect 17400 2150 17414 2202
rect 17414 2150 17426 2202
rect 17426 2150 17456 2202
rect 17480 2150 17490 2202
rect 17490 2150 17536 2202
rect 17240 2148 17296 2150
rect 17320 2148 17376 2150
rect 17400 2148 17456 2150
rect 17480 2148 17536 2150
rect 22668 2202 22724 2204
rect 22748 2202 22804 2204
rect 22828 2202 22884 2204
rect 22908 2202 22964 2204
rect 22668 2150 22714 2202
rect 22714 2150 22724 2202
rect 22748 2150 22778 2202
rect 22778 2150 22790 2202
rect 22790 2150 22804 2202
rect 22828 2150 22842 2202
rect 22842 2150 22854 2202
rect 22854 2150 22884 2202
rect 22908 2150 22918 2202
rect 22918 2150 22964 2202
rect 22668 2148 22724 2150
rect 22748 2148 22804 2150
rect 22828 2148 22884 2150
rect 22908 2148 22964 2150
<< metal3 >>
rect 6374 21792 6690 21793
rect 6374 21728 6380 21792
rect 6444 21728 6460 21792
rect 6524 21728 6540 21792
rect 6604 21728 6620 21792
rect 6684 21728 6690 21792
rect 6374 21727 6690 21728
rect 11802 21792 12118 21793
rect 11802 21728 11808 21792
rect 11872 21728 11888 21792
rect 11952 21728 11968 21792
rect 12032 21728 12048 21792
rect 12112 21728 12118 21792
rect 11802 21727 12118 21728
rect 17230 21792 17546 21793
rect 17230 21728 17236 21792
rect 17300 21728 17316 21792
rect 17380 21728 17396 21792
rect 17460 21728 17476 21792
rect 17540 21728 17546 21792
rect 17230 21727 17546 21728
rect 22658 21792 22974 21793
rect 22658 21728 22664 21792
rect 22728 21728 22744 21792
rect 22808 21728 22824 21792
rect 22888 21728 22904 21792
rect 22968 21728 22974 21792
rect 22658 21727 22974 21728
rect 3660 21248 3976 21249
rect 3660 21184 3666 21248
rect 3730 21184 3746 21248
rect 3810 21184 3826 21248
rect 3890 21184 3906 21248
rect 3970 21184 3976 21248
rect 3660 21183 3976 21184
rect 9088 21248 9404 21249
rect 9088 21184 9094 21248
rect 9158 21184 9174 21248
rect 9238 21184 9254 21248
rect 9318 21184 9334 21248
rect 9398 21184 9404 21248
rect 9088 21183 9404 21184
rect 14516 21248 14832 21249
rect 14516 21184 14522 21248
rect 14586 21184 14602 21248
rect 14666 21184 14682 21248
rect 14746 21184 14762 21248
rect 14826 21184 14832 21248
rect 14516 21183 14832 21184
rect 19944 21248 20260 21249
rect 19944 21184 19950 21248
rect 20014 21184 20030 21248
rect 20094 21184 20110 21248
rect 20174 21184 20190 21248
rect 20254 21184 20260 21248
rect 19944 21183 20260 21184
rect 16297 21042 16363 21045
rect 17309 21042 17375 21045
rect 16297 21040 17375 21042
rect 16297 20984 16302 21040
rect 16358 20984 17314 21040
rect 17370 20984 17375 21040
rect 16297 20982 17375 20984
rect 16297 20979 16363 20982
rect 17309 20979 17375 20982
rect 6374 20704 6690 20705
rect 6374 20640 6380 20704
rect 6444 20640 6460 20704
rect 6524 20640 6540 20704
rect 6604 20640 6620 20704
rect 6684 20640 6690 20704
rect 6374 20639 6690 20640
rect 11802 20704 12118 20705
rect 11802 20640 11808 20704
rect 11872 20640 11888 20704
rect 11952 20640 11968 20704
rect 12032 20640 12048 20704
rect 12112 20640 12118 20704
rect 11802 20639 12118 20640
rect 17230 20704 17546 20705
rect 17230 20640 17236 20704
rect 17300 20640 17316 20704
rect 17380 20640 17396 20704
rect 17460 20640 17476 20704
rect 17540 20640 17546 20704
rect 17230 20639 17546 20640
rect 22658 20704 22974 20705
rect 22658 20640 22664 20704
rect 22728 20640 22744 20704
rect 22808 20640 22824 20704
rect 22888 20640 22904 20704
rect 22968 20640 22974 20704
rect 22658 20639 22974 20640
rect 3660 20160 3976 20161
rect 3660 20096 3666 20160
rect 3730 20096 3746 20160
rect 3810 20096 3826 20160
rect 3890 20096 3906 20160
rect 3970 20096 3976 20160
rect 3660 20095 3976 20096
rect 9088 20160 9404 20161
rect 9088 20096 9094 20160
rect 9158 20096 9174 20160
rect 9238 20096 9254 20160
rect 9318 20096 9334 20160
rect 9398 20096 9404 20160
rect 9088 20095 9404 20096
rect 14516 20160 14832 20161
rect 14516 20096 14522 20160
rect 14586 20096 14602 20160
rect 14666 20096 14682 20160
rect 14746 20096 14762 20160
rect 14826 20096 14832 20160
rect 14516 20095 14832 20096
rect 19944 20160 20260 20161
rect 19944 20096 19950 20160
rect 20014 20096 20030 20160
rect 20094 20096 20110 20160
rect 20174 20096 20190 20160
rect 20254 20096 20260 20160
rect 19944 20095 20260 20096
rect 6374 19616 6690 19617
rect 6374 19552 6380 19616
rect 6444 19552 6460 19616
rect 6524 19552 6540 19616
rect 6604 19552 6620 19616
rect 6684 19552 6690 19616
rect 6374 19551 6690 19552
rect 11802 19616 12118 19617
rect 11802 19552 11808 19616
rect 11872 19552 11888 19616
rect 11952 19552 11968 19616
rect 12032 19552 12048 19616
rect 12112 19552 12118 19616
rect 11802 19551 12118 19552
rect 17230 19616 17546 19617
rect 17230 19552 17236 19616
rect 17300 19552 17316 19616
rect 17380 19552 17396 19616
rect 17460 19552 17476 19616
rect 17540 19552 17546 19616
rect 17230 19551 17546 19552
rect 22658 19616 22974 19617
rect 22658 19552 22664 19616
rect 22728 19552 22744 19616
rect 22808 19552 22824 19616
rect 22888 19552 22904 19616
rect 22968 19552 22974 19616
rect 22658 19551 22974 19552
rect 3660 19072 3976 19073
rect 3660 19008 3666 19072
rect 3730 19008 3746 19072
rect 3810 19008 3826 19072
rect 3890 19008 3906 19072
rect 3970 19008 3976 19072
rect 3660 19007 3976 19008
rect 9088 19072 9404 19073
rect 9088 19008 9094 19072
rect 9158 19008 9174 19072
rect 9238 19008 9254 19072
rect 9318 19008 9334 19072
rect 9398 19008 9404 19072
rect 9088 19007 9404 19008
rect 14516 19072 14832 19073
rect 14516 19008 14522 19072
rect 14586 19008 14602 19072
rect 14666 19008 14682 19072
rect 14746 19008 14762 19072
rect 14826 19008 14832 19072
rect 14516 19007 14832 19008
rect 19944 19072 20260 19073
rect 19944 19008 19950 19072
rect 20014 19008 20030 19072
rect 20094 19008 20110 19072
rect 20174 19008 20190 19072
rect 20254 19008 20260 19072
rect 19944 19007 20260 19008
rect 6374 18528 6690 18529
rect 6374 18464 6380 18528
rect 6444 18464 6460 18528
rect 6524 18464 6540 18528
rect 6604 18464 6620 18528
rect 6684 18464 6690 18528
rect 6374 18463 6690 18464
rect 11802 18528 12118 18529
rect 11802 18464 11808 18528
rect 11872 18464 11888 18528
rect 11952 18464 11968 18528
rect 12032 18464 12048 18528
rect 12112 18464 12118 18528
rect 11802 18463 12118 18464
rect 17230 18528 17546 18529
rect 17230 18464 17236 18528
rect 17300 18464 17316 18528
rect 17380 18464 17396 18528
rect 17460 18464 17476 18528
rect 17540 18464 17546 18528
rect 17230 18463 17546 18464
rect 22658 18528 22974 18529
rect 22658 18464 22664 18528
rect 22728 18464 22744 18528
rect 22808 18464 22824 18528
rect 22888 18464 22904 18528
rect 22968 18464 22974 18528
rect 22658 18463 22974 18464
rect 3660 17984 3976 17985
rect 3660 17920 3666 17984
rect 3730 17920 3746 17984
rect 3810 17920 3826 17984
rect 3890 17920 3906 17984
rect 3970 17920 3976 17984
rect 3660 17919 3976 17920
rect 9088 17984 9404 17985
rect 9088 17920 9094 17984
rect 9158 17920 9174 17984
rect 9238 17920 9254 17984
rect 9318 17920 9334 17984
rect 9398 17920 9404 17984
rect 9088 17919 9404 17920
rect 14516 17984 14832 17985
rect 14516 17920 14522 17984
rect 14586 17920 14602 17984
rect 14666 17920 14682 17984
rect 14746 17920 14762 17984
rect 14826 17920 14832 17984
rect 14516 17919 14832 17920
rect 19944 17984 20260 17985
rect 19944 17920 19950 17984
rect 20014 17920 20030 17984
rect 20094 17920 20110 17984
rect 20174 17920 20190 17984
rect 20254 17920 20260 17984
rect 19944 17919 20260 17920
rect 6374 17440 6690 17441
rect 6374 17376 6380 17440
rect 6444 17376 6460 17440
rect 6524 17376 6540 17440
rect 6604 17376 6620 17440
rect 6684 17376 6690 17440
rect 6374 17375 6690 17376
rect 11802 17440 12118 17441
rect 11802 17376 11808 17440
rect 11872 17376 11888 17440
rect 11952 17376 11968 17440
rect 12032 17376 12048 17440
rect 12112 17376 12118 17440
rect 11802 17375 12118 17376
rect 17230 17440 17546 17441
rect 17230 17376 17236 17440
rect 17300 17376 17316 17440
rect 17380 17376 17396 17440
rect 17460 17376 17476 17440
rect 17540 17376 17546 17440
rect 17230 17375 17546 17376
rect 22658 17440 22974 17441
rect 22658 17376 22664 17440
rect 22728 17376 22744 17440
rect 22808 17376 22824 17440
rect 22888 17376 22904 17440
rect 22968 17376 22974 17440
rect 22658 17375 22974 17376
rect 3660 16896 3976 16897
rect 3660 16832 3666 16896
rect 3730 16832 3746 16896
rect 3810 16832 3826 16896
rect 3890 16832 3906 16896
rect 3970 16832 3976 16896
rect 3660 16831 3976 16832
rect 9088 16896 9404 16897
rect 9088 16832 9094 16896
rect 9158 16832 9174 16896
rect 9238 16832 9254 16896
rect 9318 16832 9334 16896
rect 9398 16832 9404 16896
rect 9088 16831 9404 16832
rect 14516 16896 14832 16897
rect 14516 16832 14522 16896
rect 14586 16832 14602 16896
rect 14666 16832 14682 16896
rect 14746 16832 14762 16896
rect 14826 16832 14832 16896
rect 14516 16831 14832 16832
rect 19944 16896 20260 16897
rect 19944 16832 19950 16896
rect 20014 16832 20030 16896
rect 20094 16832 20110 16896
rect 20174 16832 20190 16896
rect 20254 16832 20260 16896
rect 19944 16831 20260 16832
rect 6374 16352 6690 16353
rect 6374 16288 6380 16352
rect 6444 16288 6460 16352
rect 6524 16288 6540 16352
rect 6604 16288 6620 16352
rect 6684 16288 6690 16352
rect 6374 16287 6690 16288
rect 11802 16352 12118 16353
rect 11802 16288 11808 16352
rect 11872 16288 11888 16352
rect 11952 16288 11968 16352
rect 12032 16288 12048 16352
rect 12112 16288 12118 16352
rect 11802 16287 12118 16288
rect 17230 16352 17546 16353
rect 17230 16288 17236 16352
rect 17300 16288 17316 16352
rect 17380 16288 17396 16352
rect 17460 16288 17476 16352
rect 17540 16288 17546 16352
rect 17230 16287 17546 16288
rect 22658 16352 22974 16353
rect 22658 16288 22664 16352
rect 22728 16288 22744 16352
rect 22808 16288 22824 16352
rect 22888 16288 22904 16352
rect 22968 16288 22974 16352
rect 22658 16287 22974 16288
rect 3660 15808 3976 15809
rect 3660 15744 3666 15808
rect 3730 15744 3746 15808
rect 3810 15744 3826 15808
rect 3890 15744 3906 15808
rect 3970 15744 3976 15808
rect 3660 15743 3976 15744
rect 9088 15808 9404 15809
rect 9088 15744 9094 15808
rect 9158 15744 9174 15808
rect 9238 15744 9254 15808
rect 9318 15744 9334 15808
rect 9398 15744 9404 15808
rect 9088 15743 9404 15744
rect 14516 15808 14832 15809
rect 14516 15744 14522 15808
rect 14586 15744 14602 15808
rect 14666 15744 14682 15808
rect 14746 15744 14762 15808
rect 14826 15744 14832 15808
rect 14516 15743 14832 15744
rect 19944 15808 20260 15809
rect 19944 15744 19950 15808
rect 20014 15744 20030 15808
rect 20094 15744 20110 15808
rect 20174 15744 20190 15808
rect 20254 15744 20260 15808
rect 19944 15743 20260 15744
rect 6374 15264 6690 15265
rect 6374 15200 6380 15264
rect 6444 15200 6460 15264
rect 6524 15200 6540 15264
rect 6604 15200 6620 15264
rect 6684 15200 6690 15264
rect 6374 15199 6690 15200
rect 11802 15264 12118 15265
rect 11802 15200 11808 15264
rect 11872 15200 11888 15264
rect 11952 15200 11968 15264
rect 12032 15200 12048 15264
rect 12112 15200 12118 15264
rect 11802 15199 12118 15200
rect 17230 15264 17546 15265
rect 17230 15200 17236 15264
rect 17300 15200 17316 15264
rect 17380 15200 17396 15264
rect 17460 15200 17476 15264
rect 17540 15200 17546 15264
rect 17230 15199 17546 15200
rect 22658 15264 22974 15265
rect 22658 15200 22664 15264
rect 22728 15200 22744 15264
rect 22808 15200 22824 15264
rect 22888 15200 22904 15264
rect 22968 15200 22974 15264
rect 22658 15199 22974 15200
rect 3660 14720 3976 14721
rect 3660 14656 3666 14720
rect 3730 14656 3746 14720
rect 3810 14656 3826 14720
rect 3890 14656 3906 14720
rect 3970 14656 3976 14720
rect 3660 14655 3976 14656
rect 9088 14720 9404 14721
rect 9088 14656 9094 14720
rect 9158 14656 9174 14720
rect 9238 14656 9254 14720
rect 9318 14656 9334 14720
rect 9398 14656 9404 14720
rect 9088 14655 9404 14656
rect 14516 14720 14832 14721
rect 14516 14656 14522 14720
rect 14586 14656 14602 14720
rect 14666 14656 14682 14720
rect 14746 14656 14762 14720
rect 14826 14656 14832 14720
rect 14516 14655 14832 14656
rect 19944 14720 20260 14721
rect 19944 14656 19950 14720
rect 20014 14656 20030 14720
rect 20094 14656 20110 14720
rect 20174 14656 20190 14720
rect 20254 14656 20260 14720
rect 19944 14655 20260 14656
rect 6374 14176 6690 14177
rect 6374 14112 6380 14176
rect 6444 14112 6460 14176
rect 6524 14112 6540 14176
rect 6604 14112 6620 14176
rect 6684 14112 6690 14176
rect 6374 14111 6690 14112
rect 11802 14176 12118 14177
rect 11802 14112 11808 14176
rect 11872 14112 11888 14176
rect 11952 14112 11968 14176
rect 12032 14112 12048 14176
rect 12112 14112 12118 14176
rect 11802 14111 12118 14112
rect 17230 14176 17546 14177
rect 17230 14112 17236 14176
rect 17300 14112 17316 14176
rect 17380 14112 17396 14176
rect 17460 14112 17476 14176
rect 17540 14112 17546 14176
rect 17230 14111 17546 14112
rect 22658 14176 22974 14177
rect 22658 14112 22664 14176
rect 22728 14112 22744 14176
rect 22808 14112 22824 14176
rect 22888 14112 22904 14176
rect 22968 14112 22974 14176
rect 22658 14111 22974 14112
rect 3660 13632 3976 13633
rect 3660 13568 3666 13632
rect 3730 13568 3746 13632
rect 3810 13568 3826 13632
rect 3890 13568 3906 13632
rect 3970 13568 3976 13632
rect 3660 13567 3976 13568
rect 9088 13632 9404 13633
rect 9088 13568 9094 13632
rect 9158 13568 9174 13632
rect 9238 13568 9254 13632
rect 9318 13568 9334 13632
rect 9398 13568 9404 13632
rect 9088 13567 9404 13568
rect 14516 13632 14832 13633
rect 14516 13568 14522 13632
rect 14586 13568 14602 13632
rect 14666 13568 14682 13632
rect 14746 13568 14762 13632
rect 14826 13568 14832 13632
rect 14516 13567 14832 13568
rect 19944 13632 20260 13633
rect 19944 13568 19950 13632
rect 20014 13568 20030 13632
rect 20094 13568 20110 13632
rect 20174 13568 20190 13632
rect 20254 13568 20260 13632
rect 19944 13567 20260 13568
rect 6374 13088 6690 13089
rect 6374 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6690 13088
rect 6374 13023 6690 13024
rect 11802 13088 12118 13089
rect 11802 13024 11808 13088
rect 11872 13024 11888 13088
rect 11952 13024 11968 13088
rect 12032 13024 12048 13088
rect 12112 13024 12118 13088
rect 11802 13023 12118 13024
rect 17230 13088 17546 13089
rect 17230 13024 17236 13088
rect 17300 13024 17316 13088
rect 17380 13024 17396 13088
rect 17460 13024 17476 13088
rect 17540 13024 17546 13088
rect 17230 13023 17546 13024
rect 22658 13088 22974 13089
rect 22658 13024 22664 13088
rect 22728 13024 22744 13088
rect 22808 13024 22824 13088
rect 22888 13024 22904 13088
rect 22968 13024 22974 13088
rect 22658 13023 22974 13024
rect 3660 12544 3976 12545
rect 3660 12480 3666 12544
rect 3730 12480 3746 12544
rect 3810 12480 3826 12544
rect 3890 12480 3906 12544
rect 3970 12480 3976 12544
rect 3660 12479 3976 12480
rect 9088 12544 9404 12545
rect 9088 12480 9094 12544
rect 9158 12480 9174 12544
rect 9238 12480 9254 12544
rect 9318 12480 9334 12544
rect 9398 12480 9404 12544
rect 9088 12479 9404 12480
rect 14516 12544 14832 12545
rect 14516 12480 14522 12544
rect 14586 12480 14602 12544
rect 14666 12480 14682 12544
rect 14746 12480 14762 12544
rect 14826 12480 14832 12544
rect 14516 12479 14832 12480
rect 19944 12544 20260 12545
rect 19944 12480 19950 12544
rect 20014 12480 20030 12544
rect 20094 12480 20110 12544
rect 20174 12480 20190 12544
rect 20254 12480 20260 12544
rect 19944 12479 20260 12480
rect 5717 12474 5783 12477
rect 5901 12474 5967 12477
rect 5717 12472 5967 12474
rect 5717 12416 5722 12472
rect 5778 12416 5906 12472
rect 5962 12416 5967 12472
rect 5717 12414 5967 12416
rect 5717 12411 5783 12414
rect 5901 12411 5967 12414
rect 6374 12000 6690 12001
rect 6374 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6690 12000
rect 6374 11935 6690 11936
rect 11802 12000 12118 12001
rect 11802 11936 11808 12000
rect 11872 11936 11888 12000
rect 11952 11936 11968 12000
rect 12032 11936 12048 12000
rect 12112 11936 12118 12000
rect 11802 11935 12118 11936
rect 17230 12000 17546 12001
rect 17230 11936 17236 12000
rect 17300 11936 17316 12000
rect 17380 11936 17396 12000
rect 17460 11936 17476 12000
rect 17540 11936 17546 12000
rect 17230 11935 17546 11936
rect 22658 12000 22974 12001
rect 22658 11936 22664 12000
rect 22728 11936 22744 12000
rect 22808 11936 22824 12000
rect 22888 11936 22904 12000
rect 22968 11936 22974 12000
rect 22658 11935 22974 11936
rect 3660 11456 3976 11457
rect 3660 11392 3666 11456
rect 3730 11392 3746 11456
rect 3810 11392 3826 11456
rect 3890 11392 3906 11456
rect 3970 11392 3976 11456
rect 3660 11391 3976 11392
rect 9088 11456 9404 11457
rect 9088 11392 9094 11456
rect 9158 11392 9174 11456
rect 9238 11392 9254 11456
rect 9318 11392 9334 11456
rect 9398 11392 9404 11456
rect 9088 11391 9404 11392
rect 14516 11456 14832 11457
rect 14516 11392 14522 11456
rect 14586 11392 14602 11456
rect 14666 11392 14682 11456
rect 14746 11392 14762 11456
rect 14826 11392 14832 11456
rect 14516 11391 14832 11392
rect 19944 11456 20260 11457
rect 19944 11392 19950 11456
rect 20014 11392 20030 11456
rect 20094 11392 20110 11456
rect 20174 11392 20190 11456
rect 20254 11392 20260 11456
rect 19944 11391 20260 11392
rect 6374 10912 6690 10913
rect 6374 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6690 10912
rect 6374 10847 6690 10848
rect 11802 10912 12118 10913
rect 11802 10848 11808 10912
rect 11872 10848 11888 10912
rect 11952 10848 11968 10912
rect 12032 10848 12048 10912
rect 12112 10848 12118 10912
rect 11802 10847 12118 10848
rect 17230 10912 17546 10913
rect 17230 10848 17236 10912
rect 17300 10848 17316 10912
rect 17380 10848 17396 10912
rect 17460 10848 17476 10912
rect 17540 10848 17546 10912
rect 17230 10847 17546 10848
rect 22658 10912 22974 10913
rect 22658 10848 22664 10912
rect 22728 10848 22744 10912
rect 22808 10848 22824 10912
rect 22888 10848 22904 10912
rect 22968 10848 22974 10912
rect 22658 10847 22974 10848
rect 9673 10706 9739 10709
rect 18229 10706 18295 10709
rect 9673 10704 18295 10706
rect 9673 10648 9678 10704
rect 9734 10648 18234 10704
rect 18290 10648 18295 10704
rect 9673 10646 18295 10648
rect 9673 10643 9739 10646
rect 18229 10643 18295 10646
rect 5901 10570 5967 10573
rect 6269 10570 6335 10573
rect 5901 10568 6335 10570
rect 5901 10512 5906 10568
rect 5962 10512 6274 10568
rect 6330 10512 6335 10568
rect 5901 10510 6335 10512
rect 5901 10507 5967 10510
rect 6269 10507 6335 10510
rect 3660 10368 3976 10369
rect 3660 10304 3666 10368
rect 3730 10304 3746 10368
rect 3810 10304 3826 10368
rect 3890 10304 3906 10368
rect 3970 10304 3976 10368
rect 3660 10303 3976 10304
rect 9088 10368 9404 10369
rect 9088 10304 9094 10368
rect 9158 10304 9174 10368
rect 9238 10304 9254 10368
rect 9318 10304 9334 10368
rect 9398 10304 9404 10368
rect 9088 10303 9404 10304
rect 14516 10368 14832 10369
rect 14516 10304 14522 10368
rect 14586 10304 14602 10368
rect 14666 10304 14682 10368
rect 14746 10304 14762 10368
rect 14826 10304 14832 10368
rect 14516 10303 14832 10304
rect 19944 10368 20260 10369
rect 19944 10304 19950 10368
rect 20014 10304 20030 10368
rect 20094 10304 20110 10368
rect 20174 10304 20190 10368
rect 20254 10304 20260 10368
rect 19944 10303 20260 10304
rect 4705 10026 4771 10029
rect 18413 10026 18479 10029
rect 4705 10024 18479 10026
rect 4705 9968 4710 10024
rect 4766 9968 18418 10024
rect 18474 9968 18479 10024
rect 4705 9966 18479 9968
rect 4705 9963 4771 9966
rect 18413 9963 18479 9966
rect 6374 9824 6690 9825
rect 6374 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6690 9824
rect 6374 9759 6690 9760
rect 11802 9824 12118 9825
rect 11802 9760 11808 9824
rect 11872 9760 11888 9824
rect 11952 9760 11968 9824
rect 12032 9760 12048 9824
rect 12112 9760 12118 9824
rect 11802 9759 12118 9760
rect 17230 9824 17546 9825
rect 17230 9760 17236 9824
rect 17300 9760 17316 9824
rect 17380 9760 17396 9824
rect 17460 9760 17476 9824
rect 17540 9760 17546 9824
rect 17230 9759 17546 9760
rect 22658 9824 22974 9825
rect 22658 9760 22664 9824
rect 22728 9760 22744 9824
rect 22808 9760 22824 9824
rect 22888 9760 22904 9824
rect 22968 9760 22974 9824
rect 22658 9759 22974 9760
rect 3660 9280 3976 9281
rect 3660 9216 3666 9280
rect 3730 9216 3746 9280
rect 3810 9216 3826 9280
rect 3890 9216 3906 9280
rect 3970 9216 3976 9280
rect 3660 9215 3976 9216
rect 9088 9280 9404 9281
rect 9088 9216 9094 9280
rect 9158 9216 9174 9280
rect 9238 9216 9254 9280
rect 9318 9216 9334 9280
rect 9398 9216 9404 9280
rect 9088 9215 9404 9216
rect 14516 9280 14832 9281
rect 14516 9216 14522 9280
rect 14586 9216 14602 9280
rect 14666 9216 14682 9280
rect 14746 9216 14762 9280
rect 14826 9216 14832 9280
rect 14516 9215 14832 9216
rect 19944 9280 20260 9281
rect 19944 9216 19950 9280
rect 20014 9216 20030 9280
rect 20094 9216 20110 9280
rect 20174 9216 20190 9280
rect 20254 9216 20260 9280
rect 19944 9215 20260 9216
rect 6374 8736 6690 8737
rect 6374 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6690 8736
rect 6374 8671 6690 8672
rect 11802 8736 12118 8737
rect 11802 8672 11808 8736
rect 11872 8672 11888 8736
rect 11952 8672 11968 8736
rect 12032 8672 12048 8736
rect 12112 8672 12118 8736
rect 11802 8671 12118 8672
rect 17230 8736 17546 8737
rect 17230 8672 17236 8736
rect 17300 8672 17316 8736
rect 17380 8672 17396 8736
rect 17460 8672 17476 8736
rect 17540 8672 17546 8736
rect 17230 8671 17546 8672
rect 22658 8736 22974 8737
rect 22658 8672 22664 8736
rect 22728 8672 22744 8736
rect 22808 8672 22824 8736
rect 22888 8672 22904 8736
rect 22968 8672 22974 8736
rect 22658 8671 22974 8672
rect 3660 8192 3976 8193
rect 3660 8128 3666 8192
rect 3730 8128 3746 8192
rect 3810 8128 3826 8192
rect 3890 8128 3906 8192
rect 3970 8128 3976 8192
rect 3660 8127 3976 8128
rect 9088 8192 9404 8193
rect 9088 8128 9094 8192
rect 9158 8128 9174 8192
rect 9238 8128 9254 8192
rect 9318 8128 9334 8192
rect 9398 8128 9404 8192
rect 9088 8127 9404 8128
rect 14516 8192 14832 8193
rect 14516 8128 14522 8192
rect 14586 8128 14602 8192
rect 14666 8128 14682 8192
rect 14746 8128 14762 8192
rect 14826 8128 14832 8192
rect 14516 8127 14832 8128
rect 19944 8192 20260 8193
rect 19944 8128 19950 8192
rect 20014 8128 20030 8192
rect 20094 8128 20110 8192
rect 20174 8128 20190 8192
rect 20254 8128 20260 8192
rect 19944 8127 20260 8128
rect 7005 7986 7071 7989
rect 16941 7986 17007 7989
rect 7005 7984 17007 7986
rect 7005 7928 7010 7984
rect 7066 7928 16946 7984
rect 17002 7928 17007 7984
rect 7005 7926 17007 7928
rect 7005 7923 7071 7926
rect 16941 7923 17007 7926
rect 6374 7648 6690 7649
rect 6374 7584 6380 7648
rect 6444 7584 6460 7648
rect 6524 7584 6540 7648
rect 6604 7584 6620 7648
rect 6684 7584 6690 7648
rect 6374 7583 6690 7584
rect 11802 7648 12118 7649
rect 11802 7584 11808 7648
rect 11872 7584 11888 7648
rect 11952 7584 11968 7648
rect 12032 7584 12048 7648
rect 12112 7584 12118 7648
rect 11802 7583 12118 7584
rect 17230 7648 17546 7649
rect 17230 7584 17236 7648
rect 17300 7584 17316 7648
rect 17380 7584 17396 7648
rect 17460 7584 17476 7648
rect 17540 7584 17546 7648
rect 17230 7583 17546 7584
rect 22658 7648 22974 7649
rect 22658 7584 22664 7648
rect 22728 7584 22744 7648
rect 22808 7584 22824 7648
rect 22888 7584 22904 7648
rect 22968 7584 22974 7648
rect 22658 7583 22974 7584
rect 3660 7104 3976 7105
rect 3660 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3976 7104
rect 3660 7039 3976 7040
rect 9088 7104 9404 7105
rect 9088 7040 9094 7104
rect 9158 7040 9174 7104
rect 9238 7040 9254 7104
rect 9318 7040 9334 7104
rect 9398 7040 9404 7104
rect 9088 7039 9404 7040
rect 14516 7104 14832 7105
rect 14516 7040 14522 7104
rect 14586 7040 14602 7104
rect 14666 7040 14682 7104
rect 14746 7040 14762 7104
rect 14826 7040 14832 7104
rect 14516 7039 14832 7040
rect 19944 7104 20260 7105
rect 19944 7040 19950 7104
rect 20014 7040 20030 7104
rect 20094 7040 20110 7104
rect 20174 7040 20190 7104
rect 20254 7040 20260 7104
rect 19944 7039 20260 7040
rect 6374 6560 6690 6561
rect 6374 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6690 6560
rect 6374 6495 6690 6496
rect 11802 6560 12118 6561
rect 11802 6496 11808 6560
rect 11872 6496 11888 6560
rect 11952 6496 11968 6560
rect 12032 6496 12048 6560
rect 12112 6496 12118 6560
rect 11802 6495 12118 6496
rect 17230 6560 17546 6561
rect 17230 6496 17236 6560
rect 17300 6496 17316 6560
rect 17380 6496 17396 6560
rect 17460 6496 17476 6560
rect 17540 6496 17546 6560
rect 17230 6495 17546 6496
rect 22658 6560 22974 6561
rect 22658 6496 22664 6560
rect 22728 6496 22744 6560
rect 22808 6496 22824 6560
rect 22888 6496 22904 6560
rect 22968 6496 22974 6560
rect 22658 6495 22974 6496
rect 3660 6016 3976 6017
rect 3660 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3976 6016
rect 3660 5951 3976 5952
rect 9088 6016 9404 6017
rect 9088 5952 9094 6016
rect 9158 5952 9174 6016
rect 9238 5952 9254 6016
rect 9318 5952 9334 6016
rect 9398 5952 9404 6016
rect 9088 5951 9404 5952
rect 14516 6016 14832 6017
rect 14516 5952 14522 6016
rect 14586 5952 14602 6016
rect 14666 5952 14682 6016
rect 14746 5952 14762 6016
rect 14826 5952 14832 6016
rect 14516 5951 14832 5952
rect 19944 6016 20260 6017
rect 19944 5952 19950 6016
rect 20014 5952 20030 6016
rect 20094 5952 20110 6016
rect 20174 5952 20190 6016
rect 20254 5952 20260 6016
rect 19944 5951 20260 5952
rect 6374 5472 6690 5473
rect 6374 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6690 5472
rect 6374 5407 6690 5408
rect 11802 5472 12118 5473
rect 11802 5408 11808 5472
rect 11872 5408 11888 5472
rect 11952 5408 11968 5472
rect 12032 5408 12048 5472
rect 12112 5408 12118 5472
rect 11802 5407 12118 5408
rect 17230 5472 17546 5473
rect 17230 5408 17236 5472
rect 17300 5408 17316 5472
rect 17380 5408 17396 5472
rect 17460 5408 17476 5472
rect 17540 5408 17546 5472
rect 17230 5407 17546 5408
rect 22658 5472 22974 5473
rect 22658 5408 22664 5472
rect 22728 5408 22744 5472
rect 22808 5408 22824 5472
rect 22888 5408 22904 5472
rect 22968 5408 22974 5472
rect 22658 5407 22974 5408
rect 3660 4928 3976 4929
rect 3660 4864 3666 4928
rect 3730 4864 3746 4928
rect 3810 4864 3826 4928
rect 3890 4864 3906 4928
rect 3970 4864 3976 4928
rect 3660 4863 3976 4864
rect 9088 4928 9404 4929
rect 9088 4864 9094 4928
rect 9158 4864 9174 4928
rect 9238 4864 9254 4928
rect 9318 4864 9334 4928
rect 9398 4864 9404 4928
rect 9088 4863 9404 4864
rect 14516 4928 14832 4929
rect 14516 4864 14522 4928
rect 14586 4864 14602 4928
rect 14666 4864 14682 4928
rect 14746 4864 14762 4928
rect 14826 4864 14832 4928
rect 14516 4863 14832 4864
rect 19944 4928 20260 4929
rect 19944 4864 19950 4928
rect 20014 4864 20030 4928
rect 20094 4864 20110 4928
rect 20174 4864 20190 4928
rect 20254 4864 20260 4928
rect 19944 4863 20260 4864
rect 6374 4384 6690 4385
rect 6374 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6690 4384
rect 6374 4319 6690 4320
rect 11802 4384 12118 4385
rect 11802 4320 11808 4384
rect 11872 4320 11888 4384
rect 11952 4320 11968 4384
rect 12032 4320 12048 4384
rect 12112 4320 12118 4384
rect 11802 4319 12118 4320
rect 17230 4384 17546 4385
rect 17230 4320 17236 4384
rect 17300 4320 17316 4384
rect 17380 4320 17396 4384
rect 17460 4320 17476 4384
rect 17540 4320 17546 4384
rect 17230 4319 17546 4320
rect 22658 4384 22974 4385
rect 22658 4320 22664 4384
rect 22728 4320 22744 4384
rect 22808 4320 22824 4384
rect 22888 4320 22904 4384
rect 22968 4320 22974 4384
rect 22658 4319 22974 4320
rect 3660 3840 3976 3841
rect 3660 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3976 3840
rect 3660 3775 3976 3776
rect 9088 3840 9404 3841
rect 9088 3776 9094 3840
rect 9158 3776 9174 3840
rect 9238 3776 9254 3840
rect 9318 3776 9334 3840
rect 9398 3776 9404 3840
rect 9088 3775 9404 3776
rect 14516 3840 14832 3841
rect 14516 3776 14522 3840
rect 14586 3776 14602 3840
rect 14666 3776 14682 3840
rect 14746 3776 14762 3840
rect 14826 3776 14832 3840
rect 14516 3775 14832 3776
rect 19944 3840 20260 3841
rect 19944 3776 19950 3840
rect 20014 3776 20030 3840
rect 20094 3776 20110 3840
rect 20174 3776 20190 3840
rect 20254 3776 20260 3840
rect 19944 3775 20260 3776
rect 6374 3296 6690 3297
rect 6374 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6690 3296
rect 6374 3231 6690 3232
rect 11802 3296 12118 3297
rect 11802 3232 11808 3296
rect 11872 3232 11888 3296
rect 11952 3232 11968 3296
rect 12032 3232 12048 3296
rect 12112 3232 12118 3296
rect 11802 3231 12118 3232
rect 17230 3296 17546 3297
rect 17230 3232 17236 3296
rect 17300 3232 17316 3296
rect 17380 3232 17396 3296
rect 17460 3232 17476 3296
rect 17540 3232 17546 3296
rect 17230 3231 17546 3232
rect 22658 3296 22974 3297
rect 22658 3232 22664 3296
rect 22728 3232 22744 3296
rect 22808 3232 22824 3296
rect 22888 3232 22904 3296
rect 22968 3232 22974 3296
rect 22658 3231 22974 3232
rect 3660 2752 3976 2753
rect 3660 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3976 2752
rect 3660 2687 3976 2688
rect 9088 2752 9404 2753
rect 9088 2688 9094 2752
rect 9158 2688 9174 2752
rect 9238 2688 9254 2752
rect 9318 2688 9334 2752
rect 9398 2688 9404 2752
rect 9088 2687 9404 2688
rect 14516 2752 14832 2753
rect 14516 2688 14522 2752
rect 14586 2688 14602 2752
rect 14666 2688 14682 2752
rect 14746 2688 14762 2752
rect 14826 2688 14832 2752
rect 14516 2687 14832 2688
rect 19944 2752 20260 2753
rect 19944 2688 19950 2752
rect 20014 2688 20030 2752
rect 20094 2688 20110 2752
rect 20174 2688 20190 2752
rect 20254 2688 20260 2752
rect 19944 2687 20260 2688
rect 6374 2208 6690 2209
rect 6374 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6690 2208
rect 6374 2143 6690 2144
rect 11802 2208 12118 2209
rect 11802 2144 11808 2208
rect 11872 2144 11888 2208
rect 11952 2144 11968 2208
rect 12032 2144 12048 2208
rect 12112 2144 12118 2208
rect 11802 2143 12118 2144
rect 17230 2208 17546 2209
rect 17230 2144 17236 2208
rect 17300 2144 17316 2208
rect 17380 2144 17396 2208
rect 17460 2144 17476 2208
rect 17540 2144 17546 2208
rect 17230 2143 17546 2144
rect 22658 2208 22974 2209
rect 22658 2144 22664 2208
rect 22728 2144 22744 2208
rect 22808 2144 22824 2208
rect 22888 2144 22904 2208
rect 22968 2144 22974 2208
rect 22658 2143 22974 2144
<< via3 >>
rect 6380 21788 6444 21792
rect 6380 21732 6384 21788
rect 6384 21732 6440 21788
rect 6440 21732 6444 21788
rect 6380 21728 6444 21732
rect 6460 21788 6524 21792
rect 6460 21732 6464 21788
rect 6464 21732 6520 21788
rect 6520 21732 6524 21788
rect 6460 21728 6524 21732
rect 6540 21788 6604 21792
rect 6540 21732 6544 21788
rect 6544 21732 6600 21788
rect 6600 21732 6604 21788
rect 6540 21728 6604 21732
rect 6620 21788 6684 21792
rect 6620 21732 6624 21788
rect 6624 21732 6680 21788
rect 6680 21732 6684 21788
rect 6620 21728 6684 21732
rect 11808 21788 11872 21792
rect 11808 21732 11812 21788
rect 11812 21732 11868 21788
rect 11868 21732 11872 21788
rect 11808 21728 11872 21732
rect 11888 21788 11952 21792
rect 11888 21732 11892 21788
rect 11892 21732 11948 21788
rect 11948 21732 11952 21788
rect 11888 21728 11952 21732
rect 11968 21788 12032 21792
rect 11968 21732 11972 21788
rect 11972 21732 12028 21788
rect 12028 21732 12032 21788
rect 11968 21728 12032 21732
rect 12048 21788 12112 21792
rect 12048 21732 12052 21788
rect 12052 21732 12108 21788
rect 12108 21732 12112 21788
rect 12048 21728 12112 21732
rect 17236 21788 17300 21792
rect 17236 21732 17240 21788
rect 17240 21732 17296 21788
rect 17296 21732 17300 21788
rect 17236 21728 17300 21732
rect 17316 21788 17380 21792
rect 17316 21732 17320 21788
rect 17320 21732 17376 21788
rect 17376 21732 17380 21788
rect 17316 21728 17380 21732
rect 17396 21788 17460 21792
rect 17396 21732 17400 21788
rect 17400 21732 17456 21788
rect 17456 21732 17460 21788
rect 17396 21728 17460 21732
rect 17476 21788 17540 21792
rect 17476 21732 17480 21788
rect 17480 21732 17536 21788
rect 17536 21732 17540 21788
rect 17476 21728 17540 21732
rect 22664 21788 22728 21792
rect 22664 21732 22668 21788
rect 22668 21732 22724 21788
rect 22724 21732 22728 21788
rect 22664 21728 22728 21732
rect 22744 21788 22808 21792
rect 22744 21732 22748 21788
rect 22748 21732 22804 21788
rect 22804 21732 22808 21788
rect 22744 21728 22808 21732
rect 22824 21788 22888 21792
rect 22824 21732 22828 21788
rect 22828 21732 22884 21788
rect 22884 21732 22888 21788
rect 22824 21728 22888 21732
rect 22904 21788 22968 21792
rect 22904 21732 22908 21788
rect 22908 21732 22964 21788
rect 22964 21732 22968 21788
rect 22904 21728 22968 21732
rect 3666 21244 3730 21248
rect 3666 21188 3670 21244
rect 3670 21188 3726 21244
rect 3726 21188 3730 21244
rect 3666 21184 3730 21188
rect 3746 21244 3810 21248
rect 3746 21188 3750 21244
rect 3750 21188 3806 21244
rect 3806 21188 3810 21244
rect 3746 21184 3810 21188
rect 3826 21244 3890 21248
rect 3826 21188 3830 21244
rect 3830 21188 3886 21244
rect 3886 21188 3890 21244
rect 3826 21184 3890 21188
rect 3906 21244 3970 21248
rect 3906 21188 3910 21244
rect 3910 21188 3966 21244
rect 3966 21188 3970 21244
rect 3906 21184 3970 21188
rect 9094 21244 9158 21248
rect 9094 21188 9098 21244
rect 9098 21188 9154 21244
rect 9154 21188 9158 21244
rect 9094 21184 9158 21188
rect 9174 21244 9238 21248
rect 9174 21188 9178 21244
rect 9178 21188 9234 21244
rect 9234 21188 9238 21244
rect 9174 21184 9238 21188
rect 9254 21244 9318 21248
rect 9254 21188 9258 21244
rect 9258 21188 9314 21244
rect 9314 21188 9318 21244
rect 9254 21184 9318 21188
rect 9334 21244 9398 21248
rect 9334 21188 9338 21244
rect 9338 21188 9394 21244
rect 9394 21188 9398 21244
rect 9334 21184 9398 21188
rect 14522 21244 14586 21248
rect 14522 21188 14526 21244
rect 14526 21188 14582 21244
rect 14582 21188 14586 21244
rect 14522 21184 14586 21188
rect 14602 21244 14666 21248
rect 14602 21188 14606 21244
rect 14606 21188 14662 21244
rect 14662 21188 14666 21244
rect 14602 21184 14666 21188
rect 14682 21244 14746 21248
rect 14682 21188 14686 21244
rect 14686 21188 14742 21244
rect 14742 21188 14746 21244
rect 14682 21184 14746 21188
rect 14762 21244 14826 21248
rect 14762 21188 14766 21244
rect 14766 21188 14822 21244
rect 14822 21188 14826 21244
rect 14762 21184 14826 21188
rect 19950 21244 20014 21248
rect 19950 21188 19954 21244
rect 19954 21188 20010 21244
rect 20010 21188 20014 21244
rect 19950 21184 20014 21188
rect 20030 21244 20094 21248
rect 20030 21188 20034 21244
rect 20034 21188 20090 21244
rect 20090 21188 20094 21244
rect 20030 21184 20094 21188
rect 20110 21244 20174 21248
rect 20110 21188 20114 21244
rect 20114 21188 20170 21244
rect 20170 21188 20174 21244
rect 20110 21184 20174 21188
rect 20190 21244 20254 21248
rect 20190 21188 20194 21244
rect 20194 21188 20250 21244
rect 20250 21188 20254 21244
rect 20190 21184 20254 21188
rect 6380 20700 6444 20704
rect 6380 20644 6384 20700
rect 6384 20644 6440 20700
rect 6440 20644 6444 20700
rect 6380 20640 6444 20644
rect 6460 20700 6524 20704
rect 6460 20644 6464 20700
rect 6464 20644 6520 20700
rect 6520 20644 6524 20700
rect 6460 20640 6524 20644
rect 6540 20700 6604 20704
rect 6540 20644 6544 20700
rect 6544 20644 6600 20700
rect 6600 20644 6604 20700
rect 6540 20640 6604 20644
rect 6620 20700 6684 20704
rect 6620 20644 6624 20700
rect 6624 20644 6680 20700
rect 6680 20644 6684 20700
rect 6620 20640 6684 20644
rect 11808 20700 11872 20704
rect 11808 20644 11812 20700
rect 11812 20644 11868 20700
rect 11868 20644 11872 20700
rect 11808 20640 11872 20644
rect 11888 20700 11952 20704
rect 11888 20644 11892 20700
rect 11892 20644 11948 20700
rect 11948 20644 11952 20700
rect 11888 20640 11952 20644
rect 11968 20700 12032 20704
rect 11968 20644 11972 20700
rect 11972 20644 12028 20700
rect 12028 20644 12032 20700
rect 11968 20640 12032 20644
rect 12048 20700 12112 20704
rect 12048 20644 12052 20700
rect 12052 20644 12108 20700
rect 12108 20644 12112 20700
rect 12048 20640 12112 20644
rect 17236 20700 17300 20704
rect 17236 20644 17240 20700
rect 17240 20644 17296 20700
rect 17296 20644 17300 20700
rect 17236 20640 17300 20644
rect 17316 20700 17380 20704
rect 17316 20644 17320 20700
rect 17320 20644 17376 20700
rect 17376 20644 17380 20700
rect 17316 20640 17380 20644
rect 17396 20700 17460 20704
rect 17396 20644 17400 20700
rect 17400 20644 17456 20700
rect 17456 20644 17460 20700
rect 17396 20640 17460 20644
rect 17476 20700 17540 20704
rect 17476 20644 17480 20700
rect 17480 20644 17536 20700
rect 17536 20644 17540 20700
rect 17476 20640 17540 20644
rect 22664 20700 22728 20704
rect 22664 20644 22668 20700
rect 22668 20644 22724 20700
rect 22724 20644 22728 20700
rect 22664 20640 22728 20644
rect 22744 20700 22808 20704
rect 22744 20644 22748 20700
rect 22748 20644 22804 20700
rect 22804 20644 22808 20700
rect 22744 20640 22808 20644
rect 22824 20700 22888 20704
rect 22824 20644 22828 20700
rect 22828 20644 22884 20700
rect 22884 20644 22888 20700
rect 22824 20640 22888 20644
rect 22904 20700 22968 20704
rect 22904 20644 22908 20700
rect 22908 20644 22964 20700
rect 22964 20644 22968 20700
rect 22904 20640 22968 20644
rect 3666 20156 3730 20160
rect 3666 20100 3670 20156
rect 3670 20100 3726 20156
rect 3726 20100 3730 20156
rect 3666 20096 3730 20100
rect 3746 20156 3810 20160
rect 3746 20100 3750 20156
rect 3750 20100 3806 20156
rect 3806 20100 3810 20156
rect 3746 20096 3810 20100
rect 3826 20156 3890 20160
rect 3826 20100 3830 20156
rect 3830 20100 3886 20156
rect 3886 20100 3890 20156
rect 3826 20096 3890 20100
rect 3906 20156 3970 20160
rect 3906 20100 3910 20156
rect 3910 20100 3966 20156
rect 3966 20100 3970 20156
rect 3906 20096 3970 20100
rect 9094 20156 9158 20160
rect 9094 20100 9098 20156
rect 9098 20100 9154 20156
rect 9154 20100 9158 20156
rect 9094 20096 9158 20100
rect 9174 20156 9238 20160
rect 9174 20100 9178 20156
rect 9178 20100 9234 20156
rect 9234 20100 9238 20156
rect 9174 20096 9238 20100
rect 9254 20156 9318 20160
rect 9254 20100 9258 20156
rect 9258 20100 9314 20156
rect 9314 20100 9318 20156
rect 9254 20096 9318 20100
rect 9334 20156 9398 20160
rect 9334 20100 9338 20156
rect 9338 20100 9394 20156
rect 9394 20100 9398 20156
rect 9334 20096 9398 20100
rect 14522 20156 14586 20160
rect 14522 20100 14526 20156
rect 14526 20100 14582 20156
rect 14582 20100 14586 20156
rect 14522 20096 14586 20100
rect 14602 20156 14666 20160
rect 14602 20100 14606 20156
rect 14606 20100 14662 20156
rect 14662 20100 14666 20156
rect 14602 20096 14666 20100
rect 14682 20156 14746 20160
rect 14682 20100 14686 20156
rect 14686 20100 14742 20156
rect 14742 20100 14746 20156
rect 14682 20096 14746 20100
rect 14762 20156 14826 20160
rect 14762 20100 14766 20156
rect 14766 20100 14822 20156
rect 14822 20100 14826 20156
rect 14762 20096 14826 20100
rect 19950 20156 20014 20160
rect 19950 20100 19954 20156
rect 19954 20100 20010 20156
rect 20010 20100 20014 20156
rect 19950 20096 20014 20100
rect 20030 20156 20094 20160
rect 20030 20100 20034 20156
rect 20034 20100 20090 20156
rect 20090 20100 20094 20156
rect 20030 20096 20094 20100
rect 20110 20156 20174 20160
rect 20110 20100 20114 20156
rect 20114 20100 20170 20156
rect 20170 20100 20174 20156
rect 20110 20096 20174 20100
rect 20190 20156 20254 20160
rect 20190 20100 20194 20156
rect 20194 20100 20250 20156
rect 20250 20100 20254 20156
rect 20190 20096 20254 20100
rect 6380 19612 6444 19616
rect 6380 19556 6384 19612
rect 6384 19556 6440 19612
rect 6440 19556 6444 19612
rect 6380 19552 6444 19556
rect 6460 19612 6524 19616
rect 6460 19556 6464 19612
rect 6464 19556 6520 19612
rect 6520 19556 6524 19612
rect 6460 19552 6524 19556
rect 6540 19612 6604 19616
rect 6540 19556 6544 19612
rect 6544 19556 6600 19612
rect 6600 19556 6604 19612
rect 6540 19552 6604 19556
rect 6620 19612 6684 19616
rect 6620 19556 6624 19612
rect 6624 19556 6680 19612
rect 6680 19556 6684 19612
rect 6620 19552 6684 19556
rect 11808 19612 11872 19616
rect 11808 19556 11812 19612
rect 11812 19556 11868 19612
rect 11868 19556 11872 19612
rect 11808 19552 11872 19556
rect 11888 19612 11952 19616
rect 11888 19556 11892 19612
rect 11892 19556 11948 19612
rect 11948 19556 11952 19612
rect 11888 19552 11952 19556
rect 11968 19612 12032 19616
rect 11968 19556 11972 19612
rect 11972 19556 12028 19612
rect 12028 19556 12032 19612
rect 11968 19552 12032 19556
rect 12048 19612 12112 19616
rect 12048 19556 12052 19612
rect 12052 19556 12108 19612
rect 12108 19556 12112 19612
rect 12048 19552 12112 19556
rect 17236 19612 17300 19616
rect 17236 19556 17240 19612
rect 17240 19556 17296 19612
rect 17296 19556 17300 19612
rect 17236 19552 17300 19556
rect 17316 19612 17380 19616
rect 17316 19556 17320 19612
rect 17320 19556 17376 19612
rect 17376 19556 17380 19612
rect 17316 19552 17380 19556
rect 17396 19612 17460 19616
rect 17396 19556 17400 19612
rect 17400 19556 17456 19612
rect 17456 19556 17460 19612
rect 17396 19552 17460 19556
rect 17476 19612 17540 19616
rect 17476 19556 17480 19612
rect 17480 19556 17536 19612
rect 17536 19556 17540 19612
rect 17476 19552 17540 19556
rect 22664 19612 22728 19616
rect 22664 19556 22668 19612
rect 22668 19556 22724 19612
rect 22724 19556 22728 19612
rect 22664 19552 22728 19556
rect 22744 19612 22808 19616
rect 22744 19556 22748 19612
rect 22748 19556 22804 19612
rect 22804 19556 22808 19612
rect 22744 19552 22808 19556
rect 22824 19612 22888 19616
rect 22824 19556 22828 19612
rect 22828 19556 22884 19612
rect 22884 19556 22888 19612
rect 22824 19552 22888 19556
rect 22904 19612 22968 19616
rect 22904 19556 22908 19612
rect 22908 19556 22964 19612
rect 22964 19556 22968 19612
rect 22904 19552 22968 19556
rect 3666 19068 3730 19072
rect 3666 19012 3670 19068
rect 3670 19012 3726 19068
rect 3726 19012 3730 19068
rect 3666 19008 3730 19012
rect 3746 19068 3810 19072
rect 3746 19012 3750 19068
rect 3750 19012 3806 19068
rect 3806 19012 3810 19068
rect 3746 19008 3810 19012
rect 3826 19068 3890 19072
rect 3826 19012 3830 19068
rect 3830 19012 3886 19068
rect 3886 19012 3890 19068
rect 3826 19008 3890 19012
rect 3906 19068 3970 19072
rect 3906 19012 3910 19068
rect 3910 19012 3966 19068
rect 3966 19012 3970 19068
rect 3906 19008 3970 19012
rect 9094 19068 9158 19072
rect 9094 19012 9098 19068
rect 9098 19012 9154 19068
rect 9154 19012 9158 19068
rect 9094 19008 9158 19012
rect 9174 19068 9238 19072
rect 9174 19012 9178 19068
rect 9178 19012 9234 19068
rect 9234 19012 9238 19068
rect 9174 19008 9238 19012
rect 9254 19068 9318 19072
rect 9254 19012 9258 19068
rect 9258 19012 9314 19068
rect 9314 19012 9318 19068
rect 9254 19008 9318 19012
rect 9334 19068 9398 19072
rect 9334 19012 9338 19068
rect 9338 19012 9394 19068
rect 9394 19012 9398 19068
rect 9334 19008 9398 19012
rect 14522 19068 14586 19072
rect 14522 19012 14526 19068
rect 14526 19012 14582 19068
rect 14582 19012 14586 19068
rect 14522 19008 14586 19012
rect 14602 19068 14666 19072
rect 14602 19012 14606 19068
rect 14606 19012 14662 19068
rect 14662 19012 14666 19068
rect 14602 19008 14666 19012
rect 14682 19068 14746 19072
rect 14682 19012 14686 19068
rect 14686 19012 14742 19068
rect 14742 19012 14746 19068
rect 14682 19008 14746 19012
rect 14762 19068 14826 19072
rect 14762 19012 14766 19068
rect 14766 19012 14822 19068
rect 14822 19012 14826 19068
rect 14762 19008 14826 19012
rect 19950 19068 20014 19072
rect 19950 19012 19954 19068
rect 19954 19012 20010 19068
rect 20010 19012 20014 19068
rect 19950 19008 20014 19012
rect 20030 19068 20094 19072
rect 20030 19012 20034 19068
rect 20034 19012 20090 19068
rect 20090 19012 20094 19068
rect 20030 19008 20094 19012
rect 20110 19068 20174 19072
rect 20110 19012 20114 19068
rect 20114 19012 20170 19068
rect 20170 19012 20174 19068
rect 20110 19008 20174 19012
rect 20190 19068 20254 19072
rect 20190 19012 20194 19068
rect 20194 19012 20250 19068
rect 20250 19012 20254 19068
rect 20190 19008 20254 19012
rect 6380 18524 6444 18528
rect 6380 18468 6384 18524
rect 6384 18468 6440 18524
rect 6440 18468 6444 18524
rect 6380 18464 6444 18468
rect 6460 18524 6524 18528
rect 6460 18468 6464 18524
rect 6464 18468 6520 18524
rect 6520 18468 6524 18524
rect 6460 18464 6524 18468
rect 6540 18524 6604 18528
rect 6540 18468 6544 18524
rect 6544 18468 6600 18524
rect 6600 18468 6604 18524
rect 6540 18464 6604 18468
rect 6620 18524 6684 18528
rect 6620 18468 6624 18524
rect 6624 18468 6680 18524
rect 6680 18468 6684 18524
rect 6620 18464 6684 18468
rect 11808 18524 11872 18528
rect 11808 18468 11812 18524
rect 11812 18468 11868 18524
rect 11868 18468 11872 18524
rect 11808 18464 11872 18468
rect 11888 18524 11952 18528
rect 11888 18468 11892 18524
rect 11892 18468 11948 18524
rect 11948 18468 11952 18524
rect 11888 18464 11952 18468
rect 11968 18524 12032 18528
rect 11968 18468 11972 18524
rect 11972 18468 12028 18524
rect 12028 18468 12032 18524
rect 11968 18464 12032 18468
rect 12048 18524 12112 18528
rect 12048 18468 12052 18524
rect 12052 18468 12108 18524
rect 12108 18468 12112 18524
rect 12048 18464 12112 18468
rect 17236 18524 17300 18528
rect 17236 18468 17240 18524
rect 17240 18468 17296 18524
rect 17296 18468 17300 18524
rect 17236 18464 17300 18468
rect 17316 18524 17380 18528
rect 17316 18468 17320 18524
rect 17320 18468 17376 18524
rect 17376 18468 17380 18524
rect 17316 18464 17380 18468
rect 17396 18524 17460 18528
rect 17396 18468 17400 18524
rect 17400 18468 17456 18524
rect 17456 18468 17460 18524
rect 17396 18464 17460 18468
rect 17476 18524 17540 18528
rect 17476 18468 17480 18524
rect 17480 18468 17536 18524
rect 17536 18468 17540 18524
rect 17476 18464 17540 18468
rect 22664 18524 22728 18528
rect 22664 18468 22668 18524
rect 22668 18468 22724 18524
rect 22724 18468 22728 18524
rect 22664 18464 22728 18468
rect 22744 18524 22808 18528
rect 22744 18468 22748 18524
rect 22748 18468 22804 18524
rect 22804 18468 22808 18524
rect 22744 18464 22808 18468
rect 22824 18524 22888 18528
rect 22824 18468 22828 18524
rect 22828 18468 22884 18524
rect 22884 18468 22888 18524
rect 22824 18464 22888 18468
rect 22904 18524 22968 18528
rect 22904 18468 22908 18524
rect 22908 18468 22964 18524
rect 22964 18468 22968 18524
rect 22904 18464 22968 18468
rect 3666 17980 3730 17984
rect 3666 17924 3670 17980
rect 3670 17924 3726 17980
rect 3726 17924 3730 17980
rect 3666 17920 3730 17924
rect 3746 17980 3810 17984
rect 3746 17924 3750 17980
rect 3750 17924 3806 17980
rect 3806 17924 3810 17980
rect 3746 17920 3810 17924
rect 3826 17980 3890 17984
rect 3826 17924 3830 17980
rect 3830 17924 3886 17980
rect 3886 17924 3890 17980
rect 3826 17920 3890 17924
rect 3906 17980 3970 17984
rect 3906 17924 3910 17980
rect 3910 17924 3966 17980
rect 3966 17924 3970 17980
rect 3906 17920 3970 17924
rect 9094 17980 9158 17984
rect 9094 17924 9098 17980
rect 9098 17924 9154 17980
rect 9154 17924 9158 17980
rect 9094 17920 9158 17924
rect 9174 17980 9238 17984
rect 9174 17924 9178 17980
rect 9178 17924 9234 17980
rect 9234 17924 9238 17980
rect 9174 17920 9238 17924
rect 9254 17980 9318 17984
rect 9254 17924 9258 17980
rect 9258 17924 9314 17980
rect 9314 17924 9318 17980
rect 9254 17920 9318 17924
rect 9334 17980 9398 17984
rect 9334 17924 9338 17980
rect 9338 17924 9394 17980
rect 9394 17924 9398 17980
rect 9334 17920 9398 17924
rect 14522 17980 14586 17984
rect 14522 17924 14526 17980
rect 14526 17924 14582 17980
rect 14582 17924 14586 17980
rect 14522 17920 14586 17924
rect 14602 17980 14666 17984
rect 14602 17924 14606 17980
rect 14606 17924 14662 17980
rect 14662 17924 14666 17980
rect 14602 17920 14666 17924
rect 14682 17980 14746 17984
rect 14682 17924 14686 17980
rect 14686 17924 14742 17980
rect 14742 17924 14746 17980
rect 14682 17920 14746 17924
rect 14762 17980 14826 17984
rect 14762 17924 14766 17980
rect 14766 17924 14822 17980
rect 14822 17924 14826 17980
rect 14762 17920 14826 17924
rect 19950 17980 20014 17984
rect 19950 17924 19954 17980
rect 19954 17924 20010 17980
rect 20010 17924 20014 17980
rect 19950 17920 20014 17924
rect 20030 17980 20094 17984
rect 20030 17924 20034 17980
rect 20034 17924 20090 17980
rect 20090 17924 20094 17980
rect 20030 17920 20094 17924
rect 20110 17980 20174 17984
rect 20110 17924 20114 17980
rect 20114 17924 20170 17980
rect 20170 17924 20174 17980
rect 20110 17920 20174 17924
rect 20190 17980 20254 17984
rect 20190 17924 20194 17980
rect 20194 17924 20250 17980
rect 20250 17924 20254 17980
rect 20190 17920 20254 17924
rect 6380 17436 6444 17440
rect 6380 17380 6384 17436
rect 6384 17380 6440 17436
rect 6440 17380 6444 17436
rect 6380 17376 6444 17380
rect 6460 17436 6524 17440
rect 6460 17380 6464 17436
rect 6464 17380 6520 17436
rect 6520 17380 6524 17436
rect 6460 17376 6524 17380
rect 6540 17436 6604 17440
rect 6540 17380 6544 17436
rect 6544 17380 6600 17436
rect 6600 17380 6604 17436
rect 6540 17376 6604 17380
rect 6620 17436 6684 17440
rect 6620 17380 6624 17436
rect 6624 17380 6680 17436
rect 6680 17380 6684 17436
rect 6620 17376 6684 17380
rect 11808 17436 11872 17440
rect 11808 17380 11812 17436
rect 11812 17380 11868 17436
rect 11868 17380 11872 17436
rect 11808 17376 11872 17380
rect 11888 17436 11952 17440
rect 11888 17380 11892 17436
rect 11892 17380 11948 17436
rect 11948 17380 11952 17436
rect 11888 17376 11952 17380
rect 11968 17436 12032 17440
rect 11968 17380 11972 17436
rect 11972 17380 12028 17436
rect 12028 17380 12032 17436
rect 11968 17376 12032 17380
rect 12048 17436 12112 17440
rect 12048 17380 12052 17436
rect 12052 17380 12108 17436
rect 12108 17380 12112 17436
rect 12048 17376 12112 17380
rect 17236 17436 17300 17440
rect 17236 17380 17240 17436
rect 17240 17380 17296 17436
rect 17296 17380 17300 17436
rect 17236 17376 17300 17380
rect 17316 17436 17380 17440
rect 17316 17380 17320 17436
rect 17320 17380 17376 17436
rect 17376 17380 17380 17436
rect 17316 17376 17380 17380
rect 17396 17436 17460 17440
rect 17396 17380 17400 17436
rect 17400 17380 17456 17436
rect 17456 17380 17460 17436
rect 17396 17376 17460 17380
rect 17476 17436 17540 17440
rect 17476 17380 17480 17436
rect 17480 17380 17536 17436
rect 17536 17380 17540 17436
rect 17476 17376 17540 17380
rect 22664 17436 22728 17440
rect 22664 17380 22668 17436
rect 22668 17380 22724 17436
rect 22724 17380 22728 17436
rect 22664 17376 22728 17380
rect 22744 17436 22808 17440
rect 22744 17380 22748 17436
rect 22748 17380 22804 17436
rect 22804 17380 22808 17436
rect 22744 17376 22808 17380
rect 22824 17436 22888 17440
rect 22824 17380 22828 17436
rect 22828 17380 22884 17436
rect 22884 17380 22888 17436
rect 22824 17376 22888 17380
rect 22904 17436 22968 17440
rect 22904 17380 22908 17436
rect 22908 17380 22964 17436
rect 22964 17380 22968 17436
rect 22904 17376 22968 17380
rect 3666 16892 3730 16896
rect 3666 16836 3670 16892
rect 3670 16836 3726 16892
rect 3726 16836 3730 16892
rect 3666 16832 3730 16836
rect 3746 16892 3810 16896
rect 3746 16836 3750 16892
rect 3750 16836 3806 16892
rect 3806 16836 3810 16892
rect 3746 16832 3810 16836
rect 3826 16892 3890 16896
rect 3826 16836 3830 16892
rect 3830 16836 3886 16892
rect 3886 16836 3890 16892
rect 3826 16832 3890 16836
rect 3906 16892 3970 16896
rect 3906 16836 3910 16892
rect 3910 16836 3966 16892
rect 3966 16836 3970 16892
rect 3906 16832 3970 16836
rect 9094 16892 9158 16896
rect 9094 16836 9098 16892
rect 9098 16836 9154 16892
rect 9154 16836 9158 16892
rect 9094 16832 9158 16836
rect 9174 16892 9238 16896
rect 9174 16836 9178 16892
rect 9178 16836 9234 16892
rect 9234 16836 9238 16892
rect 9174 16832 9238 16836
rect 9254 16892 9318 16896
rect 9254 16836 9258 16892
rect 9258 16836 9314 16892
rect 9314 16836 9318 16892
rect 9254 16832 9318 16836
rect 9334 16892 9398 16896
rect 9334 16836 9338 16892
rect 9338 16836 9394 16892
rect 9394 16836 9398 16892
rect 9334 16832 9398 16836
rect 14522 16892 14586 16896
rect 14522 16836 14526 16892
rect 14526 16836 14582 16892
rect 14582 16836 14586 16892
rect 14522 16832 14586 16836
rect 14602 16892 14666 16896
rect 14602 16836 14606 16892
rect 14606 16836 14662 16892
rect 14662 16836 14666 16892
rect 14602 16832 14666 16836
rect 14682 16892 14746 16896
rect 14682 16836 14686 16892
rect 14686 16836 14742 16892
rect 14742 16836 14746 16892
rect 14682 16832 14746 16836
rect 14762 16892 14826 16896
rect 14762 16836 14766 16892
rect 14766 16836 14822 16892
rect 14822 16836 14826 16892
rect 14762 16832 14826 16836
rect 19950 16892 20014 16896
rect 19950 16836 19954 16892
rect 19954 16836 20010 16892
rect 20010 16836 20014 16892
rect 19950 16832 20014 16836
rect 20030 16892 20094 16896
rect 20030 16836 20034 16892
rect 20034 16836 20090 16892
rect 20090 16836 20094 16892
rect 20030 16832 20094 16836
rect 20110 16892 20174 16896
rect 20110 16836 20114 16892
rect 20114 16836 20170 16892
rect 20170 16836 20174 16892
rect 20110 16832 20174 16836
rect 20190 16892 20254 16896
rect 20190 16836 20194 16892
rect 20194 16836 20250 16892
rect 20250 16836 20254 16892
rect 20190 16832 20254 16836
rect 6380 16348 6444 16352
rect 6380 16292 6384 16348
rect 6384 16292 6440 16348
rect 6440 16292 6444 16348
rect 6380 16288 6444 16292
rect 6460 16348 6524 16352
rect 6460 16292 6464 16348
rect 6464 16292 6520 16348
rect 6520 16292 6524 16348
rect 6460 16288 6524 16292
rect 6540 16348 6604 16352
rect 6540 16292 6544 16348
rect 6544 16292 6600 16348
rect 6600 16292 6604 16348
rect 6540 16288 6604 16292
rect 6620 16348 6684 16352
rect 6620 16292 6624 16348
rect 6624 16292 6680 16348
rect 6680 16292 6684 16348
rect 6620 16288 6684 16292
rect 11808 16348 11872 16352
rect 11808 16292 11812 16348
rect 11812 16292 11868 16348
rect 11868 16292 11872 16348
rect 11808 16288 11872 16292
rect 11888 16348 11952 16352
rect 11888 16292 11892 16348
rect 11892 16292 11948 16348
rect 11948 16292 11952 16348
rect 11888 16288 11952 16292
rect 11968 16348 12032 16352
rect 11968 16292 11972 16348
rect 11972 16292 12028 16348
rect 12028 16292 12032 16348
rect 11968 16288 12032 16292
rect 12048 16348 12112 16352
rect 12048 16292 12052 16348
rect 12052 16292 12108 16348
rect 12108 16292 12112 16348
rect 12048 16288 12112 16292
rect 17236 16348 17300 16352
rect 17236 16292 17240 16348
rect 17240 16292 17296 16348
rect 17296 16292 17300 16348
rect 17236 16288 17300 16292
rect 17316 16348 17380 16352
rect 17316 16292 17320 16348
rect 17320 16292 17376 16348
rect 17376 16292 17380 16348
rect 17316 16288 17380 16292
rect 17396 16348 17460 16352
rect 17396 16292 17400 16348
rect 17400 16292 17456 16348
rect 17456 16292 17460 16348
rect 17396 16288 17460 16292
rect 17476 16348 17540 16352
rect 17476 16292 17480 16348
rect 17480 16292 17536 16348
rect 17536 16292 17540 16348
rect 17476 16288 17540 16292
rect 22664 16348 22728 16352
rect 22664 16292 22668 16348
rect 22668 16292 22724 16348
rect 22724 16292 22728 16348
rect 22664 16288 22728 16292
rect 22744 16348 22808 16352
rect 22744 16292 22748 16348
rect 22748 16292 22804 16348
rect 22804 16292 22808 16348
rect 22744 16288 22808 16292
rect 22824 16348 22888 16352
rect 22824 16292 22828 16348
rect 22828 16292 22884 16348
rect 22884 16292 22888 16348
rect 22824 16288 22888 16292
rect 22904 16348 22968 16352
rect 22904 16292 22908 16348
rect 22908 16292 22964 16348
rect 22964 16292 22968 16348
rect 22904 16288 22968 16292
rect 3666 15804 3730 15808
rect 3666 15748 3670 15804
rect 3670 15748 3726 15804
rect 3726 15748 3730 15804
rect 3666 15744 3730 15748
rect 3746 15804 3810 15808
rect 3746 15748 3750 15804
rect 3750 15748 3806 15804
rect 3806 15748 3810 15804
rect 3746 15744 3810 15748
rect 3826 15804 3890 15808
rect 3826 15748 3830 15804
rect 3830 15748 3886 15804
rect 3886 15748 3890 15804
rect 3826 15744 3890 15748
rect 3906 15804 3970 15808
rect 3906 15748 3910 15804
rect 3910 15748 3966 15804
rect 3966 15748 3970 15804
rect 3906 15744 3970 15748
rect 9094 15804 9158 15808
rect 9094 15748 9098 15804
rect 9098 15748 9154 15804
rect 9154 15748 9158 15804
rect 9094 15744 9158 15748
rect 9174 15804 9238 15808
rect 9174 15748 9178 15804
rect 9178 15748 9234 15804
rect 9234 15748 9238 15804
rect 9174 15744 9238 15748
rect 9254 15804 9318 15808
rect 9254 15748 9258 15804
rect 9258 15748 9314 15804
rect 9314 15748 9318 15804
rect 9254 15744 9318 15748
rect 9334 15804 9398 15808
rect 9334 15748 9338 15804
rect 9338 15748 9394 15804
rect 9394 15748 9398 15804
rect 9334 15744 9398 15748
rect 14522 15804 14586 15808
rect 14522 15748 14526 15804
rect 14526 15748 14582 15804
rect 14582 15748 14586 15804
rect 14522 15744 14586 15748
rect 14602 15804 14666 15808
rect 14602 15748 14606 15804
rect 14606 15748 14662 15804
rect 14662 15748 14666 15804
rect 14602 15744 14666 15748
rect 14682 15804 14746 15808
rect 14682 15748 14686 15804
rect 14686 15748 14742 15804
rect 14742 15748 14746 15804
rect 14682 15744 14746 15748
rect 14762 15804 14826 15808
rect 14762 15748 14766 15804
rect 14766 15748 14822 15804
rect 14822 15748 14826 15804
rect 14762 15744 14826 15748
rect 19950 15804 20014 15808
rect 19950 15748 19954 15804
rect 19954 15748 20010 15804
rect 20010 15748 20014 15804
rect 19950 15744 20014 15748
rect 20030 15804 20094 15808
rect 20030 15748 20034 15804
rect 20034 15748 20090 15804
rect 20090 15748 20094 15804
rect 20030 15744 20094 15748
rect 20110 15804 20174 15808
rect 20110 15748 20114 15804
rect 20114 15748 20170 15804
rect 20170 15748 20174 15804
rect 20110 15744 20174 15748
rect 20190 15804 20254 15808
rect 20190 15748 20194 15804
rect 20194 15748 20250 15804
rect 20250 15748 20254 15804
rect 20190 15744 20254 15748
rect 6380 15260 6444 15264
rect 6380 15204 6384 15260
rect 6384 15204 6440 15260
rect 6440 15204 6444 15260
rect 6380 15200 6444 15204
rect 6460 15260 6524 15264
rect 6460 15204 6464 15260
rect 6464 15204 6520 15260
rect 6520 15204 6524 15260
rect 6460 15200 6524 15204
rect 6540 15260 6604 15264
rect 6540 15204 6544 15260
rect 6544 15204 6600 15260
rect 6600 15204 6604 15260
rect 6540 15200 6604 15204
rect 6620 15260 6684 15264
rect 6620 15204 6624 15260
rect 6624 15204 6680 15260
rect 6680 15204 6684 15260
rect 6620 15200 6684 15204
rect 11808 15260 11872 15264
rect 11808 15204 11812 15260
rect 11812 15204 11868 15260
rect 11868 15204 11872 15260
rect 11808 15200 11872 15204
rect 11888 15260 11952 15264
rect 11888 15204 11892 15260
rect 11892 15204 11948 15260
rect 11948 15204 11952 15260
rect 11888 15200 11952 15204
rect 11968 15260 12032 15264
rect 11968 15204 11972 15260
rect 11972 15204 12028 15260
rect 12028 15204 12032 15260
rect 11968 15200 12032 15204
rect 12048 15260 12112 15264
rect 12048 15204 12052 15260
rect 12052 15204 12108 15260
rect 12108 15204 12112 15260
rect 12048 15200 12112 15204
rect 17236 15260 17300 15264
rect 17236 15204 17240 15260
rect 17240 15204 17296 15260
rect 17296 15204 17300 15260
rect 17236 15200 17300 15204
rect 17316 15260 17380 15264
rect 17316 15204 17320 15260
rect 17320 15204 17376 15260
rect 17376 15204 17380 15260
rect 17316 15200 17380 15204
rect 17396 15260 17460 15264
rect 17396 15204 17400 15260
rect 17400 15204 17456 15260
rect 17456 15204 17460 15260
rect 17396 15200 17460 15204
rect 17476 15260 17540 15264
rect 17476 15204 17480 15260
rect 17480 15204 17536 15260
rect 17536 15204 17540 15260
rect 17476 15200 17540 15204
rect 22664 15260 22728 15264
rect 22664 15204 22668 15260
rect 22668 15204 22724 15260
rect 22724 15204 22728 15260
rect 22664 15200 22728 15204
rect 22744 15260 22808 15264
rect 22744 15204 22748 15260
rect 22748 15204 22804 15260
rect 22804 15204 22808 15260
rect 22744 15200 22808 15204
rect 22824 15260 22888 15264
rect 22824 15204 22828 15260
rect 22828 15204 22884 15260
rect 22884 15204 22888 15260
rect 22824 15200 22888 15204
rect 22904 15260 22968 15264
rect 22904 15204 22908 15260
rect 22908 15204 22964 15260
rect 22964 15204 22968 15260
rect 22904 15200 22968 15204
rect 3666 14716 3730 14720
rect 3666 14660 3670 14716
rect 3670 14660 3726 14716
rect 3726 14660 3730 14716
rect 3666 14656 3730 14660
rect 3746 14716 3810 14720
rect 3746 14660 3750 14716
rect 3750 14660 3806 14716
rect 3806 14660 3810 14716
rect 3746 14656 3810 14660
rect 3826 14716 3890 14720
rect 3826 14660 3830 14716
rect 3830 14660 3886 14716
rect 3886 14660 3890 14716
rect 3826 14656 3890 14660
rect 3906 14716 3970 14720
rect 3906 14660 3910 14716
rect 3910 14660 3966 14716
rect 3966 14660 3970 14716
rect 3906 14656 3970 14660
rect 9094 14716 9158 14720
rect 9094 14660 9098 14716
rect 9098 14660 9154 14716
rect 9154 14660 9158 14716
rect 9094 14656 9158 14660
rect 9174 14716 9238 14720
rect 9174 14660 9178 14716
rect 9178 14660 9234 14716
rect 9234 14660 9238 14716
rect 9174 14656 9238 14660
rect 9254 14716 9318 14720
rect 9254 14660 9258 14716
rect 9258 14660 9314 14716
rect 9314 14660 9318 14716
rect 9254 14656 9318 14660
rect 9334 14716 9398 14720
rect 9334 14660 9338 14716
rect 9338 14660 9394 14716
rect 9394 14660 9398 14716
rect 9334 14656 9398 14660
rect 14522 14716 14586 14720
rect 14522 14660 14526 14716
rect 14526 14660 14582 14716
rect 14582 14660 14586 14716
rect 14522 14656 14586 14660
rect 14602 14716 14666 14720
rect 14602 14660 14606 14716
rect 14606 14660 14662 14716
rect 14662 14660 14666 14716
rect 14602 14656 14666 14660
rect 14682 14716 14746 14720
rect 14682 14660 14686 14716
rect 14686 14660 14742 14716
rect 14742 14660 14746 14716
rect 14682 14656 14746 14660
rect 14762 14716 14826 14720
rect 14762 14660 14766 14716
rect 14766 14660 14822 14716
rect 14822 14660 14826 14716
rect 14762 14656 14826 14660
rect 19950 14716 20014 14720
rect 19950 14660 19954 14716
rect 19954 14660 20010 14716
rect 20010 14660 20014 14716
rect 19950 14656 20014 14660
rect 20030 14716 20094 14720
rect 20030 14660 20034 14716
rect 20034 14660 20090 14716
rect 20090 14660 20094 14716
rect 20030 14656 20094 14660
rect 20110 14716 20174 14720
rect 20110 14660 20114 14716
rect 20114 14660 20170 14716
rect 20170 14660 20174 14716
rect 20110 14656 20174 14660
rect 20190 14716 20254 14720
rect 20190 14660 20194 14716
rect 20194 14660 20250 14716
rect 20250 14660 20254 14716
rect 20190 14656 20254 14660
rect 6380 14172 6444 14176
rect 6380 14116 6384 14172
rect 6384 14116 6440 14172
rect 6440 14116 6444 14172
rect 6380 14112 6444 14116
rect 6460 14172 6524 14176
rect 6460 14116 6464 14172
rect 6464 14116 6520 14172
rect 6520 14116 6524 14172
rect 6460 14112 6524 14116
rect 6540 14172 6604 14176
rect 6540 14116 6544 14172
rect 6544 14116 6600 14172
rect 6600 14116 6604 14172
rect 6540 14112 6604 14116
rect 6620 14172 6684 14176
rect 6620 14116 6624 14172
rect 6624 14116 6680 14172
rect 6680 14116 6684 14172
rect 6620 14112 6684 14116
rect 11808 14172 11872 14176
rect 11808 14116 11812 14172
rect 11812 14116 11868 14172
rect 11868 14116 11872 14172
rect 11808 14112 11872 14116
rect 11888 14172 11952 14176
rect 11888 14116 11892 14172
rect 11892 14116 11948 14172
rect 11948 14116 11952 14172
rect 11888 14112 11952 14116
rect 11968 14172 12032 14176
rect 11968 14116 11972 14172
rect 11972 14116 12028 14172
rect 12028 14116 12032 14172
rect 11968 14112 12032 14116
rect 12048 14172 12112 14176
rect 12048 14116 12052 14172
rect 12052 14116 12108 14172
rect 12108 14116 12112 14172
rect 12048 14112 12112 14116
rect 17236 14172 17300 14176
rect 17236 14116 17240 14172
rect 17240 14116 17296 14172
rect 17296 14116 17300 14172
rect 17236 14112 17300 14116
rect 17316 14172 17380 14176
rect 17316 14116 17320 14172
rect 17320 14116 17376 14172
rect 17376 14116 17380 14172
rect 17316 14112 17380 14116
rect 17396 14172 17460 14176
rect 17396 14116 17400 14172
rect 17400 14116 17456 14172
rect 17456 14116 17460 14172
rect 17396 14112 17460 14116
rect 17476 14172 17540 14176
rect 17476 14116 17480 14172
rect 17480 14116 17536 14172
rect 17536 14116 17540 14172
rect 17476 14112 17540 14116
rect 22664 14172 22728 14176
rect 22664 14116 22668 14172
rect 22668 14116 22724 14172
rect 22724 14116 22728 14172
rect 22664 14112 22728 14116
rect 22744 14172 22808 14176
rect 22744 14116 22748 14172
rect 22748 14116 22804 14172
rect 22804 14116 22808 14172
rect 22744 14112 22808 14116
rect 22824 14172 22888 14176
rect 22824 14116 22828 14172
rect 22828 14116 22884 14172
rect 22884 14116 22888 14172
rect 22824 14112 22888 14116
rect 22904 14172 22968 14176
rect 22904 14116 22908 14172
rect 22908 14116 22964 14172
rect 22964 14116 22968 14172
rect 22904 14112 22968 14116
rect 3666 13628 3730 13632
rect 3666 13572 3670 13628
rect 3670 13572 3726 13628
rect 3726 13572 3730 13628
rect 3666 13568 3730 13572
rect 3746 13628 3810 13632
rect 3746 13572 3750 13628
rect 3750 13572 3806 13628
rect 3806 13572 3810 13628
rect 3746 13568 3810 13572
rect 3826 13628 3890 13632
rect 3826 13572 3830 13628
rect 3830 13572 3886 13628
rect 3886 13572 3890 13628
rect 3826 13568 3890 13572
rect 3906 13628 3970 13632
rect 3906 13572 3910 13628
rect 3910 13572 3966 13628
rect 3966 13572 3970 13628
rect 3906 13568 3970 13572
rect 9094 13628 9158 13632
rect 9094 13572 9098 13628
rect 9098 13572 9154 13628
rect 9154 13572 9158 13628
rect 9094 13568 9158 13572
rect 9174 13628 9238 13632
rect 9174 13572 9178 13628
rect 9178 13572 9234 13628
rect 9234 13572 9238 13628
rect 9174 13568 9238 13572
rect 9254 13628 9318 13632
rect 9254 13572 9258 13628
rect 9258 13572 9314 13628
rect 9314 13572 9318 13628
rect 9254 13568 9318 13572
rect 9334 13628 9398 13632
rect 9334 13572 9338 13628
rect 9338 13572 9394 13628
rect 9394 13572 9398 13628
rect 9334 13568 9398 13572
rect 14522 13628 14586 13632
rect 14522 13572 14526 13628
rect 14526 13572 14582 13628
rect 14582 13572 14586 13628
rect 14522 13568 14586 13572
rect 14602 13628 14666 13632
rect 14602 13572 14606 13628
rect 14606 13572 14662 13628
rect 14662 13572 14666 13628
rect 14602 13568 14666 13572
rect 14682 13628 14746 13632
rect 14682 13572 14686 13628
rect 14686 13572 14742 13628
rect 14742 13572 14746 13628
rect 14682 13568 14746 13572
rect 14762 13628 14826 13632
rect 14762 13572 14766 13628
rect 14766 13572 14822 13628
rect 14822 13572 14826 13628
rect 14762 13568 14826 13572
rect 19950 13628 20014 13632
rect 19950 13572 19954 13628
rect 19954 13572 20010 13628
rect 20010 13572 20014 13628
rect 19950 13568 20014 13572
rect 20030 13628 20094 13632
rect 20030 13572 20034 13628
rect 20034 13572 20090 13628
rect 20090 13572 20094 13628
rect 20030 13568 20094 13572
rect 20110 13628 20174 13632
rect 20110 13572 20114 13628
rect 20114 13572 20170 13628
rect 20170 13572 20174 13628
rect 20110 13568 20174 13572
rect 20190 13628 20254 13632
rect 20190 13572 20194 13628
rect 20194 13572 20250 13628
rect 20250 13572 20254 13628
rect 20190 13568 20254 13572
rect 6380 13084 6444 13088
rect 6380 13028 6384 13084
rect 6384 13028 6440 13084
rect 6440 13028 6444 13084
rect 6380 13024 6444 13028
rect 6460 13084 6524 13088
rect 6460 13028 6464 13084
rect 6464 13028 6520 13084
rect 6520 13028 6524 13084
rect 6460 13024 6524 13028
rect 6540 13084 6604 13088
rect 6540 13028 6544 13084
rect 6544 13028 6600 13084
rect 6600 13028 6604 13084
rect 6540 13024 6604 13028
rect 6620 13084 6684 13088
rect 6620 13028 6624 13084
rect 6624 13028 6680 13084
rect 6680 13028 6684 13084
rect 6620 13024 6684 13028
rect 11808 13084 11872 13088
rect 11808 13028 11812 13084
rect 11812 13028 11868 13084
rect 11868 13028 11872 13084
rect 11808 13024 11872 13028
rect 11888 13084 11952 13088
rect 11888 13028 11892 13084
rect 11892 13028 11948 13084
rect 11948 13028 11952 13084
rect 11888 13024 11952 13028
rect 11968 13084 12032 13088
rect 11968 13028 11972 13084
rect 11972 13028 12028 13084
rect 12028 13028 12032 13084
rect 11968 13024 12032 13028
rect 12048 13084 12112 13088
rect 12048 13028 12052 13084
rect 12052 13028 12108 13084
rect 12108 13028 12112 13084
rect 12048 13024 12112 13028
rect 17236 13084 17300 13088
rect 17236 13028 17240 13084
rect 17240 13028 17296 13084
rect 17296 13028 17300 13084
rect 17236 13024 17300 13028
rect 17316 13084 17380 13088
rect 17316 13028 17320 13084
rect 17320 13028 17376 13084
rect 17376 13028 17380 13084
rect 17316 13024 17380 13028
rect 17396 13084 17460 13088
rect 17396 13028 17400 13084
rect 17400 13028 17456 13084
rect 17456 13028 17460 13084
rect 17396 13024 17460 13028
rect 17476 13084 17540 13088
rect 17476 13028 17480 13084
rect 17480 13028 17536 13084
rect 17536 13028 17540 13084
rect 17476 13024 17540 13028
rect 22664 13084 22728 13088
rect 22664 13028 22668 13084
rect 22668 13028 22724 13084
rect 22724 13028 22728 13084
rect 22664 13024 22728 13028
rect 22744 13084 22808 13088
rect 22744 13028 22748 13084
rect 22748 13028 22804 13084
rect 22804 13028 22808 13084
rect 22744 13024 22808 13028
rect 22824 13084 22888 13088
rect 22824 13028 22828 13084
rect 22828 13028 22884 13084
rect 22884 13028 22888 13084
rect 22824 13024 22888 13028
rect 22904 13084 22968 13088
rect 22904 13028 22908 13084
rect 22908 13028 22964 13084
rect 22964 13028 22968 13084
rect 22904 13024 22968 13028
rect 3666 12540 3730 12544
rect 3666 12484 3670 12540
rect 3670 12484 3726 12540
rect 3726 12484 3730 12540
rect 3666 12480 3730 12484
rect 3746 12540 3810 12544
rect 3746 12484 3750 12540
rect 3750 12484 3806 12540
rect 3806 12484 3810 12540
rect 3746 12480 3810 12484
rect 3826 12540 3890 12544
rect 3826 12484 3830 12540
rect 3830 12484 3886 12540
rect 3886 12484 3890 12540
rect 3826 12480 3890 12484
rect 3906 12540 3970 12544
rect 3906 12484 3910 12540
rect 3910 12484 3966 12540
rect 3966 12484 3970 12540
rect 3906 12480 3970 12484
rect 9094 12540 9158 12544
rect 9094 12484 9098 12540
rect 9098 12484 9154 12540
rect 9154 12484 9158 12540
rect 9094 12480 9158 12484
rect 9174 12540 9238 12544
rect 9174 12484 9178 12540
rect 9178 12484 9234 12540
rect 9234 12484 9238 12540
rect 9174 12480 9238 12484
rect 9254 12540 9318 12544
rect 9254 12484 9258 12540
rect 9258 12484 9314 12540
rect 9314 12484 9318 12540
rect 9254 12480 9318 12484
rect 9334 12540 9398 12544
rect 9334 12484 9338 12540
rect 9338 12484 9394 12540
rect 9394 12484 9398 12540
rect 9334 12480 9398 12484
rect 14522 12540 14586 12544
rect 14522 12484 14526 12540
rect 14526 12484 14582 12540
rect 14582 12484 14586 12540
rect 14522 12480 14586 12484
rect 14602 12540 14666 12544
rect 14602 12484 14606 12540
rect 14606 12484 14662 12540
rect 14662 12484 14666 12540
rect 14602 12480 14666 12484
rect 14682 12540 14746 12544
rect 14682 12484 14686 12540
rect 14686 12484 14742 12540
rect 14742 12484 14746 12540
rect 14682 12480 14746 12484
rect 14762 12540 14826 12544
rect 14762 12484 14766 12540
rect 14766 12484 14822 12540
rect 14822 12484 14826 12540
rect 14762 12480 14826 12484
rect 19950 12540 20014 12544
rect 19950 12484 19954 12540
rect 19954 12484 20010 12540
rect 20010 12484 20014 12540
rect 19950 12480 20014 12484
rect 20030 12540 20094 12544
rect 20030 12484 20034 12540
rect 20034 12484 20090 12540
rect 20090 12484 20094 12540
rect 20030 12480 20094 12484
rect 20110 12540 20174 12544
rect 20110 12484 20114 12540
rect 20114 12484 20170 12540
rect 20170 12484 20174 12540
rect 20110 12480 20174 12484
rect 20190 12540 20254 12544
rect 20190 12484 20194 12540
rect 20194 12484 20250 12540
rect 20250 12484 20254 12540
rect 20190 12480 20254 12484
rect 6380 11996 6444 12000
rect 6380 11940 6384 11996
rect 6384 11940 6440 11996
rect 6440 11940 6444 11996
rect 6380 11936 6444 11940
rect 6460 11996 6524 12000
rect 6460 11940 6464 11996
rect 6464 11940 6520 11996
rect 6520 11940 6524 11996
rect 6460 11936 6524 11940
rect 6540 11996 6604 12000
rect 6540 11940 6544 11996
rect 6544 11940 6600 11996
rect 6600 11940 6604 11996
rect 6540 11936 6604 11940
rect 6620 11996 6684 12000
rect 6620 11940 6624 11996
rect 6624 11940 6680 11996
rect 6680 11940 6684 11996
rect 6620 11936 6684 11940
rect 11808 11996 11872 12000
rect 11808 11940 11812 11996
rect 11812 11940 11868 11996
rect 11868 11940 11872 11996
rect 11808 11936 11872 11940
rect 11888 11996 11952 12000
rect 11888 11940 11892 11996
rect 11892 11940 11948 11996
rect 11948 11940 11952 11996
rect 11888 11936 11952 11940
rect 11968 11996 12032 12000
rect 11968 11940 11972 11996
rect 11972 11940 12028 11996
rect 12028 11940 12032 11996
rect 11968 11936 12032 11940
rect 12048 11996 12112 12000
rect 12048 11940 12052 11996
rect 12052 11940 12108 11996
rect 12108 11940 12112 11996
rect 12048 11936 12112 11940
rect 17236 11996 17300 12000
rect 17236 11940 17240 11996
rect 17240 11940 17296 11996
rect 17296 11940 17300 11996
rect 17236 11936 17300 11940
rect 17316 11996 17380 12000
rect 17316 11940 17320 11996
rect 17320 11940 17376 11996
rect 17376 11940 17380 11996
rect 17316 11936 17380 11940
rect 17396 11996 17460 12000
rect 17396 11940 17400 11996
rect 17400 11940 17456 11996
rect 17456 11940 17460 11996
rect 17396 11936 17460 11940
rect 17476 11996 17540 12000
rect 17476 11940 17480 11996
rect 17480 11940 17536 11996
rect 17536 11940 17540 11996
rect 17476 11936 17540 11940
rect 22664 11996 22728 12000
rect 22664 11940 22668 11996
rect 22668 11940 22724 11996
rect 22724 11940 22728 11996
rect 22664 11936 22728 11940
rect 22744 11996 22808 12000
rect 22744 11940 22748 11996
rect 22748 11940 22804 11996
rect 22804 11940 22808 11996
rect 22744 11936 22808 11940
rect 22824 11996 22888 12000
rect 22824 11940 22828 11996
rect 22828 11940 22884 11996
rect 22884 11940 22888 11996
rect 22824 11936 22888 11940
rect 22904 11996 22968 12000
rect 22904 11940 22908 11996
rect 22908 11940 22964 11996
rect 22964 11940 22968 11996
rect 22904 11936 22968 11940
rect 3666 11452 3730 11456
rect 3666 11396 3670 11452
rect 3670 11396 3726 11452
rect 3726 11396 3730 11452
rect 3666 11392 3730 11396
rect 3746 11452 3810 11456
rect 3746 11396 3750 11452
rect 3750 11396 3806 11452
rect 3806 11396 3810 11452
rect 3746 11392 3810 11396
rect 3826 11452 3890 11456
rect 3826 11396 3830 11452
rect 3830 11396 3886 11452
rect 3886 11396 3890 11452
rect 3826 11392 3890 11396
rect 3906 11452 3970 11456
rect 3906 11396 3910 11452
rect 3910 11396 3966 11452
rect 3966 11396 3970 11452
rect 3906 11392 3970 11396
rect 9094 11452 9158 11456
rect 9094 11396 9098 11452
rect 9098 11396 9154 11452
rect 9154 11396 9158 11452
rect 9094 11392 9158 11396
rect 9174 11452 9238 11456
rect 9174 11396 9178 11452
rect 9178 11396 9234 11452
rect 9234 11396 9238 11452
rect 9174 11392 9238 11396
rect 9254 11452 9318 11456
rect 9254 11396 9258 11452
rect 9258 11396 9314 11452
rect 9314 11396 9318 11452
rect 9254 11392 9318 11396
rect 9334 11452 9398 11456
rect 9334 11396 9338 11452
rect 9338 11396 9394 11452
rect 9394 11396 9398 11452
rect 9334 11392 9398 11396
rect 14522 11452 14586 11456
rect 14522 11396 14526 11452
rect 14526 11396 14582 11452
rect 14582 11396 14586 11452
rect 14522 11392 14586 11396
rect 14602 11452 14666 11456
rect 14602 11396 14606 11452
rect 14606 11396 14662 11452
rect 14662 11396 14666 11452
rect 14602 11392 14666 11396
rect 14682 11452 14746 11456
rect 14682 11396 14686 11452
rect 14686 11396 14742 11452
rect 14742 11396 14746 11452
rect 14682 11392 14746 11396
rect 14762 11452 14826 11456
rect 14762 11396 14766 11452
rect 14766 11396 14822 11452
rect 14822 11396 14826 11452
rect 14762 11392 14826 11396
rect 19950 11452 20014 11456
rect 19950 11396 19954 11452
rect 19954 11396 20010 11452
rect 20010 11396 20014 11452
rect 19950 11392 20014 11396
rect 20030 11452 20094 11456
rect 20030 11396 20034 11452
rect 20034 11396 20090 11452
rect 20090 11396 20094 11452
rect 20030 11392 20094 11396
rect 20110 11452 20174 11456
rect 20110 11396 20114 11452
rect 20114 11396 20170 11452
rect 20170 11396 20174 11452
rect 20110 11392 20174 11396
rect 20190 11452 20254 11456
rect 20190 11396 20194 11452
rect 20194 11396 20250 11452
rect 20250 11396 20254 11452
rect 20190 11392 20254 11396
rect 6380 10908 6444 10912
rect 6380 10852 6384 10908
rect 6384 10852 6440 10908
rect 6440 10852 6444 10908
rect 6380 10848 6444 10852
rect 6460 10908 6524 10912
rect 6460 10852 6464 10908
rect 6464 10852 6520 10908
rect 6520 10852 6524 10908
rect 6460 10848 6524 10852
rect 6540 10908 6604 10912
rect 6540 10852 6544 10908
rect 6544 10852 6600 10908
rect 6600 10852 6604 10908
rect 6540 10848 6604 10852
rect 6620 10908 6684 10912
rect 6620 10852 6624 10908
rect 6624 10852 6680 10908
rect 6680 10852 6684 10908
rect 6620 10848 6684 10852
rect 11808 10908 11872 10912
rect 11808 10852 11812 10908
rect 11812 10852 11868 10908
rect 11868 10852 11872 10908
rect 11808 10848 11872 10852
rect 11888 10908 11952 10912
rect 11888 10852 11892 10908
rect 11892 10852 11948 10908
rect 11948 10852 11952 10908
rect 11888 10848 11952 10852
rect 11968 10908 12032 10912
rect 11968 10852 11972 10908
rect 11972 10852 12028 10908
rect 12028 10852 12032 10908
rect 11968 10848 12032 10852
rect 12048 10908 12112 10912
rect 12048 10852 12052 10908
rect 12052 10852 12108 10908
rect 12108 10852 12112 10908
rect 12048 10848 12112 10852
rect 17236 10908 17300 10912
rect 17236 10852 17240 10908
rect 17240 10852 17296 10908
rect 17296 10852 17300 10908
rect 17236 10848 17300 10852
rect 17316 10908 17380 10912
rect 17316 10852 17320 10908
rect 17320 10852 17376 10908
rect 17376 10852 17380 10908
rect 17316 10848 17380 10852
rect 17396 10908 17460 10912
rect 17396 10852 17400 10908
rect 17400 10852 17456 10908
rect 17456 10852 17460 10908
rect 17396 10848 17460 10852
rect 17476 10908 17540 10912
rect 17476 10852 17480 10908
rect 17480 10852 17536 10908
rect 17536 10852 17540 10908
rect 17476 10848 17540 10852
rect 22664 10908 22728 10912
rect 22664 10852 22668 10908
rect 22668 10852 22724 10908
rect 22724 10852 22728 10908
rect 22664 10848 22728 10852
rect 22744 10908 22808 10912
rect 22744 10852 22748 10908
rect 22748 10852 22804 10908
rect 22804 10852 22808 10908
rect 22744 10848 22808 10852
rect 22824 10908 22888 10912
rect 22824 10852 22828 10908
rect 22828 10852 22884 10908
rect 22884 10852 22888 10908
rect 22824 10848 22888 10852
rect 22904 10908 22968 10912
rect 22904 10852 22908 10908
rect 22908 10852 22964 10908
rect 22964 10852 22968 10908
rect 22904 10848 22968 10852
rect 3666 10364 3730 10368
rect 3666 10308 3670 10364
rect 3670 10308 3726 10364
rect 3726 10308 3730 10364
rect 3666 10304 3730 10308
rect 3746 10364 3810 10368
rect 3746 10308 3750 10364
rect 3750 10308 3806 10364
rect 3806 10308 3810 10364
rect 3746 10304 3810 10308
rect 3826 10364 3890 10368
rect 3826 10308 3830 10364
rect 3830 10308 3886 10364
rect 3886 10308 3890 10364
rect 3826 10304 3890 10308
rect 3906 10364 3970 10368
rect 3906 10308 3910 10364
rect 3910 10308 3966 10364
rect 3966 10308 3970 10364
rect 3906 10304 3970 10308
rect 9094 10364 9158 10368
rect 9094 10308 9098 10364
rect 9098 10308 9154 10364
rect 9154 10308 9158 10364
rect 9094 10304 9158 10308
rect 9174 10364 9238 10368
rect 9174 10308 9178 10364
rect 9178 10308 9234 10364
rect 9234 10308 9238 10364
rect 9174 10304 9238 10308
rect 9254 10364 9318 10368
rect 9254 10308 9258 10364
rect 9258 10308 9314 10364
rect 9314 10308 9318 10364
rect 9254 10304 9318 10308
rect 9334 10364 9398 10368
rect 9334 10308 9338 10364
rect 9338 10308 9394 10364
rect 9394 10308 9398 10364
rect 9334 10304 9398 10308
rect 14522 10364 14586 10368
rect 14522 10308 14526 10364
rect 14526 10308 14582 10364
rect 14582 10308 14586 10364
rect 14522 10304 14586 10308
rect 14602 10364 14666 10368
rect 14602 10308 14606 10364
rect 14606 10308 14662 10364
rect 14662 10308 14666 10364
rect 14602 10304 14666 10308
rect 14682 10364 14746 10368
rect 14682 10308 14686 10364
rect 14686 10308 14742 10364
rect 14742 10308 14746 10364
rect 14682 10304 14746 10308
rect 14762 10364 14826 10368
rect 14762 10308 14766 10364
rect 14766 10308 14822 10364
rect 14822 10308 14826 10364
rect 14762 10304 14826 10308
rect 19950 10364 20014 10368
rect 19950 10308 19954 10364
rect 19954 10308 20010 10364
rect 20010 10308 20014 10364
rect 19950 10304 20014 10308
rect 20030 10364 20094 10368
rect 20030 10308 20034 10364
rect 20034 10308 20090 10364
rect 20090 10308 20094 10364
rect 20030 10304 20094 10308
rect 20110 10364 20174 10368
rect 20110 10308 20114 10364
rect 20114 10308 20170 10364
rect 20170 10308 20174 10364
rect 20110 10304 20174 10308
rect 20190 10364 20254 10368
rect 20190 10308 20194 10364
rect 20194 10308 20250 10364
rect 20250 10308 20254 10364
rect 20190 10304 20254 10308
rect 6380 9820 6444 9824
rect 6380 9764 6384 9820
rect 6384 9764 6440 9820
rect 6440 9764 6444 9820
rect 6380 9760 6444 9764
rect 6460 9820 6524 9824
rect 6460 9764 6464 9820
rect 6464 9764 6520 9820
rect 6520 9764 6524 9820
rect 6460 9760 6524 9764
rect 6540 9820 6604 9824
rect 6540 9764 6544 9820
rect 6544 9764 6600 9820
rect 6600 9764 6604 9820
rect 6540 9760 6604 9764
rect 6620 9820 6684 9824
rect 6620 9764 6624 9820
rect 6624 9764 6680 9820
rect 6680 9764 6684 9820
rect 6620 9760 6684 9764
rect 11808 9820 11872 9824
rect 11808 9764 11812 9820
rect 11812 9764 11868 9820
rect 11868 9764 11872 9820
rect 11808 9760 11872 9764
rect 11888 9820 11952 9824
rect 11888 9764 11892 9820
rect 11892 9764 11948 9820
rect 11948 9764 11952 9820
rect 11888 9760 11952 9764
rect 11968 9820 12032 9824
rect 11968 9764 11972 9820
rect 11972 9764 12028 9820
rect 12028 9764 12032 9820
rect 11968 9760 12032 9764
rect 12048 9820 12112 9824
rect 12048 9764 12052 9820
rect 12052 9764 12108 9820
rect 12108 9764 12112 9820
rect 12048 9760 12112 9764
rect 17236 9820 17300 9824
rect 17236 9764 17240 9820
rect 17240 9764 17296 9820
rect 17296 9764 17300 9820
rect 17236 9760 17300 9764
rect 17316 9820 17380 9824
rect 17316 9764 17320 9820
rect 17320 9764 17376 9820
rect 17376 9764 17380 9820
rect 17316 9760 17380 9764
rect 17396 9820 17460 9824
rect 17396 9764 17400 9820
rect 17400 9764 17456 9820
rect 17456 9764 17460 9820
rect 17396 9760 17460 9764
rect 17476 9820 17540 9824
rect 17476 9764 17480 9820
rect 17480 9764 17536 9820
rect 17536 9764 17540 9820
rect 17476 9760 17540 9764
rect 22664 9820 22728 9824
rect 22664 9764 22668 9820
rect 22668 9764 22724 9820
rect 22724 9764 22728 9820
rect 22664 9760 22728 9764
rect 22744 9820 22808 9824
rect 22744 9764 22748 9820
rect 22748 9764 22804 9820
rect 22804 9764 22808 9820
rect 22744 9760 22808 9764
rect 22824 9820 22888 9824
rect 22824 9764 22828 9820
rect 22828 9764 22884 9820
rect 22884 9764 22888 9820
rect 22824 9760 22888 9764
rect 22904 9820 22968 9824
rect 22904 9764 22908 9820
rect 22908 9764 22964 9820
rect 22964 9764 22968 9820
rect 22904 9760 22968 9764
rect 3666 9276 3730 9280
rect 3666 9220 3670 9276
rect 3670 9220 3726 9276
rect 3726 9220 3730 9276
rect 3666 9216 3730 9220
rect 3746 9276 3810 9280
rect 3746 9220 3750 9276
rect 3750 9220 3806 9276
rect 3806 9220 3810 9276
rect 3746 9216 3810 9220
rect 3826 9276 3890 9280
rect 3826 9220 3830 9276
rect 3830 9220 3886 9276
rect 3886 9220 3890 9276
rect 3826 9216 3890 9220
rect 3906 9276 3970 9280
rect 3906 9220 3910 9276
rect 3910 9220 3966 9276
rect 3966 9220 3970 9276
rect 3906 9216 3970 9220
rect 9094 9276 9158 9280
rect 9094 9220 9098 9276
rect 9098 9220 9154 9276
rect 9154 9220 9158 9276
rect 9094 9216 9158 9220
rect 9174 9276 9238 9280
rect 9174 9220 9178 9276
rect 9178 9220 9234 9276
rect 9234 9220 9238 9276
rect 9174 9216 9238 9220
rect 9254 9276 9318 9280
rect 9254 9220 9258 9276
rect 9258 9220 9314 9276
rect 9314 9220 9318 9276
rect 9254 9216 9318 9220
rect 9334 9276 9398 9280
rect 9334 9220 9338 9276
rect 9338 9220 9394 9276
rect 9394 9220 9398 9276
rect 9334 9216 9398 9220
rect 14522 9276 14586 9280
rect 14522 9220 14526 9276
rect 14526 9220 14582 9276
rect 14582 9220 14586 9276
rect 14522 9216 14586 9220
rect 14602 9276 14666 9280
rect 14602 9220 14606 9276
rect 14606 9220 14662 9276
rect 14662 9220 14666 9276
rect 14602 9216 14666 9220
rect 14682 9276 14746 9280
rect 14682 9220 14686 9276
rect 14686 9220 14742 9276
rect 14742 9220 14746 9276
rect 14682 9216 14746 9220
rect 14762 9276 14826 9280
rect 14762 9220 14766 9276
rect 14766 9220 14822 9276
rect 14822 9220 14826 9276
rect 14762 9216 14826 9220
rect 19950 9276 20014 9280
rect 19950 9220 19954 9276
rect 19954 9220 20010 9276
rect 20010 9220 20014 9276
rect 19950 9216 20014 9220
rect 20030 9276 20094 9280
rect 20030 9220 20034 9276
rect 20034 9220 20090 9276
rect 20090 9220 20094 9276
rect 20030 9216 20094 9220
rect 20110 9276 20174 9280
rect 20110 9220 20114 9276
rect 20114 9220 20170 9276
rect 20170 9220 20174 9276
rect 20110 9216 20174 9220
rect 20190 9276 20254 9280
rect 20190 9220 20194 9276
rect 20194 9220 20250 9276
rect 20250 9220 20254 9276
rect 20190 9216 20254 9220
rect 6380 8732 6444 8736
rect 6380 8676 6384 8732
rect 6384 8676 6440 8732
rect 6440 8676 6444 8732
rect 6380 8672 6444 8676
rect 6460 8732 6524 8736
rect 6460 8676 6464 8732
rect 6464 8676 6520 8732
rect 6520 8676 6524 8732
rect 6460 8672 6524 8676
rect 6540 8732 6604 8736
rect 6540 8676 6544 8732
rect 6544 8676 6600 8732
rect 6600 8676 6604 8732
rect 6540 8672 6604 8676
rect 6620 8732 6684 8736
rect 6620 8676 6624 8732
rect 6624 8676 6680 8732
rect 6680 8676 6684 8732
rect 6620 8672 6684 8676
rect 11808 8732 11872 8736
rect 11808 8676 11812 8732
rect 11812 8676 11868 8732
rect 11868 8676 11872 8732
rect 11808 8672 11872 8676
rect 11888 8732 11952 8736
rect 11888 8676 11892 8732
rect 11892 8676 11948 8732
rect 11948 8676 11952 8732
rect 11888 8672 11952 8676
rect 11968 8732 12032 8736
rect 11968 8676 11972 8732
rect 11972 8676 12028 8732
rect 12028 8676 12032 8732
rect 11968 8672 12032 8676
rect 12048 8732 12112 8736
rect 12048 8676 12052 8732
rect 12052 8676 12108 8732
rect 12108 8676 12112 8732
rect 12048 8672 12112 8676
rect 17236 8732 17300 8736
rect 17236 8676 17240 8732
rect 17240 8676 17296 8732
rect 17296 8676 17300 8732
rect 17236 8672 17300 8676
rect 17316 8732 17380 8736
rect 17316 8676 17320 8732
rect 17320 8676 17376 8732
rect 17376 8676 17380 8732
rect 17316 8672 17380 8676
rect 17396 8732 17460 8736
rect 17396 8676 17400 8732
rect 17400 8676 17456 8732
rect 17456 8676 17460 8732
rect 17396 8672 17460 8676
rect 17476 8732 17540 8736
rect 17476 8676 17480 8732
rect 17480 8676 17536 8732
rect 17536 8676 17540 8732
rect 17476 8672 17540 8676
rect 22664 8732 22728 8736
rect 22664 8676 22668 8732
rect 22668 8676 22724 8732
rect 22724 8676 22728 8732
rect 22664 8672 22728 8676
rect 22744 8732 22808 8736
rect 22744 8676 22748 8732
rect 22748 8676 22804 8732
rect 22804 8676 22808 8732
rect 22744 8672 22808 8676
rect 22824 8732 22888 8736
rect 22824 8676 22828 8732
rect 22828 8676 22884 8732
rect 22884 8676 22888 8732
rect 22824 8672 22888 8676
rect 22904 8732 22968 8736
rect 22904 8676 22908 8732
rect 22908 8676 22964 8732
rect 22964 8676 22968 8732
rect 22904 8672 22968 8676
rect 3666 8188 3730 8192
rect 3666 8132 3670 8188
rect 3670 8132 3726 8188
rect 3726 8132 3730 8188
rect 3666 8128 3730 8132
rect 3746 8188 3810 8192
rect 3746 8132 3750 8188
rect 3750 8132 3806 8188
rect 3806 8132 3810 8188
rect 3746 8128 3810 8132
rect 3826 8188 3890 8192
rect 3826 8132 3830 8188
rect 3830 8132 3886 8188
rect 3886 8132 3890 8188
rect 3826 8128 3890 8132
rect 3906 8188 3970 8192
rect 3906 8132 3910 8188
rect 3910 8132 3966 8188
rect 3966 8132 3970 8188
rect 3906 8128 3970 8132
rect 9094 8188 9158 8192
rect 9094 8132 9098 8188
rect 9098 8132 9154 8188
rect 9154 8132 9158 8188
rect 9094 8128 9158 8132
rect 9174 8188 9238 8192
rect 9174 8132 9178 8188
rect 9178 8132 9234 8188
rect 9234 8132 9238 8188
rect 9174 8128 9238 8132
rect 9254 8188 9318 8192
rect 9254 8132 9258 8188
rect 9258 8132 9314 8188
rect 9314 8132 9318 8188
rect 9254 8128 9318 8132
rect 9334 8188 9398 8192
rect 9334 8132 9338 8188
rect 9338 8132 9394 8188
rect 9394 8132 9398 8188
rect 9334 8128 9398 8132
rect 14522 8188 14586 8192
rect 14522 8132 14526 8188
rect 14526 8132 14582 8188
rect 14582 8132 14586 8188
rect 14522 8128 14586 8132
rect 14602 8188 14666 8192
rect 14602 8132 14606 8188
rect 14606 8132 14662 8188
rect 14662 8132 14666 8188
rect 14602 8128 14666 8132
rect 14682 8188 14746 8192
rect 14682 8132 14686 8188
rect 14686 8132 14742 8188
rect 14742 8132 14746 8188
rect 14682 8128 14746 8132
rect 14762 8188 14826 8192
rect 14762 8132 14766 8188
rect 14766 8132 14822 8188
rect 14822 8132 14826 8188
rect 14762 8128 14826 8132
rect 19950 8188 20014 8192
rect 19950 8132 19954 8188
rect 19954 8132 20010 8188
rect 20010 8132 20014 8188
rect 19950 8128 20014 8132
rect 20030 8188 20094 8192
rect 20030 8132 20034 8188
rect 20034 8132 20090 8188
rect 20090 8132 20094 8188
rect 20030 8128 20094 8132
rect 20110 8188 20174 8192
rect 20110 8132 20114 8188
rect 20114 8132 20170 8188
rect 20170 8132 20174 8188
rect 20110 8128 20174 8132
rect 20190 8188 20254 8192
rect 20190 8132 20194 8188
rect 20194 8132 20250 8188
rect 20250 8132 20254 8188
rect 20190 8128 20254 8132
rect 6380 7644 6444 7648
rect 6380 7588 6384 7644
rect 6384 7588 6440 7644
rect 6440 7588 6444 7644
rect 6380 7584 6444 7588
rect 6460 7644 6524 7648
rect 6460 7588 6464 7644
rect 6464 7588 6520 7644
rect 6520 7588 6524 7644
rect 6460 7584 6524 7588
rect 6540 7644 6604 7648
rect 6540 7588 6544 7644
rect 6544 7588 6600 7644
rect 6600 7588 6604 7644
rect 6540 7584 6604 7588
rect 6620 7644 6684 7648
rect 6620 7588 6624 7644
rect 6624 7588 6680 7644
rect 6680 7588 6684 7644
rect 6620 7584 6684 7588
rect 11808 7644 11872 7648
rect 11808 7588 11812 7644
rect 11812 7588 11868 7644
rect 11868 7588 11872 7644
rect 11808 7584 11872 7588
rect 11888 7644 11952 7648
rect 11888 7588 11892 7644
rect 11892 7588 11948 7644
rect 11948 7588 11952 7644
rect 11888 7584 11952 7588
rect 11968 7644 12032 7648
rect 11968 7588 11972 7644
rect 11972 7588 12028 7644
rect 12028 7588 12032 7644
rect 11968 7584 12032 7588
rect 12048 7644 12112 7648
rect 12048 7588 12052 7644
rect 12052 7588 12108 7644
rect 12108 7588 12112 7644
rect 12048 7584 12112 7588
rect 17236 7644 17300 7648
rect 17236 7588 17240 7644
rect 17240 7588 17296 7644
rect 17296 7588 17300 7644
rect 17236 7584 17300 7588
rect 17316 7644 17380 7648
rect 17316 7588 17320 7644
rect 17320 7588 17376 7644
rect 17376 7588 17380 7644
rect 17316 7584 17380 7588
rect 17396 7644 17460 7648
rect 17396 7588 17400 7644
rect 17400 7588 17456 7644
rect 17456 7588 17460 7644
rect 17396 7584 17460 7588
rect 17476 7644 17540 7648
rect 17476 7588 17480 7644
rect 17480 7588 17536 7644
rect 17536 7588 17540 7644
rect 17476 7584 17540 7588
rect 22664 7644 22728 7648
rect 22664 7588 22668 7644
rect 22668 7588 22724 7644
rect 22724 7588 22728 7644
rect 22664 7584 22728 7588
rect 22744 7644 22808 7648
rect 22744 7588 22748 7644
rect 22748 7588 22804 7644
rect 22804 7588 22808 7644
rect 22744 7584 22808 7588
rect 22824 7644 22888 7648
rect 22824 7588 22828 7644
rect 22828 7588 22884 7644
rect 22884 7588 22888 7644
rect 22824 7584 22888 7588
rect 22904 7644 22968 7648
rect 22904 7588 22908 7644
rect 22908 7588 22964 7644
rect 22964 7588 22968 7644
rect 22904 7584 22968 7588
rect 3666 7100 3730 7104
rect 3666 7044 3670 7100
rect 3670 7044 3726 7100
rect 3726 7044 3730 7100
rect 3666 7040 3730 7044
rect 3746 7100 3810 7104
rect 3746 7044 3750 7100
rect 3750 7044 3806 7100
rect 3806 7044 3810 7100
rect 3746 7040 3810 7044
rect 3826 7100 3890 7104
rect 3826 7044 3830 7100
rect 3830 7044 3886 7100
rect 3886 7044 3890 7100
rect 3826 7040 3890 7044
rect 3906 7100 3970 7104
rect 3906 7044 3910 7100
rect 3910 7044 3966 7100
rect 3966 7044 3970 7100
rect 3906 7040 3970 7044
rect 9094 7100 9158 7104
rect 9094 7044 9098 7100
rect 9098 7044 9154 7100
rect 9154 7044 9158 7100
rect 9094 7040 9158 7044
rect 9174 7100 9238 7104
rect 9174 7044 9178 7100
rect 9178 7044 9234 7100
rect 9234 7044 9238 7100
rect 9174 7040 9238 7044
rect 9254 7100 9318 7104
rect 9254 7044 9258 7100
rect 9258 7044 9314 7100
rect 9314 7044 9318 7100
rect 9254 7040 9318 7044
rect 9334 7100 9398 7104
rect 9334 7044 9338 7100
rect 9338 7044 9394 7100
rect 9394 7044 9398 7100
rect 9334 7040 9398 7044
rect 14522 7100 14586 7104
rect 14522 7044 14526 7100
rect 14526 7044 14582 7100
rect 14582 7044 14586 7100
rect 14522 7040 14586 7044
rect 14602 7100 14666 7104
rect 14602 7044 14606 7100
rect 14606 7044 14662 7100
rect 14662 7044 14666 7100
rect 14602 7040 14666 7044
rect 14682 7100 14746 7104
rect 14682 7044 14686 7100
rect 14686 7044 14742 7100
rect 14742 7044 14746 7100
rect 14682 7040 14746 7044
rect 14762 7100 14826 7104
rect 14762 7044 14766 7100
rect 14766 7044 14822 7100
rect 14822 7044 14826 7100
rect 14762 7040 14826 7044
rect 19950 7100 20014 7104
rect 19950 7044 19954 7100
rect 19954 7044 20010 7100
rect 20010 7044 20014 7100
rect 19950 7040 20014 7044
rect 20030 7100 20094 7104
rect 20030 7044 20034 7100
rect 20034 7044 20090 7100
rect 20090 7044 20094 7100
rect 20030 7040 20094 7044
rect 20110 7100 20174 7104
rect 20110 7044 20114 7100
rect 20114 7044 20170 7100
rect 20170 7044 20174 7100
rect 20110 7040 20174 7044
rect 20190 7100 20254 7104
rect 20190 7044 20194 7100
rect 20194 7044 20250 7100
rect 20250 7044 20254 7100
rect 20190 7040 20254 7044
rect 6380 6556 6444 6560
rect 6380 6500 6384 6556
rect 6384 6500 6440 6556
rect 6440 6500 6444 6556
rect 6380 6496 6444 6500
rect 6460 6556 6524 6560
rect 6460 6500 6464 6556
rect 6464 6500 6520 6556
rect 6520 6500 6524 6556
rect 6460 6496 6524 6500
rect 6540 6556 6604 6560
rect 6540 6500 6544 6556
rect 6544 6500 6600 6556
rect 6600 6500 6604 6556
rect 6540 6496 6604 6500
rect 6620 6556 6684 6560
rect 6620 6500 6624 6556
rect 6624 6500 6680 6556
rect 6680 6500 6684 6556
rect 6620 6496 6684 6500
rect 11808 6556 11872 6560
rect 11808 6500 11812 6556
rect 11812 6500 11868 6556
rect 11868 6500 11872 6556
rect 11808 6496 11872 6500
rect 11888 6556 11952 6560
rect 11888 6500 11892 6556
rect 11892 6500 11948 6556
rect 11948 6500 11952 6556
rect 11888 6496 11952 6500
rect 11968 6556 12032 6560
rect 11968 6500 11972 6556
rect 11972 6500 12028 6556
rect 12028 6500 12032 6556
rect 11968 6496 12032 6500
rect 12048 6556 12112 6560
rect 12048 6500 12052 6556
rect 12052 6500 12108 6556
rect 12108 6500 12112 6556
rect 12048 6496 12112 6500
rect 17236 6556 17300 6560
rect 17236 6500 17240 6556
rect 17240 6500 17296 6556
rect 17296 6500 17300 6556
rect 17236 6496 17300 6500
rect 17316 6556 17380 6560
rect 17316 6500 17320 6556
rect 17320 6500 17376 6556
rect 17376 6500 17380 6556
rect 17316 6496 17380 6500
rect 17396 6556 17460 6560
rect 17396 6500 17400 6556
rect 17400 6500 17456 6556
rect 17456 6500 17460 6556
rect 17396 6496 17460 6500
rect 17476 6556 17540 6560
rect 17476 6500 17480 6556
rect 17480 6500 17536 6556
rect 17536 6500 17540 6556
rect 17476 6496 17540 6500
rect 22664 6556 22728 6560
rect 22664 6500 22668 6556
rect 22668 6500 22724 6556
rect 22724 6500 22728 6556
rect 22664 6496 22728 6500
rect 22744 6556 22808 6560
rect 22744 6500 22748 6556
rect 22748 6500 22804 6556
rect 22804 6500 22808 6556
rect 22744 6496 22808 6500
rect 22824 6556 22888 6560
rect 22824 6500 22828 6556
rect 22828 6500 22884 6556
rect 22884 6500 22888 6556
rect 22824 6496 22888 6500
rect 22904 6556 22968 6560
rect 22904 6500 22908 6556
rect 22908 6500 22964 6556
rect 22964 6500 22968 6556
rect 22904 6496 22968 6500
rect 3666 6012 3730 6016
rect 3666 5956 3670 6012
rect 3670 5956 3726 6012
rect 3726 5956 3730 6012
rect 3666 5952 3730 5956
rect 3746 6012 3810 6016
rect 3746 5956 3750 6012
rect 3750 5956 3806 6012
rect 3806 5956 3810 6012
rect 3746 5952 3810 5956
rect 3826 6012 3890 6016
rect 3826 5956 3830 6012
rect 3830 5956 3886 6012
rect 3886 5956 3890 6012
rect 3826 5952 3890 5956
rect 3906 6012 3970 6016
rect 3906 5956 3910 6012
rect 3910 5956 3966 6012
rect 3966 5956 3970 6012
rect 3906 5952 3970 5956
rect 9094 6012 9158 6016
rect 9094 5956 9098 6012
rect 9098 5956 9154 6012
rect 9154 5956 9158 6012
rect 9094 5952 9158 5956
rect 9174 6012 9238 6016
rect 9174 5956 9178 6012
rect 9178 5956 9234 6012
rect 9234 5956 9238 6012
rect 9174 5952 9238 5956
rect 9254 6012 9318 6016
rect 9254 5956 9258 6012
rect 9258 5956 9314 6012
rect 9314 5956 9318 6012
rect 9254 5952 9318 5956
rect 9334 6012 9398 6016
rect 9334 5956 9338 6012
rect 9338 5956 9394 6012
rect 9394 5956 9398 6012
rect 9334 5952 9398 5956
rect 14522 6012 14586 6016
rect 14522 5956 14526 6012
rect 14526 5956 14582 6012
rect 14582 5956 14586 6012
rect 14522 5952 14586 5956
rect 14602 6012 14666 6016
rect 14602 5956 14606 6012
rect 14606 5956 14662 6012
rect 14662 5956 14666 6012
rect 14602 5952 14666 5956
rect 14682 6012 14746 6016
rect 14682 5956 14686 6012
rect 14686 5956 14742 6012
rect 14742 5956 14746 6012
rect 14682 5952 14746 5956
rect 14762 6012 14826 6016
rect 14762 5956 14766 6012
rect 14766 5956 14822 6012
rect 14822 5956 14826 6012
rect 14762 5952 14826 5956
rect 19950 6012 20014 6016
rect 19950 5956 19954 6012
rect 19954 5956 20010 6012
rect 20010 5956 20014 6012
rect 19950 5952 20014 5956
rect 20030 6012 20094 6016
rect 20030 5956 20034 6012
rect 20034 5956 20090 6012
rect 20090 5956 20094 6012
rect 20030 5952 20094 5956
rect 20110 6012 20174 6016
rect 20110 5956 20114 6012
rect 20114 5956 20170 6012
rect 20170 5956 20174 6012
rect 20110 5952 20174 5956
rect 20190 6012 20254 6016
rect 20190 5956 20194 6012
rect 20194 5956 20250 6012
rect 20250 5956 20254 6012
rect 20190 5952 20254 5956
rect 6380 5468 6444 5472
rect 6380 5412 6384 5468
rect 6384 5412 6440 5468
rect 6440 5412 6444 5468
rect 6380 5408 6444 5412
rect 6460 5468 6524 5472
rect 6460 5412 6464 5468
rect 6464 5412 6520 5468
rect 6520 5412 6524 5468
rect 6460 5408 6524 5412
rect 6540 5468 6604 5472
rect 6540 5412 6544 5468
rect 6544 5412 6600 5468
rect 6600 5412 6604 5468
rect 6540 5408 6604 5412
rect 6620 5468 6684 5472
rect 6620 5412 6624 5468
rect 6624 5412 6680 5468
rect 6680 5412 6684 5468
rect 6620 5408 6684 5412
rect 11808 5468 11872 5472
rect 11808 5412 11812 5468
rect 11812 5412 11868 5468
rect 11868 5412 11872 5468
rect 11808 5408 11872 5412
rect 11888 5468 11952 5472
rect 11888 5412 11892 5468
rect 11892 5412 11948 5468
rect 11948 5412 11952 5468
rect 11888 5408 11952 5412
rect 11968 5468 12032 5472
rect 11968 5412 11972 5468
rect 11972 5412 12028 5468
rect 12028 5412 12032 5468
rect 11968 5408 12032 5412
rect 12048 5468 12112 5472
rect 12048 5412 12052 5468
rect 12052 5412 12108 5468
rect 12108 5412 12112 5468
rect 12048 5408 12112 5412
rect 17236 5468 17300 5472
rect 17236 5412 17240 5468
rect 17240 5412 17296 5468
rect 17296 5412 17300 5468
rect 17236 5408 17300 5412
rect 17316 5468 17380 5472
rect 17316 5412 17320 5468
rect 17320 5412 17376 5468
rect 17376 5412 17380 5468
rect 17316 5408 17380 5412
rect 17396 5468 17460 5472
rect 17396 5412 17400 5468
rect 17400 5412 17456 5468
rect 17456 5412 17460 5468
rect 17396 5408 17460 5412
rect 17476 5468 17540 5472
rect 17476 5412 17480 5468
rect 17480 5412 17536 5468
rect 17536 5412 17540 5468
rect 17476 5408 17540 5412
rect 22664 5468 22728 5472
rect 22664 5412 22668 5468
rect 22668 5412 22724 5468
rect 22724 5412 22728 5468
rect 22664 5408 22728 5412
rect 22744 5468 22808 5472
rect 22744 5412 22748 5468
rect 22748 5412 22804 5468
rect 22804 5412 22808 5468
rect 22744 5408 22808 5412
rect 22824 5468 22888 5472
rect 22824 5412 22828 5468
rect 22828 5412 22884 5468
rect 22884 5412 22888 5468
rect 22824 5408 22888 5412
rect 22904 5468 22968 5472
rect 22904 5412 22908 5468
rect 22908 5412 22964 5468
rect 22964 5412 22968 5468
rect 22904 5408 22968 5412
rect 3666 4924 3730 4928
rect 3666 4868 3670 4924
rect 3670 4868 3726 4924
rect 3726 4868 3730 4924
rect 3666 4864 3730 4868
rect 3746 4924 3810 4928
rect 3746 4868 3750 4924
rect 3750 4868 3806 4924
rect 3806 4868 3810 4924
rect 3746 4864 3810 4868
rect 3826 4924 3890 4928
rect 3826 4868 3830 4924
rect 3830 4868 3886 4924
rect 3886 4868 3890 4924
rect 3826 4864 3890 4868
rect 3906 4924 3970 4928
rect 3906 4868 3910 4924
rect 3910 4868 3966 4924
rect 3966 4868 3970 4924
rect 3906 4864 3970 4868
rect 9094 4924 9158 4928
rect 9094 4868 9098 4924
rect 9098 4868 9154 4924
rect 9154 4868 9158 4924
rect 9094 4864 9158 4868
rect 9174 4924 9238 4928
rect 9174 4868 9178 4924
rect 9178 4868 9234 4924
rect 9234 4868 9238 4924
rect 9174 4864 9238 4868
rect 9254 4924 9318 4928
rect 9254 4868 9258 4924
rect 9258 4868 9314 4924
rect 9314 4868 9318 4924
rect 9254 4864 9318 4868
rect 9334 4924 9398 4928
rect 9334 4868 9338 4924
rect 9338 4868 9394 4924
rect 9394 4868 9398 4924
rect 9334 4864 9398 4868
rect 14522 4924 14586 4928
rect 14522 4868 14526 4924
rect 14526 4868 14582 4924
rect 14582 4868 14586 4924
rect 14522 4864 14586 4868
rect 14602 4924 14666 4928
rect 14602 4868 14606 4924
rect 14606 4868 14662 4924
rect 14662 4868 14666 4924
rect 14602 4864 14666 4868
rect 14682 4924 14746 4928
rect 14682 4868 14686 4924
rect 14686 4868 14742 4924
rect 14742 4868 14746 4924
rect 14682 4864 14746 4868
rect 14762 4924 14826 4928
rect 14762 4868 14766 4924
rect 14766 4868 14822 4924
rect 14822 4868 14826 4924
rect 14762 4864 14826 4868
rect 19950 4924 20014 4928
rect 19950 4868 19954 4924
rect 19954 4868 20010 4924
rect 20010 4868 20014 4924
rect 19950 4864 20014 4868
rect 20030 4924 20094 4928
rect 20030 4868 20034 4924
rect 20034 4868 20090 4924
rect 20090 4868 20094 4924
rect 20030 4864 20094 4868
rect 20110 4924 20174 4928
rect 20110 4868 20114 4924
rect 20114 4868 20170 4924
rect 20170 4868 20174 4924
rect 20110 4864 20174 4868
rect 20190 4924 20254 4928
rect 20190 4868 20194 4924
rect 20194 4868 20250 4924
rect 20250 4868 20254 4924
rect 20190 4864 20254 4868
rect 6380 4380 6444 4384
rect 6380 4324 6384 4380
rect 6384 4324 6440 4380
rect 6440 4324 6444 4380
rect 6380 4320 6444 4324
rect 6460 4380 6524 4384
rect 6460 4324 6464 4380
rect 6464 4324 6520 4380
rect 6520 4324 6524 4380
rect 6460 4320 6524 4324
rect 6540 4380 6604 4384
rect 6540 4324 6544 4380
rect 6544 4324 6600 4380
rect 6600 4324 6604 4380
rect 6540 4320 6604 4324
rect 6620 4380 6684 4384
rect 6620 4324 6624 4380
rect 6624 4324 6680 4380
rect 6680 4324 6684 4380
rect 6620 4320 6684 4324
rect 11808 4380 11872 4384
rect 11808 4324 11812 4380
rect 11812 4324 11868 4380
rect 11868 4324 11872 4380
rect 11808 4320 11872 4324
rect 11888 4380 11952 4384
rect 11888 4324 11892 4380
rect 11892 4324 11948 4380
rect 11948 4324 11952 4380
rect 11888 4320 11952 4324
rect 11968 4380 12032 4384
rect 11968 4324 11972 4380
rect 11972 4324 12028 4380
rect 12028 4324 12032 4380
rect 11968 4320 12032 4324
rect 12048 4380 12112 4384
rect 12048 4324 12052 4380
rect 12052 4324 12108 4380
rect 12108 4324 12112 4380
rect 12048 4320 12112 4324
rect 17236 4380 17300 4384
rect 17236 4324 17240 4380
rect 17240 4324 17296 4380
rect 17296 4324 17300 4380
rect 17236 4320 17300 4324
rect 17316 4380 17380 4384
rect 17316 4324 17320 4380
rect 17320 4324 17376 4380
rect 17376 4324 17380 4380
rect 17316 4320 17380 4324
rect 17396 4380 17460 4384
rect 17396 4324 17400 4380
rect 17400 4324 17456 4380
rect 17456 4324 17460 4380
rect 17396 4320 17460 4324
rect 17476 4380 17540 4384
rect 17476 4324 17480 4380
rect 17480 4324 17536 4380
rect 17536 4324 17540 4380
rect 17476 4320 17540 4324
rect 22664 4380 22728 4384
rect 22664 4324 22668 4380
rect 22668 4324 22724 4380
rect 22724 4324 22728 4380
rect 22664 4320 22728 4324
rect 22744 4380 22808 4384
rect 22744 4324 22748 4380
rect 22748 4324 22804 4380
rect 22804 4324 22808 4380
rect 22744 4320 22808 4324
rect 22824 4380 22888 4384
rect 22824 4324 22828 4380
rect 22828 4324 22884 4380
rect 22884 4324 22888 4380
rect 22824 4320 22888 4324
rect 22904 4380 22968 4384
rect 22904 4324 22908 4380
rect 22908 4324 22964 4380
rect 22964 4324 22968 4380
rect 22904 4320 22968 4324
rect 3666 3836 3730 3840
rect 3666 3780 3670 3836
rect 3670 3780 3726 3836
rect 3726 3780 3730 3836
rect 3666 3776 3730 3780
rect 3746 3836 3810 3840
rect 3746 3780 3750 3836
rect 3750 3780 3806 3836
rect 3806 3780 3810 3836
rect 3746 3776 3810 3780
rect 3826 3836 3890 3840
rect 3826 3780 3830 3836
rect 3830 3780 3886 3836
rect 3886 3780 3890 3836
rect 3826 3776 3890 3780
rect 3906 3836 3970 3840
rect 3906 3780 3910 3836
rect 3910 3780 3966 3836
rect 3966 3780 3970 3836
rect 3906 3776 3970 3780
rect 9094 3836 9158 3840
rect 9094 3780 9098 3836
rect 9098 3780 9154 3836
rect 9154 3780 9158 3836
rect 9094 3776 9158 3780
rect 9174 3836 9238 3840
rect 9174 3780 9178 3836
rect 9178 3780 9234 3836
rect 9234 3780 9238 3836
rect 9174 3776 9238 3780
rect 9254 3836 9318 3840
rect 9254 3780 9258 3836
rect 9258 3780 9314 3836
rect 9314 3780 9318 3836
rect 9254 3776 9318 3780
rect 9334 3836 9398 3840
rect 9334 3780 9338 3836
rect 9338 3780 9394 3836
rect 9394 3780 9398 3836
rect 9334 3776 9398 3780
rect 14522 3836 14586 3840
rect 14522 3780 14526 3836
rect 14526 3780 14582 3836
rect 14582 3780 14586 3836
rect 14522 3776 14586 3780
rect 14602 3836 14666 3840
rect 14602 3780 14606 3836
rect 14606 3780 14662 3836
rect 14662 3780 14666 3836
rect 14602 3776 14666 3780
rect 14682 3836 14746 3840
rect 14682 3780 14686 3836
rect 14686 3780 14742 3836
rect 14742 3780 14746 3836
rect 14682 3776 14746 3780
rect 14762 3836 14826 3840
rect 14762 3780 14766 3836
rect 14766 3780 14822 3836
rect 14822 3780 14826 3836
rect 14762 3776 14826 3780
rect 19950 3836 20014 3840
rect 19950 3780 19954 3836
rect 19954 3780 20010 3836
rect 20010 3780 20014 3836
rect 19950 3776 20014 3780
rect 20030 3836 20094 3840
rect 20030 3780 20034 3836
rect 20034 3780 20090 3836
rect 20090 3780 20094 3836
rect 20030 3776 20094 3780
rect 20110 3836 20174 3840
rect 20110 3780 20114 3836
rect 20114 3780 20170 3836
rect 20170 3780 20174 3836
rect 20110 3776 20174 3780
rect 20190 3836 20254 3840
rect 20190 3780 20194 3836
rect 20194 3780 20250 3836
rect 20250 3780 20254 3836
rect 20190 3776 20254 3780
rect 6380 3292 6444 3296
rect 6380 3236 6384 3292
rect 6384 3236 6440 3292
rect 6440 3236 6444 3292
rect 6380 3232 6444 3236
rect 6460 3292 6524 3296
rect 6460 3236 6464 3292
rect 6464 3236 6520 3292
rect 6520 3236 6524 3292
rect 6460 3232 6524 3236
rect 6540 3292 6604 3296
rect 6540 3236 6544 3292
rect 6544 3236 6600 3292
rect 6600 3236 6604 3292
rect 6540 3232 6604 3236
rect 6620 3292 6684 3296
rect 6620 3236 6624 3292
rect 6624 3236 6680 3292
rect 6680 3236 6684 3292
rect 6620 3232 6684 3236
rect 11808 3292 11872 3296
rect 11808 3236 11812 3292
rect 11812 3236 11868 3292
rect 11868 3236 11872 3292
rect 11808 3232 11872 3236
rect 11888 3292 11952 3296
rect 11888 3236 11892 3292
rect 11892 3236 11948 3292
rect 11948 3236 11952 3292
rect 11888 3232 11952 3236
rect 11968 3292 12032 3296
rect 11968 3236 11972 3292
rect 11972 3236 12028 3292
rect 12028 3236 12032 3292
rect 11968 3232 12032 3236
rect 12048 3292 12112 3296
rect 12048 3236 12052 3292
rect 12052 3236 12108 3292
rect 12108 3236 12112 3292
rect 12048 3232 12112 3236
rect 17236 3292 17300 3296
rect 17236 3236 17240 3292
rect 17240 3236 17296 3292
rect 17296 3236 17300 3292
rect 17236 3232 17300 3236
rect 17316 3292 17380 3296
rect 17316 3236 17320 3292
rect 17320 3236 17376 3292
rect 17376 3236 17380 3292
rect 17316 3232 17380 3236
rect 17396 3292 17460 3296
rect 17396 3236 17400 3292
rect 17400 3236 17456 3292
rect 17456 3236 17460 3292
rect 17396 3232 17460 3236
rect 17476 3292 17540 3296
rect 17476 3236 17480 3292
rect 17480 3236 17536 3292
rect 17536 3236 17540 3292
rect 17476 3232 17540 3236
rect 22664 3292 22728 3296
rect 22664 3236 22668 3292
rect 22668 3236 22724 3292
rect 22724 3236 22728 3292
rect 22664 3232 22728 3236
rect 22744 3292 22808 3296
rect 22744 3236 22748 3292
rect 22748 3236 22804 3292
rect 22804 3236 22808 3292
rect 22744 3232 22808 3236
rect 22824 3292 22888 3296
rect 22824 3236 22828 3292
rect 22828 3236 22884 3292
rect 22884 3236 22888 3292
rect 22824 3232 22888 3236
rect 22904 3292 22968 3296
rect 22904 3236 22908 3292
rect 22908 3236 22964 3292
rect 22964 3236 22968 3292
rect 22904 3232 22968 3236
rect 3666 2748 3730 2752
rect 3666 2692 3670 2748
rect 3670 2692 3726 2748
rect 3726 2692 3730 2748
rect 3666 2688 3730 2692
rect 3746 2748 3810 2752
rect 3746 2692 3750 2748
rect 3750 2692 3806 2748
rect 3806 2692 3810 2748
rect 3746 2688 3810 2692
rect 3826 2748 3890 2752
rect 3826 2692 3830 2748
rect 3830 2692 3886 2748
rect 3886 2692 3890 2748
rect 3826 2688 3890 2692
rect 3906 2748 3970 2752
rect 3906 2692 3910 2748
rect 3910 2692 3966 2748
rect 3966 2692 3970 2748
rect 3906 2688 3970 2692
rect 9094 2748 9158 2752
rect 9094 2692 9098 2748
rect 9098 2692 9154 2748
rect 9154 2692 9158 2748
rect 9094 2688 9158 2692
rect 9174 2748 9238 2752
rect 9174 2692 9178 2748
rect 9178 2692 9234 2748
rect 9234 2692 9238 2748
rect 9174 2688 9238 2692
rect 9254 2748 9318 2752
rect 9254 2692 9258 2748
rect 9258 2692 9314 2748
rect 9314 2692 9318 2748
rect 9254 2688 9318 2692
rect 9334 2748 9398 2752
rect 9334 2692 9338 2748
rect 9338 2692 9394 2748
rect 9394 2692 9398 2748
rect 9334 2688 9398 2692
rect 14522 2748 14586 2752
rect 14522 2692 14526 2748
rect 14526 2692 14582 2748
rect 14582 2692 14586 2748
rect 14522 2688 14586 2692
rect 14602 2748 14666 2752
rect 14602 2692 14606 2748
rect 14606 2692 14662 2748
rect 14662 2692 14666 2748
rect 14602 2688 14666 2692
rect 14682 2748 14746 2752
rect 14682 2692 14686 2748
rect 14686 2692 14742 2748
rect 14742 2692 14746 2748
rect 14682 2688 14746 2692
rect 14762 2748 14826 2752
rect 14762 2692 14766 2748
rect 14766 2692 14822 2748
rect 14822 2692 14826 2748
rect 14762 2688 14826 2692
rect 19950 2748 20014 2752
rect 19950 2692 19954 2748
rect 19954 2692 20010 2748
rect 20010 2692 20014 2748
rect 19950 2688 20014 2692
rect 20030 2748 20094 2752
rect 20030 2692 20034 2748
rect 20034 2692 20090 2748
rect 20090 2692 20094 2748
rect 20030 2688 20094 2692
rect 20110 2748 20174 2752
rect 20110 2692 20114 2748
rect 20114 2692 20170 2748
rect 20170 2692 20174 2748
rect 20110 2688 20174 2692
rect 20190 2748 20254 2752
rect 20190 2692 20194 2748
rect 20194 2692 20250 2748
rect 20250 2692 20254 2748
rect 20190 2688 20254 2692
rect 6380 2204 6444 2208
rect 6380 2148 6384 2204
rect 6384 2148 6440 2204
rect 6440 2148 6444 2204
rect 6380 2144 6444 2148
rect 6460 2204 6524 2208
rect 6460 2148 6464 2204
rect 6464 2148 6520 2204
rect 6520 2148 6524 2204
rect 6460 2144 6524 2148
rect 6540 2204 6604 2208
rect 6540 2148 6544 2204
rect 6544 2148 6600 2204
rect 6600 2148 6604 2204
rect 6540 2144 6604 2148
rect 6620 2204 6684 2208
rect 6620 2148 6624 2204
rect 6624 2148 6680 2204
rect 6680 2148 6684 2204
rect 6620 2144 6684 2148
rect 11808 2204 11872 2208
rect 11808 2148 11812 2204
rect 11812 2148 11868 2204
rect 11868 2148 11872 2204
rect 11808 2144 11872 2148
rect 11888 2204 11952 2208
rect 11888 2148 11892 2204
rect 11892 2148 11948 2204
rect 11948 2148 11952 2204
rect 11888 2144 11952 2148
rect 11968 2204 12032 2208
rect 11968 2148 11972 2204
rect 11972 2148 12028 2204
rect 12028 2148 12032 2204
rect 11968 2144 12032 2148
rect 12048 2204 12112 2208
rect 12048 2148 12052 2204
rect 12052 2148 12108 2204
rect 12108 2148 12112 2204
rect 12048 2144 12112 2148
rect 17236 2204 17300 2208
rect 17236 2148 17240 2204
rect 17240 2148 17296 2204
rect 17296 2148 17300 2204
rect 17236 2144 17300 2148
rect 17316 2204 17380 2208
rect 17316 2148 17320 2204
rect 17320 2148 17376 2204
rect 17376 2148 17380 2204
rect 17316 2144 17380 2148
rect 17396 2204 17460 2208
rect 17396 2148 17400 2204
rect 17400 2148 17456 2204
rect 17456 2148 17460 2204
rect 17396 2144 17460 2148
rect 17476 2204 17540 2208
rect 17476 2148 17480 2204
rect 17480 2148 17536 2204
rect 17536 2148 17540 2204
rect 17476 2144 17540 2148
rect 22664 2204 22728 2208
rect 22664 2148 22668 2204
rect 22668 2148 22724 2204
rect 22724 2148 22728 2204
rect 22664 2144 22728 2148
rect 22744 2204 22808 2208
rect 22744 2148 22748 2204
rect 22748 2148 22804 2204
rect 22804 2148 22808 2204
rect 22744 2144 22808 2148
rect 22824 2204 22888 2208
rect 22824 2148 22828 2204
rect 22828 2148 22884 2204
rect 22884 2148 22888 2204
rect 22824 2144 22888 2148
rect 22904 2204 22968 2208
rect 22904 2148 22908 2204
rect 22908 2148 22964 2204
rect 22964 2148 22968 2204
rect 22904 2144 22968 2148
<< metal4 >>
rect 3658 21248 3978 21808
rect 3658 21184 3666 21248
rect 3730 21184 3746 21248
rect 3810 21184 3826 21248
rect 3890 21184 3906 21248
rect 3970 21184 3978 21248
rect 3658 20160 3978 21184
rect 3658 20096 3666 20160
rect 3730 20096 3746 20160
rect 3810 20096 3826 20160
rect 3890 20096 3906 20160
rect 3970 20096 3978 20160
rect 3658 19072 3978 20096
rect 3658 19008 3666 19072
rect 3730 19008 3746 19072
rect 3810 19008 3826 19072
rect 3890 19008 3906 19072
rect 3970 19008 3978 19072
rect 3658 17984 3978 19008
rect 3658 17920 3666 17984
rect 3730 17920 3746 17984
rect 3810 17920 3826 17984
rect 3890 17920 3906 17984
rect 3970 17920 3978 17984
rect 3658 16896 3978 17920
rect 3658 16832 3666 16896
rect 3730 16832 3746 16896
rect 3810 16832 3826 16896
rect 3890 16832 3906 16896
rect 3970 16832 3978 16896
rect 3658 15808 3978 16832
rect 3658 15744 3666 15808
rect 3730 15744 3746 15808
rect 3810 15744 3826 15808
rect 3890 15744 3906 15808
rect 3970 15744 3978 15808
rect 3658 14720 3978 15744
rect 3658 14656 3666 14720
rect 3730 14656 3746 14720
rect 3810 14656 3826 14720
rect 3890 14656 3906 14720
rect 3970 14656 3978 14720
rect 3658 13632 3978 14656
rect 3658 13568 3666 13632
rect 3730 13568 3746 13632
rect 3810 13568 3826 13632
rect 3890 13568 3906 13632
rect 3970 13568 3978 13632
rect 3658 12544 3978 13568
rect 3658 12480 3666 12544
rect 3730 12480 3746 12544
rect 3810 12480 3826 12544
rect 3890 12480 3906 12544
rect 3970 12480 3978 12544
rect 3658 11456 3978 12480
rect 3658 11392 3666 11456
rect 3730 11392 3746 11456
rect 3810 11392 3826 11456
rect 3890 11392 3906 11456
rect 3970 11392 3978 11456
rect 3658 10368 3978 11392
rect 3658 10304 3666 10368
rect 3730 10304 3746 10368
rect 3810 10304 3826 10368
rect 3890 10304 3906 10368
rect 3970 10304 3978 10368
rect 3658 9280 3978 10304
rect 3658 9216 3666 9280
rect 3730 9216 3746 9280
rect 3810 9216 3826 9280
rect 3890 9216 3906 9280
rect 3970 9216 3978 9280
rect 3658 8192 3978 9216
rect 3658 8128 3666 8192
rect 3730 8128 3746 8192
rect 3810 8128 3826 8192
rect 3890 8128 3906 8192
rect 3970 8128 3978 8192
rect 3658 7104 3978 8128
rect 3658 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3978 7104
rect 3658 6016 3978 7040
rect 3658 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3978 6016
rect 3658 4928 3978 5952
rect 3658 4864 3666 4928
rect 3730 4864 3746 4928
rect 3810 4864 3826 4928
rect 3890 4864 3906 4928
rect 3970 4864 3978 4928
rect 3658 3840 3978 4864
rect 3658 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3978 3840
rect 3658 2752 3978 3776
rect 3658 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3978 2752
rect 3658 2128 3978 2688
rect 6372 21792 6692 21808
rect 6372 21728 6380 21792
rect 6444 21728 6460 21792
rect 6524 21728 6540 21792
rect 6604 21728 6620 21792
rect 6684 21728 6692 21792
rect 6372 20704 6692 21728
rect 6372 20640 6380 20704
rect 6444 20640 6460 20704
rect 6524 20640 6540 20704
rect 6604 20640 6620 20704
rect 6684 20640 6692 20704
rect 6372 19616 6692 20640
rect 6372 19552 6380 19616
rect 6444 19552 6460 19616
rect 6524 19552 6540 19616
rect 6604 19552 6620 19616
rect 6684 19552 6692 19616
rect 6372 18528 6692 19552
rect 6372 18464 6380 18528
rect 6444 18464 6460 18528
rect 6524 18464 6540 18528
rect 6604 18464 6620 18528
rect 6684 18464 6692 18528
rect 6372 17440 6692 18464
rect 6372 17376 6380 17440
rect 6444 17376 6460 17440
rect 6524 17376 6540 17440
rect 6604 17376 6620 17440
rect 6684 17376 6692 17440
rect 6372 16352 6692 17376
rect 6372 16288 6380 16352
rect 6444 16288 6460 16352
rect 6524 16288 6540 16352
rect 6604 16288 6620 16352
rect 6684 16288 6692 16352
rect 6372 15264 6692 16288
rect 6372 15200 6380 15264
rect 6444 15200 6460 15264
rect 6524 15200 6540 15264
rect 6604 15200 6620 15264
rect 6684 15200 6692 15264
rect 6372 14176 6692 15200
rect 6372 14112 6380 14176
rect 6444 14112 6460 14176
rect 6524 14112 6540 14176
rect 6604 14112 6620 14176
rect 6684 14112 6692 14176
rect 6372 13088 6692 14112
rect 6372 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6692 13088
rect 6372 12000 6692 13024
rect 6372 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6692 12000
rect 6372 10912 6692 11936
rect 6372 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6692 10912
rect 6372 9824 6692 10848
rect 6372 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6692 9824
rect 6372 8736 6692 9760
rect 6372 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6692 8736
rect 6372 7648 6692 8672
rect 6372 7584 6380 7648
rect 6444 7584 6460 7648
rect 6524 7584 6540 7648
rect 6604 7584 6620 7648
rect 6684 7584 6692 7648
rect 6372 6560 6692 7584
rect 6372 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6692 6560
rect 6372 5472 6692 6496
rect 6372 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6692 5472
rect 6372 4384 6692 5408
rect 6372 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6692 4384
rect 6372 3296 6692 4320
rect 6372 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6692 3296
rect 6372 2208 6692 3232
rect 6372 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6692 2208
rect 6372 2128 6692 2144
rect 9086 21248 9406 21808
rect 9086 21184 9094 21248
rect 9158 21184 9174 21248
rect 9238 21184 9254 21248
rect 9318 21184 9334 21248
rect 9398 21184 9406 21248
rect 9086 20160 9406 21184
rect 9086 20096 9094 20160
rect 9158 20096 9174 20160
rect 9238 20096 9254 20160
rect 9318 20096 9334 20160
rect 9398 20096 9406 20160
rect 9086 19072 9406 20096
rect 9086 19008 9094 19072
rect 9158 19008 9174 19072
rect 9238 19008 9254 19072
rect 9318 19008 9334 19072
rect 9398 19008 9406 19072
rect 9086 17984 9406 19008
rect 9086 17920 9094 17984
rect 9158 17920 9174 17984
rect 9238 17920 9254 17984
rect 9318 17920 9334 17984
rect 9398 17920 9406 17984
rect 9086 16896 9406 17920
rect 9086 16832 9094 16896
rect 9158 16832 9174 16896
rect 9238 16832 9254 16896
rect 9318 16832 9334 16896
rect 9398 16832 9406 16896
rect 9086 15808 9406 16832
rect 9086 15744 9094 15808
rect 9158 15744 9174 15808
rect 9238 15744 9254 15808
rect 9318 15744 9334 15808
rect 9398 15744 9406 15808
rect 9086 14720 9406 15744
rect 9086 14656 9094 14720
rect 9158 14656 9174 14720
rect 9238 14656 9254 14720
rect 9318 14656 9334 14720
rect 9398 14656 9406 14720
rect 9086 13632 9406 14656
rect 9086 13568 9094 13632
rect 9158 13568 9174 13632
rect 9238 13568 9254 13632
rect 9318 13568 9334 13632
rect 9398 13568 9406 13632
rect 9086 12544 9406 13568
rect 9086 12480 9094 12544
rect 9158 12480 9174 12544
rect 9238 12480 9254 12544
rect 9318 12480 9334 12544
rect 9398 12480 9406 12544
rect 9086 11456 9406 12480
rect 9086 11392 9094 11456
rect 9158 11392 9174 11456
rect 9238 11392 9254 11456
rect 9318 11392 9334 11456
rect 9398 11392 9406 11456
rect 9086 10368 9406 11392
rect 9086 10304 9094 10368
rect 9158 10304 9174 10368
rect 9238 10304 9254 10368
rect 9318 10304 9334 10368
rect 9398 10304 9406 10368
rect 9086 9280 9406 10304
rect 9086 9216 9094 9280
rect 9158 9216 9174 9280
rect 9238 9216 9254 9280
rect 9318 9216 9334 9280
rect 9398 9216 9406 9280
rect 9086 8192 9406 9216
rect 9086 8128 9094 8192
rect 9158 8128 9174 8192
rect 9238 8128 9254 8192
rect 9318 8128 9334 8192
rect 9398 8128 9406 8192
rect 9086 7104 9406 8128
rect 9086 7040 9094 7104
rect 9158 7040 9174 7104
rect 9238 7040 9254 7104
rect 9318 7040 9334 7104
rect 9398 7040 9406 7104
rect 9086 6016 9406 7040
rect 9086 5952 9094 6016
rect 9158 5952 9174 6016
rect 9238 5952 9254 6016
rect 9318 5952 9334 6016
rect 9398 5952 9406 6016
rect 9086 4928 9406 5952
rect 9086 4864 9094 4928
rect 9158 4864 9174 4928
rect 9238 4864 9254 4928
rect 9318 4864 9334 4928
rect 9398 4864 9406 4928
rect 9086 3840 9406 4864
rect 9086 3776 9094 3840
rect 9158 3776 9174 3840
rect 9238 3776 9254 3840
rect 9318 3776 9334 3840
rect 9398 3776 9406 3840
rect 9086 2752 9406 3776
rect 9086 2688 9094 2752
rect 9158 2688 9174 2752
rect 9238 2688 9254 2752
rect 9318 2688 9334 2752
rect 9398 2688 9406 2752
rect 9086 2128 9406 2688
rect 11800 21792 12120 21808
rect 11800 21728 11808 21792
rect 11872 21728 11888 21792
rect 11952 21728 11968 21792
rect 12032 21728 12048 21792
rect 12112 21728 12120 21792
rect 11800 20704 12120 21728
rect 11800 20640 11808 20704
rect 11872 20640 11888 20704
rect 11952 20640 11968 20704
rect 12032 20640 12048 20704
rect 12112 20640 12120 20704
rect 11800 19616 12120 20640
rect 11800 19552 11808 19616
rect 11872 19552 11888 19616
rect 11952 19552 11968 19616
rect 12032 19552 12048 19616
rect 12112 19552 12120 19616
rect 11800 18528 12120 19552
rect 11800 18464 11808 18528
rect 11872 18464 11888 18528
rect 11952 18464 11968 18528
rect 12032 18464 12048 18528
rect 12112 18464 12120 18528
rect 11800 17440 12120 18464
rect 11800 17376 11808 17440
rect 11872 17376 11888 17440
rect 11952 17376 11968 17440
rect 12032 17376 12048 17440
rect 12112 17376 12120 17440
rect 11800 16352 12120 17376
rect 11800 16288 11808 16352
rect 11872 16288 11888 16352
rect 11952 16288 11968 16352
rect 12032 16288 12048 16352
rect 12112 16288 12120 16352
rect 11800 15264 12120 16288
rect 11800 15200 11808 15264
rect 11872 15200 11888 15264
rect 11952 15200 11968 15264
rect 12032 15200 12048 15264
rect 12112 15200 12120 15264
rect 11800 14176 12120 15200
rect 11800 14112 11808 14176
rect 11872 14112 11888 14176
rect 11952 14112 11968 14176
rect 12032 14112 12048 14176
rect 12112 14112 12120 14176
rect 11800 13088 12120 14112
rect 11800 13024 11808 13088
rect 11872 13024 11888 13088
rect 11952 13024 11968 13088
rect 12032 13024 12048 13088
rect 12112 13024 12120 13088
rect 11800 12000 12120 13024
rect 11800 11936 11808 12000
rect 11872 11936 11888 12000
rect 11952 11936 11968 12000
rect 12032 11936 12048 12000
rect 12112 11936 12120 12000
rect 11800 10912 12120 11936
rect 11800 10848 11808 10912
rect 11872 10848 11888 10912
rect 11952 10848 11968 10912
rect 12032 10848 12048 10912
rect 12112 10848 12120 10912
rect 11800 9824 12120 10848
rect 11800 9760 11808 9824
rect 11872 9760 11888 9824
rect 11952 9760 11968 9824
rect 12032 9760 12048 9824
rect 12112 9760 12120 9824
rect 11800 8736 12120 9760
rect 11800 8672 11808 8736
rect 11872 8672 11888 8736
rect 11952 8672 11968 8736
rect 12032 8672 12048 8736
rect 12112 8672 12120 8736
rect 11800 7648 12120 8672
rect 11800 7584 11808 7648
rect 11872 7584 11888 7648
rect 11952 7584 11968 7648
rect 12032 7584 12048 7648
rect 12112 7584 12120 7648
rect 11800 6560 12120 7584
rect 11800 6496 11808 6560
rect 11872 6496 11888 6560
rect 11952 6496 11968 6560
rect 12032 6496 12048 6560
rect 12112 6496 12120 6560
rect 11800 5472 12120 6496
rect 11800 5408 11808 5472
rect 11872 5408 11888 5472
rect 11952 5408 11968 5472
rect 12032 5408 12048 5472
rect 12112 5408 12120 5472
rect 11800 4384 12120 5408
rect 11800 4320 11808 4384
rect 11872 4320 11888 4384
rect 11952 4320 11968 4384
rect 12032 4320 12048 4384
rect 12112 4320 12120 4384
rect 11800 3296 12120 4320
rect 11800 3232 11808 3296
rect 11872 3232 11888 3296
rect 11952 3232 11968 3296
rect 12032 3232 12048 3296
rect 12112 3232 12120 3296
rect 11800 2208 12120 3232
rect 11800 2144 11808 2208
rect 11872 2144 11888 2208
rect 11952 2144 11968 2208
rect 12032 2144 12048 2208
rect 12112 2144 12120 2208
rect 11800 2128 12120 2144
rect 14514 21248 14834 21808
rect 14514 21184 14522 21248
rect 14586 21184 14602 21248
rect 14666 21184 14682 21248
rect 14746 21184 14762 21248
rect 14826 21184 14834 21248
rect 14514 20160 14834 21184
rect 14514 20096 14522 20160
rect 14586 20096 14602 20160
rect 14666 20096 14682 20160
rect 14746 20096 14762 20160
rect 14826 20096 14834 20160
rect 14514 19072 14834 20096
rect 14514 19008 14522 19072
rect 14586 19008 14602 19072
rect 14666 19008 14682 19072
rect 14746 19008 14762 19072
rect 14826 19008 14834 19072
rect 14514 17984 14834 19008
rect 14514 17920 14522 17984
rect 14586 17920 14602 17984
rect 14666 17920 14682 17984
rect 14746 17920 14762 17984
rect 14826 17920 14834 17984
rect 14514 16896 14834 17920
rect 14514 16832 14522 16896
rect 14586 16832 14602 16896
rect 14666 16832 14682 16896
rect 14746 16832 14762 16896
rect 14826 16832 14834 16896
rect 14514 15808 14834 16832
rect 14514 15744 14522 15808
rect 14586 15744 14602 15808
rect 14666 15744 14682 15808
rect 14746 15744 14762 15808
rect 14826 15744 14834 15808
rect 14514 14720 14834 15744
rect 14514 14656 14522 14720
rect 14586 14656 14602 14720
rect 14666 14656 14682 14720
rect 14746 14656 14762 14720
rect 14826 14656 14834 14720
rect 14514 13632 14834 14656
rect 14514 13568 14522 13632
rect 14586 13568 14602 13632
rect 14666 13568 14682 13632
rect 14746 13568 14762 13632
rect 14826 13568 14834 13632
rect 14514 12544 14834 13568
rect 14514 12480 14522 12544
rect 14586 12480 14602 12544
rect 14666 12480 14682 12544
rect 14746 12480 14762 12544
rect 14826 12480 14834 12544
rect 14514 11456 14834 12480
rect 14514 11392 14522 11456
rect 14586 11392 14602 11456
rect 14666 11392 14682 11456
rect 14746 11392 14762 11456
rect 14826 11392 14834 11456
rect 14514 10368 14834 11392
rect 14514 10304 14522 10368
rect 14586 10304 14602 10368
rect 14666 10304 14682 10368
rect 14746 10304 14762 10368
rect 14826 10304 14834 10368
rect 14514 9280 14834 10304
rect 14514 9216 14522 9280
rect 14586 9216 14602 9280
rect 14666 9216 14682 9280
rect 14746 9216 14762 9280
rect 14826 9216 14834 9280
rect 14514 8192 14834 9216
rect 14514 8128 14522 8192
rect 14586 8128 14602 8192
rect 14666 8128 14682 8192
rect 14746 8128 14762 8192
rect 14826 8128 14834 8192
rect 14514 7104 14834 8128
rect 14514 7040 14522 7104
rect 14586 7040 14602 7104
rect 14666 7040 14682 7104
rect 14746 7040 14762 7104
rect 14826 7040 14834 7104
rect 14514 6016 14834 7040
rect 14514 5952 14522 6016
rect 14586 5952 14602 6016
rect 14666 5952 14682 6016
rect 14746 5952 14762 6016
rect 14826 5952 14834 6016
rect 14514 4928 14834 5952
rect 14514 4864 14522 4928
rect 14586 4864 14602 4928
rect 14666 4864 14682 4928
rect 14746 4864 14762 4928
rect 14826 4864 14834 4928
rect 14514 3840 14834 4864
rect 14514 3776 14522 3840
rect 14586 3776 14602 3840
rect 14666 3776 14682 3840
rect 14746 3776 14762 3840
rect 14826 3776 14834 3840
rect 14514 2752 14834 3776
rect 14514 2688 14522 2752
rect 14586 2688 14602 2752
rect 14666 2688 14682 2752
rect 14746 2688 14762 2752
rect 14826 2688 14834 2752
rect 14514 2128 14834 2688
rect 17228 21792 17548 21808
rect 17228 21728 17236 21792
rect 17300 21728 17316 21792
rect 17380 21728 17396 21792
rect 17460 21728 17476 21792
rect 17540 21728 17548 21792
rect 17228 20704 17548 21728
rect 17228 20640 17236 20704
rect 17300 20640 17316 20704
rect 17380 20640 17396 20704
rect 17460 20640 17476 20704
rect 17540 20640 17548 20704
rect 17228 19616 17548 20640
rect 17228 19552 17236 19616
rect 17300 19552 17316 19616
rect 17380 19552 17396 19616
rect 17460 19552 17476 19616
rect 17540 19552 17548 19616
rect 17228 18528 17548 19552
rect 17228 18464 17236 18528
rect 17300 18464 17316 18528
rect 17380 18464 17396 18528
rect 17460 18464 17476 18528
rect 17540 18464 17548 18528
rect 17228 17440 17548 18464
rect 17228 17376 17236 17440
rect 17300 17376 17316 17440
rect 17380 17376 17396 17440
rect 17460 17376 17476 17440
rect 17540 17376 17548 17440
rect 17228 16352 17548 17376
rect 17228 16288 17236 16352
rect 17300 16288 17316 16352
rect 17380 16288 17396 16352
rect 17460 16288 17476 16352
rect 17540 16288 17548 16352
rect 17228 15264 17548 16288
rect 17228 15200 17236 15264
rect 17300 15200 17316 15264
rect 17380 15200 17396 15264
rect 17460 15200 17476 15264
rect 17540 15200 17548 15264
rect 17228 14176 17548 15200
rect 17228 14112 17236 14176
rect 17300 14112 17316 14176
rect 17380 14112 17396 14176
rect 17460 14112 17476 14176
rect 17540 14112 17548 14176
rect 17228 13088 17548 14112
rect 17228 13024 17236 13088
rect 17300 13024 17316 13088
rect 17380 13024 17396 13088
rect 17460 13024 17476 13088
rect 17540 13024 17548 13088
rect 17228 12000 17548 13024
rect 17228 11936 17236 12000
rect 17300 11936 17316 12000
rect 17380 11936 17396 12000
rect 17460 11936 17476 12000
rect 17540 11936 17548 12000
rect 17228 10912 17548 11936
rect 17228 10848 17236 10912
rect 17300 10848 17316 10912
rect 17380 10848 17396 10912
rect 17460 10848 17476 10912
rect 17540 10848 17548 10912
rect 17228 9824 17548 10848
rect 17228 9760 17236 9824
rect 17300 9760 17316 9824
rect 17380 9760 17396 9824
rect 17460 9760 17476 9824
rect 17540 9760 17548 9824
rect 17228 8736 17548 9760
rect 17228 8672 17236 8736
rect 17300 8672 17316 8736
rect 17380 8672 17396 8736
rect 17460 8672 17476 8736
rect 17540 8672 17548 8736
rect 17228 7648 17548 8672
rect 17228 7584 17236 7648
rect 17300 7584 17316 7648
rect 17380 7584 17396 7648
rect 17460 7584 17476 7648
rect 17540 7584 17548 7648
rect 17228 6560 17548 7584
rect 17228 6496 17236 6560
rect 17300 6496 17316 6560
rect 17380 6496 17396 6560
rect 17460 6496 17476 6560
rect 17540 6496 17548 6560
rect 17228 5472 17548 6496
rect 17228 5408 17236 5472
rect 17300 5408 17316 5472
rect 17380 5408 17396 5472
rect 17460 5408 17476 5472
rect 17540 5408 17548 5472
rect 17228 4384 17548 5408
rect 17228 4320 17236 4384
rect 17300 4320 17316 4384
rect 17380 4320 17396 4384
rect 17460 4320 17476 4384
rect 17540 4320 17548 4384
rect 17228 3296 17548 4320
rect 17228 3232 17236 3296
rect 17300 3232 17316 3296
rect 17380 3232 17396 3296
rect 17460 3232 17476 3296
rect 17540 3232 17548 3296
rect 17228 2208 17548 3232
rect 17228 2144 17236 2208
rect 17300 2144 17316 2208
rect 17380 2144 17396 2208
rect 17460 2144 17476 2208
rect 17540 2144 17548 2208
rect 17228 2128 17548 2144
rect 19942 21248 20262 21808
rect 19942 21184 19950 21248
rect 20014 21184 20030 21248
rect 20094 21184 20110 21248
rect 20174 21184 20190 21248
rect 20254 21184 20262 21248
rect 19942 20160 20262 21184
rect 19942 20096 19950 20160
rect 20014 20096 20030 20160
rect 20094 20096 20110 20160
rect 20174 20096 20190 20160
rect 20254 20096 20262 20160
rect 19942 19072 20262 20096
rect 19942 19008 19950 19072
rect 20014 19008 20030 19072
rect 20094 19008 20110 19072
rect 20174 19008 20190 19072
rect 20254 19008 20262 19072
rect 19942 17984 20262 19008
rect 19942 17920 19950 17984
rect 20014 17920 20030 17984
rect 20094 17920 20110 17984
rect 20174 17920 20190 17984
rect 20254 17920 20262 17984
rect 19942 16896 20262 17920
rect 19942 16832 19950 16896
rect 20014 16832 20030 16896
rect 20094 16832 20110 16896
rect 20174 16832 20190 16896
rect 20254 16832 20262 16896
rect 19942 15808 20262 16832
rect 19942 15744 19950 15808
rect 20014 15744 20030 15808
rect 20094 15744 20110 15808
rect 20174 15744 20190 15808
rect 20254 15744 20262 15808
rect 19942 14720 20262 15744
rect 19942 14656 19950 14720
rect 20014 14656 20030 14720
rect 20094 14656 20110 14720
rect 20174 14656 20190 14720
rect 20254 14656 20262 14720
rect 19942 13632 20262 14656
rect 19942 13568 19950 13632
rect 20014 13568 20030 13632
rect 20094 13568 20110 13632
rect 20174 13568 20190 13632
rect 20254 13568 20262 13632
rect 19942 12544 20262 13568
rect 19942 12480 19950 12544
rect 20014 12480 20030 12544
rect 20094 12480 20110 12544
rect 20174 12480 20190 12544
rect 20254 12480 20262 12544
rect 19942 11456 20262 12480
rect 19942 11392 19950 11456
rect 20014 11392 20030 11456
rect 20094 11392 20110 11456
rect 20174 11392 20190 11456
rect 20254 11392 20262 11456
rect 19942 10368 20262 11392
rect 19942 10304 19950 10368
rect 20014 10304 20030 10368
rect 20094 10304 20110 10368
rect 20174 10304 20190 10368
rect 20254 10304 20262 10368
rect 19942 9280 20262 10304
rect 19942 9216 19950 9280
rect 20014 9216 20030 9280
rect 20094 9216 20110 9280
rect 20174 9216 20190 9280
rect 20254 9216 20262 9280
rect 19942 8192 20262 9216
rect 19942 8128 19950 8192
rect 20014 8128 20030 8192
rect 20094 8128 20110 8192
rect 20174 8128 20190 8192
rect 20254 8128 20262 8192
rect 19942 7104 20262 8128
rect 19942 7040 19950 7104
rect 20014 7040 20030 7104
rect 20094 7040 20110 7104
rect 20174 7040 20190 7104
rect 20254 7040 20262 7104
rect 19942 6016 20262 7040
rect 19942 5952 19950 6016
rect 20014 5952 20030 6016
rect 20094 5952 20110 6016
rect 20174 5952 20190 6016
rect 20254 5952 20262 6016
rect 19942 4928 20262 5952
rect 19942 4864 19950 4928
rect 20014 4864 20030 4928
rect 20094 4864 20110 4928
rect 20174 4864 20190 4928
rect 20254 4864 20262 4928
rect 19942 3840 20262 4864
rect 19942 3776 19950 3840
rect 20014 3776 20030 3840
rect 20094 3776 20110 3840
rect 20174 3776 20190 3840
rect 20254 3776 20262 3840
rect 19942 2752 20262 3776
rect 19942 2688 19950 2752
rect 20014 2688 20030 2752
rect 20094 2688 20110 2752
rect 20174 2688 20190 2752
rect 20254 2688 20262 2752
rect 19942 2128 20262 2688
rect 22656 21792 22976 21808
rect 22656 21728 22664 21792
rect 22728 21728 22744 21792
rect 22808 21728 22824 21792
rect 22888 21728 22904 21792
rect 22968 21728 22976 21792
rect 22656 20704 22976 21728
rect 22656 20640 22664 20704
rect 22728 20640 22744 20704
rect 22808 20640 22824 20704
rect 22888 20640 22904 20704
rect 22968 20640 22976 20704
rect 22656 19616 22976 20640
rect 22656 19552 22664 19616
rect 22728 19552 22744 19616
rect 22808 19552 22824 19616
rect 22888 19552 22904 19616
rect 22968 19552 22976 19616
rect 22656 18528 22976 19552
rect 22656 18464 22664 18528
rect 22728 18464 22744 18528
rect 22808 18464 22824 18528
rect 22888 18464 22904 18528
rect 22968 18464 22976 18528
rect 22656 17440 22976 18464
rect 22656 17376 22664 17440
rect 22728 17376 22744 17440
rect 22808 17376 22824 17440
rect 22888 17376 22904 17440
rect 22968 17376 22976 17440
rect 22656 16352 22976 17376
rect 22656 16288 22664 16352
rect 22728 16288 22744 16352
rect 22808 16288 22824 16352
rect 22888 16288 22904 16352
rect 22968 16288 22976 16352
rect 22656 15264 22976 16288
rect 22656 15200 22664 15264
rect 22728 15200 22744 15264
rect 22808 15200 22824 15264
rect 22888 15200 22904 15264
rect 22968 15200 22976 15264
rect 22656 14176 22976 15200
rect 22656 14112 22664 14176
rect 22728 14112 22744 14176
rect 22808 14112 22824 14176
rect 22888 14112 22904 14176
rect 22968 14112 22976 14176
rect 22656 13088 22976 14112
rect 22656 13024 22664 13088
rect 22728 13024 22744 13088
rect 22808 13024 22824 13088
rect 22888 13024 22904 13088
rect 22968 13024 22976 13088
rect 22656 12000 22976 13024
rect 22656 11936 22664 12000
rect 22728 11936 22744 12000
rect 22808 11936 22824 12000
rect 22888 11936 22904 12000
rect 22968 11936 22976 12000
rect 22656 10912 22976 11936
rect 22656 10848 22664 10912
rect 22728 10848 22744 10912
rect 22808 10848 22824 10912
rect 22888 10848 22904 10912
rect 22968 10848 22976 10912
rect 22656 9824 22976 10848
rect 22656 9760 22664 9824
rect 22728 9760 22744 9824
rect 22808 9760 22824 9824
rect 22888 9760 22904 9824
rect 22968 9760 22976 9824
rect 22656 8736 22976 9760
rect 22656 8672 22664 8736
rect 22728 8672 22744 8736
rect 22808 8672 22824 8736
rect 22888 8672 22904 8736
rect 22968 8672 22976 8736
rect 22656 7648 22976 8672
rect 22656 7584 22664 7648
rect 22728 7584 22744 7648
rect 22808 7584 22824 7648
rect 22888 7584 22904 7648
rect 22968 7584 22976 7648
rect 22656 6560 22976 7584
rect 22656 6496 22664 6560
rect 22728 6496 22744 6560
rect 22808 6496 22824 6560
rect 22888 6496 22904 6560
rect 22968 6496 22976 6560
rect 22656 5472 22976 6496
rect 22656 5408 22664 5472
rect 22728 5408 22744 5472
rect 22808 5408 22824 5472
rect 22888 5408 22904 5472
rect 22968 5408 22976 5472
rect 22656 4384 22976 5408
rect 22656 4320 22664 4384
rect 22728 4320 22744 4384
rect 22808 4320 22824 4384
rect 22888 4320 22904 4384
rect 22968 4320 22976 4384
rect 22656 3296 22976 4320
rect 22656 3232 22664 3296
rect 22728 3232 22744 3296
rect 22808 3232 22824 3296
rect 22888 3232 22904 3296
rect 22968 3232 22976 3296
rect 22656 2208 22976 3232
rect 22656 2144 22664 2208
rect 22728 2144 22744 2208
rect 22808 2144 22824 2208
rect 22888 2144 22904 2208
rect 22968 2144 22976 2208
rect 22656 2128 22976 2144
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45
timestamp 1676037725
transform 1 0 5244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1676037725
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_177
timestamp 1676037725
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1676037725
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1676037725
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_205
timestamp 1676037725
transform 1 0 19964 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_213
timestamp 1676037725
transform 1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_159
timestamp 1676037725
transform 1 0 15732 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_37
timestamp 1676037725
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1676037725
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_64
timestamp 1676037725
transform 1 0 6992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_72
timestamp 1676037725
transform 1 0 7728 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_79
timestamp 1676037725
transform 1 0 8372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_91
timestamp 1676037725
transform 1 0 9476 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_97
timestamp 1676037725
transform 1 0 10028 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_121
timestamp 1676037725
transform 1 0 12236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_133
timestamp 1676037725
transform 1 0 13340 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_144
timestamp 1676037725
transform 1 0 14352 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_156
timestamp 1676037725
transform 1 0 15456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1676037725
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_173
timestamp 1676037725
transform 1 0 17020 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_180
timestamp 1676037725
transform 1 0 17664 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_194
timestamp 1676037725
transform 1 0 18952 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_206
timestamp 1676037725
transform 1 0 20056 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_218
timestamp 1676037725
transform 1 0 21160 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1676037725
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_39
timestamp 1676037725
transform 1 0 4692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_49
timestamp 1676037725
transform 1 0 5612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_60
timestamp 1676037725
transform 1 0 6624 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_71
timestamp 1676037725
transform 1 0 7636 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1676037725
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_100
timestamp 1676037725
transform 1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_111
timestamp 1676037725
transform 1 0 11316 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_119
timestamp 1676037725
transform 1 0 12052 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_126
timestamp 1676037725
transform 1 0 12696 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_152
timestamp 1676037725
transform 1 0 15088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_161
timestamp 1676037725
transform 1 0 15916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_168
timestamp 1676037725
transform 1 0 16560 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_180
timestamp 1676037725
transform 1 0 17664 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1676037725
transform 1 0 18676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_204
timestamp 1676037725
transform 1 0 19872 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_216
timestamp 1676037725
transform 1 0 20976 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_228
timestamp 1676037725
transform 1 0 22080 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_232
timestamp 1676037725
transform 1 0 22448 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_19
timestamp 1676037725
transform 1 0 2852 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_23
timestamp 1676037725
transform 1 0 3220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_35
timestamp 1676037725
transform 1 0 4324 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_44
timestamp 1676037725
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_64
timestamp 1676037725
transform 1 0 6992 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_75
timestamp 1676037725
transform 1 0 8004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_85
timestamp 1676037725
transform 1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_97
timestamp 1676037725
transform 1 0 10028 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_103
timestamp 1676037725
transform 1 0 10580 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_124
timestamp 1676037725
transform 1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_131
timestamp 1676037725
transform 1 0 13156 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_141
timestamp 1676037725
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_148
timestamp 1676037725
transform 1 0 14720 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_156
timestamp 1676037725
transform 1 0 15456 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 1676037725
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_184
timestamp 1676037725
transform 1 0 18032 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_192
timestamp 1676037725
transform 1 0 18768 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_202
timestamp 1676037725
transform 1 0 19688 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_214
timestamp 1676037725
transform 1 0 20792 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp 1676037725
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_37
timestamp 1676037725
transform 1 0 4508 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_49
timestamp 1676037725
transform 1 0 5612 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_61
timestamp 1676037725
transform 1 0 6716 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_72
timestamp 1676037725
transform 1 0 7728 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_126
timestamp 1676037725
transform 1 0 12696 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_130
timestamp 1676037725
transform 1 0 13064 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1676037725
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_166
timestamp 1676037725
transform 1 0 16376 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_178
timestamp 1676037725
transform 1 0 17480 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_186
timestamp 1676037725
transform 1 0 18216 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_11
timestamp 1676037725
transform 1 0 2116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_23
timestamp 1676037725
transform 1 0 3220 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_35
timestamp 1676037725
transform 1 0 4324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_47
timestamp 1676037725
transform 1 0 5428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_64
timestamp 1676037725
transform 1 0 6992 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_72
timestamp 1676037725
transform 1 0 7728 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_79
timestamp 1676037725
transform 1 0 8372 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_90
timestamp 1676037725
transform 1 0 9384 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_102
timestamp 1676037725
transform 1 0 10488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1676037725
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_119
timestamp 1676037725
transform 1 0 12052 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_131
timestamp 1676037725
transform 1 0 13156 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_139
timestamp 1676037725
transform 1 0 13892 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_151
timestamp 1676037725
transform 1 0 14996 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_157
timestamp 1676037725
transform 1 0 15548 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_198
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_210
timestamp 1676037725
transform 1 0 20424 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_14
timestamp 1676037725
transform 1 0 2392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1676037725
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_49
timestamp 1676037725
transform 1 0 5612 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1676037725
transform 1 0 6440 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_76
timestamp 1676037725
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_96
timestamp 1676037725
transform 1 0 9936 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_106
timestamp 1676037725
transform 1 0 10856 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_115
timestamp 1676037725
transform 1 0 11684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_124
timestamp 1676037725
transform 1 0 12512 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_151
timestamp 1676037725
transform 1 0 14996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_163
timestamp 1676037725
transform 1 0 16100 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_176
timestamp 1676037725
transform 1 0 17296 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_182
timestamp 1676037725
transform 1 0 17848 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_207
timestamp 1676037725
transform 1 0 20148 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_219
timestamp 1676037725
transform 1 0 21252 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_231
timestamp 1676037725
transform 1 0 22356 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1676037725
transform 1 0 1748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_12
timestamp 1676037725
transform 1 0 2208 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_22
timestamp 1676037725
transform 1 0 3128 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_30
timestamp 1676037725
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_42
timestamp 1676037725
transform 1 0 4968 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1676037725
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1676037725
transform 1 0 6808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_71
timestamp 1676037725
transform 1 0 7636 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_77
timestamp 1676037725
transform 1 0 8188 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_129
timestamp 1676037725
transform 1 0 12972 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_134
timestamp 1676037725
transform 1 0 13432 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_141
timestamp 1676037725
transform 1 0 14076 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1676037725
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_157
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1676037725
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_185
timestamp 1676037725
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_195
timestamp 1676037725
transform 1 0 19044 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_206
timestamp 1676037725
transform 1 0 20056 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1676037725
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_72
timestamp 1676037725
transform 1 0 7728 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_188
timestamp 1676037725
transform 1 0 18400 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1676037725
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_16
timestamp 1676037725
transform 1 0 2576 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_23
timestamp 1676037725
transform 1 0 3220 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_31
timestamp 1676037725
transform 1 0 3956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_50
timestamp 1676037725
transform 1 0 5704 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_77
timestamp 1676037725
transform 1 0 8188 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_94
timestamp 1676037725
transform 1 0 9752 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_106
timestamp 1676037725
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_141
timestamp 1676037725
transform 1 0 14076 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1676037725
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_157
timestamp 1676037725
transform 1 0 15548 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1676037725
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_177
timestamp 1676037725
transform 1 0 17388 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_185
timestamp 1676037725
transform 1 0 18124 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_204
timestamp 1676037725
transform 1 0 19872 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_216
timestamp 1676037725
transform 1 0 20976 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_11
timestamp 1676037725
transform 1 0 2116 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1676037725
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_50
timestamp 1676037725
transform 1 0 5704 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_56
timestamp 1676037725
transform 1 0 6256 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_73
timestamp 1676037725
transform 1 0 7820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp 1676037725
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_107
timestamp 1676037725
transform 1 0 10948 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_128
timestamp 1676037725
transform 1 0 12880 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_159
timestamp 1676037725
transform 1 0 15732 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_172
timestamp 1676037725
transform 1 0 16928 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_184
timestamp 1676037725
transform 1 0 18032 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_208
timestamp 1676037725
transform 1 0 20240 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_220
timestamp 1676037725
transform 1 0 21344 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_232
timestamp 1676037725
transform 1 0 22448 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1676037725
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_73
timestamp 1676037725
transform 1 0 7820 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_90
timestamp 1676037725
transform 1 0 9384 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_141
timestamp 1676037725
transform 1 0 14076 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_153
timestamp 1676037725
transform 1 0 15180 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_163
timestamp 1676037725
transform 1 0 16100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_198
timestamp 1676037725
transform 1 0 19320 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_206
timestamp 1676037725
transform 1 0 20056 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1676037725
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_153
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_161
timestamp 1676037725
transform 1 0 15916 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_171
timestamp 1676037725
transform 1 0 16836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_183
timestamp 1676037725
transform 1 0 17940 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_206
timestamp 1676037725
transform 1 0 20056 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_218
timestamp 1676037725
transform 1 0 21160 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_230
timestamp 1676037725
transform 1 0 22264 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1676037725
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_16
timestamp 1676037725
transform 1 0 2576 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_28
timestamp 1676037725
transform 1 0 3680 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_50
timestamp 1676037725
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_65
timestamp 1676037725
transform 1 0 7084 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_83
timestamp 1676037725
transform 1 0 8740 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_91
timestamp 1676037725
transform 1 0 9476 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_121
timestamp 1676037725
transform 1 0 12236 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_140
timestamp 1676037725
transform 1 0 13984 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_146
timestamp 1676037725
transform 1 0 14536 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_151
timestamp 1676037725
transform 1 0 14996 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1676037725
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_174
timestamp 1676037725
transform 1 0 17112 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_186
timestamp 1676037725
transform 1 0 18216 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_195
timestamp 1676037725
transform 1 0 19044 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1676037725
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1676037725
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1676037725
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_33
timestamp 1676037725
transform 1 0 4140 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_50
timestamp 1676037725
transform 1 0 5704 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_58
timestamp 1676037725
transform 1 0 6440 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_110
timestamp 1676037725
transform 1 0 11224 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_159
timestamp 1676037725
transform 1 0 15732 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_164
timestamp 1676037725
transform 1 0 16192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_175
timestamp 1676037725
transform 1 0 17204 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_182
timestamp 1676037725
transform 1 0 17848 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_191
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_204
timestamp 1676037725
transform 1 0 19872 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_216
timestamp 1676037725
transform 1 0 20976 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_228
timestamp 1676037725
transform 1 0 22080 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_232
timestamp 1676037725
transform 1 0 22448 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_11
timestamp 1676037725
transform 1 0 2116 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp 1676037725
transform 1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_31
timestamp 1676037725
transform 1 0 3956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_35
timestamp 1676037725
transform 1 0 4324 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1676037725
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_87
timestamp 1676037725
transform 1 0 9108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_99
timestamp 1676037725
transform 1 0 10212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1676037725
transform 1 0 12236 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_139
timestamp 1676037725
transform 1 0 13892 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_151
timestamp 1676037725
transform 1 0 14996 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_176
timestamp 1676037725
transform 1 0 17296 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_188
timestamp 1676037725
transform 1 0 18400 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_202
timestamp 1676037725
transform 1 0 19688 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_210
timestamp 1676037725
transform 1 0 20424 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_18
timestamp 1676037725
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1676037725
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1676037725
transform 1 0 9476 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_108
timestamp 1676037725
transform 1 0 11040 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_120
timestamp 1676037725
transform 1 0 12144 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_159
timestamp 1676037725
transform 1 0 15732 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_169
timestamp 1676037725
transform 1 0 16652 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_178
timestamp 1676037725
transform 1 0 17480 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp 1676037725
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_203
timestamp 1676037725
transform 1 0 19780 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_215
timestamp 1676037725
transform 1 0 20884 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_227
timestamp 1676037725
transform 1 0 21988 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_11
timestamp 1676037725
transform 1 0 2116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1676037725
transform 1 0 3036 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_28
timestamp 1676037725
transform 1 0 3680 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_40
timestamp 1676037725
transform 1 0 4784 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1676037725
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1676037725
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_144
timestamp 1676037725
transform 1 0 14352 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_156
timestamp 1676037725
transform 1 0 15456 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_178
timestamp 1676037725
transform 1 0 17480 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_186
timestamp 1676037725
transform 1 0 18216 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1676037725
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_11
timestamp 1676037725
transform 1 0 2116 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1676037725
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_61
timestamp 1676037725
transform 1 0 6716 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1676037725
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_93
timestamp 1676037725
transform 1 0 9660 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_110
timestamp 1676037725
transform 1 0 11224 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_118
timestamp 1676037725
transform 1 0 11960 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1676037725
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_156
timestamp 1676037725
transform 1 0 15456 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_168
timestamp 1676037725
transform 1 0 16560 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_172
timestamp 1676037725
transform 1 0 16928 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_181
timestamp 1676037725
transform 1 0 17756 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1676037725
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_206
timestamp 1676037725
transform 1 0 20056 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_218
timestamp 1676037725
transform 1 0 21160 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_230
timestamp 1676037725
transform 1 0 22264 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_17
timestamp 1676037725
transform 1 0 2668 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_24
timestamp 1676037725
transform 1 0 3312 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_36
timestamp 1676037725
transform 1 0 4416 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1676037725
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_65
timestamp 1676037725
transform 1 0 7084 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_84
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_92
timestamp 1676037725
transform 1 0 9568 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1676037725
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_144
timestamp 1676037725
transform 1 0 14352 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_156
timestamp 1676037725
transform 1 0 15456 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_184
timestamp 1676037725
transform 1 0 18032 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_188
timestamp 1676037725
transform 1 0 18400 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_203
timestamp 1676037725
transform 1 0 19780 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_210
timestamp 1676037725
transform 1 0 20424 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1676037725
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1676037725
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_22
timestamp 1676037725
transform 1 0 3128 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1676037725
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_160
timestamp 1676037725
transform 1 0 15824 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_167
timestamp 1676037725
transform 1 0 16468 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_179
timestamp 1676037725
transform 1 0 17572 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_191
timestamp 1676037725
transform 1 0 18676 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1676037725
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_204
timestamp 1676037725
transform 1 0 19872 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_216
timestamp 1676037725
transform 1 0 20976 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_228
timestamp 1676037725
transform 1 0 22080 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_232
timestamp 1676037725
transform 1 0 22448 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_10
timestamp 1676037725
transform 1 0 2024 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_17
timestamp 1676037725
transform 1 0 2668 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_25
timestamp 1676037725
transform 1 0 3404 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_33
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1676037725
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_65
timestamp 1676037725
transform 1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_84
timestamp 1676037725
transform 1 0 8832 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_96
timestamp 1676037725
transform 1 0 9936 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1676037725
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_153
timestamp 1676037725
transform 1 0 15180 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_160
timestamp 1676037725
transform 1 0 15824 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_194
timestamp 1676037725
transform 1 0 18952 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_201
timestamp 1676037725
transform 1 0 19596 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_213
timestamp 1676037725
transform 1 0 20700 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1676037725
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1676037725
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_73
timestamp 1676037725
transform 1 0 7820 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1676037725
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_105
timestamp 1676037725
transform 1 0 10764 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_117
timestamp 1676037725
transform 1 0 11868 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_172
timestamp 1676037725
transform 1 0 16928 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_184
timestamp 1676037725
transform 1 0 18032 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_188
timestamp 1676037725
transform 1 0 18400 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_202
timestamp 1676037725
transform 1 0 19688 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_219
timestamp 1676037725
transform 1 0 21252 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_231
timestamp 1676037725
transform 1 0 22356 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_16
timestamp 1676037725
transform 1 0 2576 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_28
timestamp 1676037725
transform 1 0 3680 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_36
timestamp 1676037725
transform 1 0 4416 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1676037725
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_79
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_107
timestamp 1676037725
transform 1 0 10948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_135
timestamp 1676037725
transform 1 0 13524 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_152
timestamp 1676037725
transform 1 0 15088 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_160
timestamp 1676037725
transform 1 0 15824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_178
timestamp 1676037725
transform 1 0 17480 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_190
timestamp 1676037725
transform 1 0 18584 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_196
timestamp 1676037725
transform 1 0 19136 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1676037725
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1676037725
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1676037725
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1676037725
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_35
timestamp 1676037725
transform 1 0 4324 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_52
timestamp 1676037725
transform 1 0 5888 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_64
timestamp 1676037725
transform 1 0 6992 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_76
timestamp 1676037725
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_117
timestamp 1676037725
transform 1 0 11868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1676037725
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_149
timestamp 1676037725
transform 1 0 14812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_158
timestamp 1676037725
transform 1 0 15640 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_167
timestamp 1676037725
transform 1 0 16468 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_179
timestamp 1676037725
transform 1 0 17572 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1676037725
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1676037725
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1676037725
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1676037725
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_11
timestamp 1676037725
transform 1 0 2116 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_20
timestamp 1676037725
transform 1 0 2944 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_32
timestamp 1676037725
transform 1 0 4048 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_63
timestamp 1676037725
transform 1 0 6900 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_80
timestamp 1676037725
transform 1 0 8464 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_92
timestamp 1676037725
transform 1 0 9568 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1676037725
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_121
timestamp 1676037725
transform 1 0 12236 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_139
timestamp 1676037725
transform 1 0 13892 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_143
timestamp 1676037725
transform 1 0 14260 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_155
timestamp 1676037725
transform 1 0 15364 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1676037725
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_185
timestamp 1676037725
transform 1 0 18124 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_198
timestamp 1676037725
transform 1 0 19320 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_210
timestamp 1676037725
transform 1 0 20424 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_14
timestamp 1676037725
transform 1 0 2392 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_23
timestamp 1676037725
transform 1 0 3220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_51
timestamp 1676037725
transform 1 0 5796 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_63
timestamp 1676037725
transform 1 0 6900 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1676037725
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_92
timestamp 1676037725
transform 1 0 9568 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_117
timestamp 1676037725
transform 1 0 11868 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_159
timestamp 1676037725
transform 1 0 15732 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_169
timestamp 1676037725
transform 1 0 16652 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_177
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1676037725
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_29
timestamp 1676037725
transform 1 0 3772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_41
timestamp 1676037725
transform 1 0 4876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1676037725
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_85
timestamp 1676037725
transform 1 0 8924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_97
timestamp 1676037725
transform 1 0 10028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_109
timestamp 1676037725
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_123
timestamp 1676037725
transform 1 0 12420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_135
timestamp 1676037725
transform 1 0 13524 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_139
timestamp 1676037725
transform 1 0 13892 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_141
timestamp 1676037725
transform 1 0 14076 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_157
timestamp 1676037725
transform 1 0 15548 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1676037725
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_193
timestamp 1676037725
transform 1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_197
timestamp 1676037725
transform 1 0 19228 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_204
timestamp 1676037725
transform 1 0 19872 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_212
timestamp 1676037725
transform 1 0 20608 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 22816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 22816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 22816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 22816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 22816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 22816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 22816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 22816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 22816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 22816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 22816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 22816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 22816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 22816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 22816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 22816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 22816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 22816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 22816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 22816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 22816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 22816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 22816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 22816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 22816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 22816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 22816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 22816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 22816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 22816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 8832 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 13984 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 19136 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16192 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1676037725
transform 1 0 8096 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1676037725
transform -1 0 14076 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1676037725
transform -1 0 7084 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1676037725
transform 1 0 2300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19872 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _188_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_2  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19504 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18676 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16928 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _193_
timestamp 1676037725
transform 1 0 17756 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20792 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19872 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18952 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17664 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _198_
timestamp 1676037725
transform 1 0 17112 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18032 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _200_
timestamp 1676037725
transform 1 0 7268 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _201_
timestamp 1676037725
transform -1 0 2484 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16284 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1676037725
transform -1 0 17112 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _204_
timestamp 1676037725
transform -1 0 4508 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _205_
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20056 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15732 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19044 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _209_
timestamp 1676037725
transform -1 0 11224 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _210_
timestamp 1676037725
transform -1 0 16284 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14352 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _212_
timestamp 1676037725
transform -1 0 11316 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _213_
timestamp 1676037725
transform -1 0 13892 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1676037725
transform 1 0 13800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18400 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _216_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17296 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8004 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4876 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or4b_4  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17940 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__o21ai_1  _220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13800 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10028 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8924 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8004 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9476 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _225_
timestamp 1676037725
transform -1 0 16376 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16192 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15364 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16100 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _229_
timestamp 1676037725
transform -1 0 20056 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_4  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18124 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_4  _231_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18308 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__or4_4  _233_
timestamp 1676037725
transform -1 0 19320 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18492 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19136 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _236_
timestamp 1676037725
transform -1 0 18952 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _237_
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _238_
timestamp 1676037725
transform 1 0 19320 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _240_
timestamp 1676037725
transform -1 0 17480 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_4  _241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18492 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1676037725
transform -1 0 3128 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19320 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _244_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16560 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18124 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _246_
timestamp 1676037725
transform 1 0 20148 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20056 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_2  _248_
timestamp 1676037725
transform 1 0 17020 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__o31a_1  _250_
timestamp 1676037725
transform -1 0 18768 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_4  _251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19780 0 -1 17408
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_1  _252_
timestamp 1676037725
transform 1 0 1748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1676037725
transform 1 0 2392 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _254_
timestamp 1676037725
transform -1 0 3312 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2484 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _257_
timestamp 1676037725
transform 1 0 2116 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _258_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _259_
timestamp 1676037725
transform 1 0 2208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _260_
timestamp 1676037725
transform -1 0 3036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _261_
timestamp 1676037725
transform 1 0 2116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _262_
timestamp 1676037725
transform 1 0 3404 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _263_
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14812 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15272 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _267_
timestamp 1676037725
transform 1 0 16560 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _268_
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _269_
timestamp 1676037725
transform 1 0 16100 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _270_
timestamp 1676037725
transform 1 0 15272 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18032 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _272_
timestamp 1676037725
transform 1 0 18400 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _273_
timestamp 1676037725
transform 1 0 18492 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _274_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _275_
timestamp 1676037725
transform -1 0 17848 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17480 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _277_
timestamp 1676037725
transform 1 0 16560 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _278_
timestamp 1676037725
transform 1 0 15824 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _279_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16836 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _282_
timestamp 1676037725
transform -1 0 14996 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_2  _283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15364 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and4_2  _284_
timestamp 1676037725
transform -1 0 13800 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _286_
timestamp 1676037725
transform 1 0 13064 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _287_
timestamp 1676037725
transform 1 0 10580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _288_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10856 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _289_
timestamp 1676037725
transform -1 0 12512 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _290_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _291_
timestamp 1676037725
transform -1 0 11684 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _292_
timestamp 1676037725
transform -1 0 19688 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _293_
timestamp 1676037725
transform -1 0 16560 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _294_
timestamp 1676037725
transform -1 0 16284 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _295_
timestamp 1676037725
transform -1 0 16284 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _296_
timestamp 1676037725
transform -1 0 18032 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _297_
timestamp 1676037725
transform -1 0 18952 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20148 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _299_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _300_
timestamp 1676037725
transform -1 0 19780 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _301_
timestamp 1676037725
transform 1 0 20056 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _302_
timestamp 1676037725
transform -1 0 15916 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _303_
timestamp 1676037725
transform -1 0 14720 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _304_
timestamp 1676037725
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _305_
timestamp 1676037725
transform -1 0 13616 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _306_
timestamp 1676037725
transform 1 0 12420 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _307_
timestamp 1676037725
transform -1 0 13156 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12512 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _309_
timestamp 1676037725
transform 1 0 11684 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and4_4  _310_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _311_
timestamp 1676037725
transform -1 0 10764 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _312_
timestamp 1676037725
transform -1 0 7728 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _313_
timestamp 1676037725
transform -1 0 6992 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _314_
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _315_
timestamp 1676037725
transform -1 0 6992 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _316_
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _317_
timestamp 1676037725
transform 1 0 6992 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _318_
timestamp 1676037725
transform 1 0 3036 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _319_
timestamp 1676037725
transform 1 0 5060 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _320_
timestamp 1676037725
transform 1 0 3864 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _321_
timestamp 1676037725
transform -1 0 4692 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1676037725
transform 1 0 2944 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _323_
timestamp 1676037725
transform -1 0 4324 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _324_
timestamp 1676037725
transform -1 0 3220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _325_
timestamp 1676037725
transform -1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _326_
timestamp 1676037725
transform -1 0 2116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _327_
timestamp 1676037725
transform 1 0 1932 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _328_
timestamp 1676037725
transform -1 0 2208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _329_
timestamp 1676037725
transform 1 0 2760 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and4_2  _330_
timestamp 1676037725
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _331_
timestamp 1676037725
transform 1 0 3496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _332_
timestamp 1676037725
transform 1 0 5612 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _333_
timestamp 1676037725
transform -1 0 6808 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _334_
timestamp 1676037725
transform -1 0 6992 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _335_
timestamp 1676037725
transform 1 0 5704 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _336_
timestamp 1676037725
transform -1 0 6440 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _337_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7176 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7452 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8372 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _340_
timestamp 1676037725
transform -1 0 9384 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1676037725
transform 1 0 9108 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _342_
timestamp 1676037725
transform -1 0 8556 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _343_
timestamp 1676037725
transform -1 0 15732 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _344_
timestamp 1676037725
transform -1 0 16468 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _345_
timestamp 1676037725
transform -1 0 15088 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _346_
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _347_
timestamp 1676037725
transform 1 0 9108 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _348_
timestamp 1676037725
transform 1 0 1932 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _349_
timestamp 1676037725
transform -1 0 3220 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _350_
timestamp 1676037725
transform -1 0 3496 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _351_
timestamp 1676037725
transform 1 0 3680 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _352_
timestamp 1676037725
transform 1 0 3036 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _353_
timestamp 1676037725
transform -1 0 2116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _354_
timestamp 1676037725
transform -1 0 2484 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _355_
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _356_
timestamp 1676037725
transform -1 0 17388 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _357_
timestamp 1676037725
transform 1 0 16100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _358_
timestamp 1676037725
transform -1 0 15548 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _359_
timestamp 1676037725
transform 1 0 15732 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _360_
timestamp 1676037725
transform 1 0 8004 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _361_
timestamp 1676037725
transform 1 0 2116 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6992 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _363_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _364_
timestamp 1676037725
transform 1 0 12052 0 1 18496
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _365_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12144 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _366_
timestamp 1676037725
transform 1 0 4508 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _367_
timestamp 1676037725
transform -1 0 6072 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _368_
timestamp 1676037725
transform 1 0 7360 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _369_
timestamp 1676037725
transform 1 0 7636 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _370_
timestamp 1676037725
transform 1 0 4416 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _371_
timestamp 1676037725
transform 1 0 9568 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _372_
timestamp 1676037725
transform 1 0 12328 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _373_
timestamp 1676037725
transform 1 0 12512 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _374_
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _375_
timestamp 1676037725
transform 1 0 12328 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _376_
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _377_
timestamp 1676037725
transform 1 0 9476 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _378_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _379_
timestamp 1676037725
transform 1 0 9200 0 1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _380_
timestamp 1676037725
transform 1 0 11316 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _381_
timestamp 1676037725
transform 1 0 12328 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _382_
timestamp 1676037725
transform 1 0 12052 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _383_
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _384_
timestamp 1676037725
transform 1 0 9752 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _385_
timestamp 1676037725
transform 1 0 9752 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _386_
timestamp 1676037725
transform 1 0 7268 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _387_
timestamp 1676037725
transform -1 0 8188 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _388_
timestamp 1676037725
transform 1 0 4232 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _389_
timestamp 1676037725
transform -1 0 5704 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _390_
timestamp 1676037725
transform -1 0 5704 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _391_
timestamp 1676037725
transform 1 0 4232 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _392_
timestamp 1676037725
transform -1 0 5612 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _393_
timestamp 1676037725
transform 1 0 6256 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _394_
timestamp 1676037725
transform 1 0 6348 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _395_
timestamp 1676037725
transform 1 0 8280 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _396_
timestamp 1676037725
transform 1 0 7912 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _397_
timestamp 1676037725
transform -1 0 11868 0 1 20672
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _398_
timestamp 1676037725
transform 1 0 12236 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _399_
timestamp 1676037725
transform 1 0 9292 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1676037725
transform 1 0 12052 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _401_
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _402_
timestamp 1676037725
transform 1 0 6992 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _403_
timestamp 1676037725
transform -1 0 5796 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _404_
timestamp 1676037725
transform -1 0 5796 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _405_
timestamp 1676037725
transform -1 0 5980 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _406_
timestamp 1676037725
transform -1 0 5980 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _407_
timestamp 1676037725
transform -1 0 6072 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _408_
timestamp 1676037725
transform -1 0 5888 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _409_
timestamp 1676037725
transform -1 0 8648 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _410_
timestamp 1676037725
transform 1 0 12420 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _411_
timestamp 1676037725
transform 1 0 9476 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _412_
timestamp 1676037725
transform 1 0 6900 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _413_
timestamp 1676037725
transform 1 0 9752 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _414_
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _415_
timestamp 1676037725
transform 1 0 7360 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9292 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1676037725
transform -1 0 7084 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1676037725
transform -1 0 7084 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1676037725
transform 1 0 10396 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1676037725
transform 1 0 10396 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3036 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout12
timestamp 1676037725
transform 1 0 3404 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout13
timestamp 1676037725
transform -1 0 8924 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 1676037725
transform 1 0 12144 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15824 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout16
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15364 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  fanout18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18400 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19688 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19964 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1676037725
transform -1 0 20608 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1676037725
transform 1 0 12052 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output3
timestamp 1676037725
transform -1 0 2300 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output4
timestamp 1676037725
transform -1 0 5244 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output5
timestamp 1676037725
transform -1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output6
timestamp 1676037725
transform 1 0 10580 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output7
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output8
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output9
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output10
timestamp 1676037725
transform 1 0 20976 0 1 2176
box -38 -48 590 592
<< labels >>
flabel metal2 s 3974 23200 4030 24000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 19982 23200 20038 24000 0 FreeSans 224 90 0 0 io_in
port 1 nsew signal input
flabel metal2 s 1674 0 1730 800 0 FreeSans 224 90 0 0 io_out[0]
port 2 nsew signal tristate
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 io_out[1]
port 3 nsew signal tristate
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 io_out[2]
port 4 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 io_out[3]
port 5 nsew signal tristate
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 io_out[4]
port 6 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 io_out[5]
port 7 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 io_out[6]
port 8 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 io_out[7]
port 9 nsew signal tristate
flabel metal2 s 11978 23200 12034 24000 0 FreeSans 224 90 0 0 rst
port 10 nsew signal input
flabel metal4 s 3658 2128 3978 21808 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 9086 2128 9406 21808 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 14514 2128 14834 21808 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 19942 2128 20262 21808 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 6372 2128 6692 21808 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 11800 2128 12120 21808 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 17228 2128 17548 21808 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 22656 2128 22976 21808 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 24000 24000
<< end >>
