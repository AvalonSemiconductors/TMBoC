magic
tech sky130B
magscale 1 2
timestamp 1683541467
<< nwell >>
rect 1066 37253 38862 37574
rect 1066 36165 38862 36731
rect 1066 35077 38862 35643
rect 1066 33989 38862 34555
rect 1066 32901 38862 33467
rect 1066 31813 38862 32379
rect 1066 30725 38862 31291
rect 1066 29637 38862 30203
rect 1066 28549 38862 29115
rect 1066 27461 38862 28027
rect 1066 26373 38862 26939
rect 1066 25285 38862 25851
rect 1066 24197 38862 24763
rect 1066 23109 38862 23675
rect 1066 22021 38862 22587
rect 1066 20933 38862 21499
rect 1066 19845 38862 20411
rect 1066 18757 38862 19323
rect 1066 17669 38862 18235
rect 1066 16581 38862 17147
rect 1066 15493 38862 16059
rect 1066 14405 38862 14971
rect 1066 13317 38862 13883
rect 1066 12229 38862 12795
rect 1066 11141 38862 11707
rect 1066 10053 38862 10619
rect 1066 8965 38862 9531
rect 1066 7877 38862 8443
rect 1066 6789 38862 7355
rect 1066 5701 38862 6267
rect 1066 4613 38862 5179
rect 1066 3525 38862 4091
rect 1066 2437 38862 3003
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 1104 2128 39086 39160
<< metal2 >>
rect 1766 39200 1822 40000
rect 5078 39200 5134 40000
rect 8390 39200 8446 40000
rect 11702 39200 11758 40000
rect 15014 39200 15070 40000
rect 18326 39200 18382 40000
rect 21638 39200 21694 40000
rect 24950 39200 25006 40000
rect 28262 39200 28318 40000
rect 31574 39200 31630 40000
rect 34886 39200 34942 40000
rect 38198 39200 38254 40000
<< obsm2 >>
rect 1878 39144 5022 39200
rect 5190 39144 8334 39200
rect 8502 39144 11646 39200
rect 11814 39144 14958 39200
rect 15126 39144 18270 39200
rect 18438 39144 21582 39200
rect 21750 39144 24894 39200
rect 25062 39144 28206 39200
rect 28374 39144 31518 39200
rect 31686 39144 34830 39200
rect 34998 39144 38142 39200
rect 38310 39144 39082 39200
rect 1768 1527 39082 39144
<< metal3 >>
rect 39200 38224 40000 38344
rect 39200 36864 40000 36984
rect 39200 35504 40000 35624
rect 39200 34144 40000 34264
rect 39200 32784 40000 32904
rect 39200 31424 40000 31544
rect 39200 30064 40000 30184
rect 39200 28704 40000 28824
rect 39200 27344 40000 27464
rect 39200 25984 40000 26104
rect 39200 24624 40000 24744
rect 39200 23264 40000 23384
rect 39200 21904 40000 22024
rect 39200 20544 40000 20664
rect 39200 19184 40000 19304
rect 39200 17824 40000 17944
rect 39200 16464 40000 16584
rect 39200 15104 40000 15224
rect 39200 13744 40000 13864
rect 39200 12384 40000 12504
rect 39200 11024 40000 11144
rect 39200 9664 40000 9784
rect 39200 8304 40000 8424
rect 39200 6944 40000 7064
rect 39200 5584 40000 5704
rect 39200 4224 40000 4344
rect 39200 2864 40000 2984
rect 39200 1504 40000 1624
<< obsm3 >>
rect 4210 38144 39120 38317
rect 4210 37064 39200 38144
rect 4210 36784 39120 37064
rect 4210 35704 39200 36784
rect 4210 35424 39120 35704
rect 4210 34344 39200 35424
rect 4210 34064 39120 34344
rect 4210 32984 39200 34064
rect 4210 32704 39120 32984
rect 4210 31624 39200 32704
rect 4210 31344 39120 31624
rect 4210 30264 39200 31344
rect 4210 29984 39120 30264
rect 4210 28904 39200 29984
rect 4210 28624 39120 28904
rect 4210 27544 39200 28624
rect 4210 27264 39120 27544
rect 4210 26184 39200 27264
rect 4210 25904 39120 26184
rect 4210 24824 39200 25904
rect 4210 24544 39120 24824
rect 4210 23464 39200 24544
rect 4210 23184 39120 23464
rect 4210 22104 39200 23184
rect 4210 21824 39120 22104
rect 4210 20744 39200 21824
rect 4210 20464 39120 20744
rect 4210 19384 39200 20464
rect 4210 19104 39120 19384
rect 4210 18024 39200 19104
rect 4210 17744 39120 18024
rect 4210 16664 39200 17744
rect 4210 16384 39120 16664
rect 4210 15304 39200 16384
rect 4210 15024 39120 15304
rect 4210 13944 39200 15024
rect 4210 13664 39120 13944
rect 4210 12584 39200 13664
rect 4210 12304 39120 12584
rect 4210 11224 39200 12304
rect 4210 10944 39120 11224
rect 4210 9864 39200 10944
rect 4210 9584 39120 9864
rect 4210 8504 39200 9584
rect 4210 8224 39120 8504
rect 4210 7144 39200 8224
rect 4210 6864 39120 7144
rect 4210 5784 39200 6864
rect 4210 5504 39120 5784
rect 4210 4424 39200 5504
rect 4210 4144 39120 4424
rect 4210 3064 39200 4144
rect 4210 2784 39120 3064
rect 4210 1704 39200 2784
rect 4210 1531 39120 1704
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 5579 3979 19488 36277
rect 19968 3979 34533 36277
<< labels >>
rlabel metal2 s 34886 39200 34942 40000 6 clk
port 1 nsew signal input
rlabel metal2 s 1766 39200 1822 40000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 5078 39200 5134 40000 6 io_in[1]
port 3 nsew signal input
rlabel metal2 s 8390 39200 8446 40000 6 io_in[2]
port 4 nsew signal input
rlabel metal2 s 11702 39200 11758 40000 6 io_in[3]
port 5 nsew signal input
rlabel metal2 s 15014 39200 15070 40000 6 io_in[4]
port 6 nsew signal input
rlabel metal2 s 18326 39200 18382 40000 6 io_in[5]
port 7 nsew signal input
rlabel metal2 s 21638 39200 21694 40000 6 io_in[6]
port 8 nsew signal input
rlabel metal2 s 24950 39200 25006 40000 6 io_in[7]
port 9 nsew signal input
rlabel metal2 s 28262 39200 28318 40000 6 io_in[8]
port 10 nsew signal input
rlabel metal2 s 31574 39200 31630 40000 6 io_in[9]
port 11 nsew signal input
rlabel metal3 s 39200 38224 40000 38344 6 io_oeb
port 12 nsew signal output
rlabel metal3 s 39200 1504 40000 1624 6 io_out[0]
port 13 nsew signal output
rlabel metal3 s 39200 15104 40000 15224 6 io_out[10]
port 14 nsew signal output
rlabel metal3 s 39200 16464 40000 16584 6 io_out[11]
port 15 nsew signal output
rlabel metal3 s 39200 17824 40000 17944 6 io_out[12]
port 16 nsew signal output
rlabel metal3 s 39200 19184 40000 19304 6 io_out[13]
port 17 nsew signal output
rlabel metal3 s 39200 20544 40000 20664 6 io_out[14]
port 18 nsew signal output
rlabel metal3 s 39200 21904 40000 22024 6 io_out[15]
port 19 nsew signal output
rlabel metal3 s 39200 23264 40000 23384 6 io_out[16]
port 20 nsew signal output
rlabel metal3 s 39200 24624 40000 24744 6 io_out[17]
port 21 nsew signal output
rlabel metal3 s 39200 25984 40000 26104 6 io_out[18]
port 22 nsew signal output
rlabel metal3 s 39200 27344 40000 27464 6 io_out[19]
port 23 nsew signal output
rlabel metal3 s 39200 2864 40000 2984 6 io_out[1]
port 24 nsew signal output
rlabel metal3 s 39200 28704 40000 28824 6 io_out[20]
port 25 nsew signal output
rlabel metal3 s 39200 30064 40000 30184 6 io_out[21]
port 26 nsew signal output
rlabel metal3 s 39200 31424 40000 31544 6 io_out[22]
port 27 nsew signal output
rlabel metal3 s 39200 32784 40000 32904 6 io_out[23]
port 28 nsew signal output
rlabel metal3 s 39200 34144 40000 34264 6 io_out[24]
port 29 nsew signal output
rlabel metal3 s 39200 35504 40000 35624 6 io_out[25]
port 30 nsew signal output
rlabel metal3 s 39200 36864 40000 36984 6 io_out[26]
port 31 nsew signal output
rlabel metal3 s 39200 4224 40000 4344 6 io_out[2]
port 32 nsew signal output
rlabel metal3 s 39200 5584 40000 5704 6 io_out[3]
port 33 nsew signal output
rlabel metal3 s 39200 6944 40000 7064 6 io_out[4]
port 34 nsew signal output
rlabel metal3 s 39200 8304 40000 8424 6 io_out[5]
port 35 nsew signal output
rlabel metal3 s 39200 9664 40000 9784 6 io_out[6]
port 36 nsew signal output
rlabel metal3 s 39200 11024 40000 11144 6 io_out[7]
port 37 nsew signal output
rlabel metal3 s 39200 12384 40000 12504 6 io_out[8]
port 38 nsew signal output
rlabel metal3 s 39200 13744 40000 13864 6 io_out[9]
port 39 nsew signal output
rlabel metal2 s 38198 39200 38254 40000 6 rst
port 40 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 42 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4112314
string GDS_FILE /media/lucah/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/MOS6502/runs/23_05_08_12_20/results/signoff/wrapped_6502.magic.gds
string GDS_START 1064460
<< end >>

