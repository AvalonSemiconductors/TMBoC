VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiplexer
  CLASS BLOCK ;
  FOREIGN multiplexer ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN design_clk_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END design_clk_o
  PIN dsi_all[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END dsi_all[0]
  PIN dsi_all[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END dsi_all[10]
  PIN dsi_all[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END dsi_all[11]
  PIN dsi_all[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END dsi_all[12]
  PIN dsi_all[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END dsi_all[13]
  PIN dsi_all[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END dsi_all[14]
  PIN dsi_all[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END dsi_all[15]
  PIN dsi_all[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END dsi_all[16]
  PIN dsi_all[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END dsi_all[17]
  PIN dsi_all[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END dsi_all[18]
  PIN dsi_all[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END dsi_all[19]
  PIN dsi_all[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END dsi_all[1]
  PIN dsi_all[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END dsi_all[20]
  PIN dsi_all[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END dsi_all[21]
  PIN dsi_all[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END dsi_all[22]
  PIN dsi_all[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END dsi_all[23]
  PIN dsi_all[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END dsi_all[24]
  PIN dsi_all[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END dsi_all[25]
  PIN dsi_all[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END dsi_all[26]
  PIN dsi_all[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END dsi_all[27]
  PIN dsi_all[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END dsi_all[2]
  PIN dsi_all[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END dsi_all[3]
  PIN dsi_all[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END dsi_all[4]
  PIN dsi_all[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END dsi_all[5]
  PIN dsi_all[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END dsi_all[6]
  PIN dsi_all[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END dsi_all[7]
  PIN dsi_all[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END dsi_all[8]
  PIN dsi_all[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END dsi_all[9]
  PIN dso_6502[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END dso_6502[0]
  PIN dso_6502[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END dso_6502[10]
  PIN dso_6502[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END dso_6502[11]
  PIN dso_6502[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END dso_6502[12]
  PIN dso_6502[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END dso_6502[13]
  PIN dso_6502[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END dso_6502[14]
  PIN dso_6502[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END dso_6502[15]
  PIN dso_6502[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END dso_6502[16]
  PIN dso_6502[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END dso_6502[17]
  PIN dso_6502[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END dso_6502[18]
  PIN dso_6502[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END dso_6502[19]
  PIN dso_6502[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END dso_6502[1]
  PIN dso_6502[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END dso_6502[20]
  PIN dso_6502[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END dso_6502[21]
  PIN dso_6502[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END dso_6502[22]
  PIN dso_6502[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END dso_6502[23]
  PIN dso_6502[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 0.000 227.150 4.000 ;
    END
  END dso_6502[24]
  PIN dso_6502[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END dso_6502[25]
  PIN dso_6502[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END dso_6502[26]
  PIN dso_6502[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END dso_6502[2]
  PIN dso_6502[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END dso_6502[3]
  PIN dso_6502[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END dso_6502[4]
  PIN dso_6502[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END dso_6502[5]
  PIN dso_6502[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END dso_6502[6]
  PIN dso_6502[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END dso_6502[7]
  PIN dso_6502[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END dso_6502[8]
  PIN dso_6502[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END dso_6502[9]
  PIN dso_LCD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END dso_LCD[0]
  PIN dso_LCD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END dso_LCD[1]
  PIN dso_LCD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END dso_LCD[2]
  PIN dso_LCD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END dso_LCD[3]
  PIN dso_LCD[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END dso_LCD[4]
  PIN dso_LCD[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END dso_LCD[5]
  PIN dso_LCD[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END dso_LCD[6]
  PIN dso_LCD[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END dso_LCD[7]
  PIN dso_as1802[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END dso_as1802[0]
  PIN dso_as1802[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END dso_as1802[10]
  PIN dso_as1802[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END dso_as1802[11]
  PIN dso_as1802[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END dso_as1802[12]
  PIN dso_as1802[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END dso_as1802[13]
  PIN dso_as1802[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END dso_as1802[14]
  PIN dso_as1802[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END dso_as1802[15]
  PIN dso_as1802[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END dso_as1802[16]
  PIN dso_as1802[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END dso_as1802[17]
  PIN dso_as1802[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END dso_as1802[18]
  PIN dso_as1802[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END dso_as1802[19]
  PIN dso_as1802[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END dso_as1802[1]
  PIN dso_as1802[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END dso_as1802[20]
  PIN dso_as1802[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END dso_as1802[21]
  PIN dso_as1802[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END dso_as1802[22]
  PIN dso_as1802[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END dso_as1802[23]
  PIN dso_as1802[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END dso_as1802[24]
  PIN dso_as1802[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END dso_as1802[25]
  PIN dso_as1802[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END dso_as1802[26]
  PIN dso_as1802[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END dso_as1802[2]
  PIN dso_as1802[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END dso_as1802[3]
  PIN dso_as1802[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END dso_as1802[4]
  PIN dso_as1802[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END dso_as1802[5]
  PIN dso_as1802[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END dso_as1802[6]
  PIN dso_as1802[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END dso_as1802[7]
  PIN dso_as1802[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END dso_as1802[8]
  PIN dso_as1802[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END dso_as1802[9]
  PIN dso_as2650[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 296.000 120.890 300.000 ;
    END
  END dso_as2650[0]
  PIN dso_as2650[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 296.000 185.290 300.000 ;
    END
  END dso_as2650[10]
  PIN dso_as2650[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 296.000 191.730 300.000 ;
    END
  END dso_as2650[11]
  PIN dso_as2650[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 296.000 198.170 300.000 ;
    END
  END dso_as2650[12]
  PIN dso_as2650[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 296.000 204.610 300.000 ;
    END
  END dso_as2650[13]
  PIN dso_as2650[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 296.000 211.050 300.000 ;
    END
  END dso_as2650[14]
  PIN dso_as2650[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 296.000 217.490 300.000 ;
    END
  END dso_as2650[15]
  PIN dso_as2650[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 296.000 223.930 300.000 ;
    END
  END dso_as2650[16]
  PIN dso_as2650[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 296.000 230.370 300.000 ;
    END
  END dso_as2650[17]
  PIN dso_as2650[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 296.000 236.810 300.000 ;
    END
  END dso_as2650[18]
  PIN dso_as2650[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 296.000 243.250 300.000 ;
    END
  END dso_as2650[19]
  PIN dso_as2650[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 296.000 127.330 300.000 ;
    END
  END dso_as2650[1]
  PIN dso_as2650[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 296.000 249.690 300.000 ;
    END
  END dso_as2650[20]
  PIN dso_as2650[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 296.000 256.130 300.000 ;
    END
  END dso_as2650[21]
  PIN dso_as2650[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 296.000 262.570 300.000 ;
    END
  END dso_as2650[22]
  PIN dso_as2650[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 296.000 269.010 300.000 ;
    END
  END dso_as2650[23]
  PIN dso_as2650[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 296.000 275.450 300.000 ;
    END
  END dso_as2650[24]
  PIN dso_as2650[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 296.000 281.890 300.000 ;
    END
  END dso_as2650[25]
  PIN dso_as2650[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 296.000 288.330 300.000 ;
    END
  END dso_as2650[26]
  PIN dso_as2650[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 296.000 133.770 300.000 ;
    END
  END dso_as2650[2]
  PIN dso_as2650[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 296.000 140.210 300.000 ;
    END
  END dso_as2650[3]
  PIN dso_as2650[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 296.000 146.650 300.000 ;
    END
  END dso_as2650[4]
  PIN dso_as2650[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 296.000 153.090 300.000 ;
    END
  END dso_as2650[5]
  PIN dso_as2650[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 296.000 159.530 300.000 ;
    END
  END dso_as2650[6]
  PIN dso_as2650[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 296.000 165.970 300.000 ;
    END
  END dso_as2650[7]
  PIN dso_as2650[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 296.000 172.410 300.000 ;
    END
  END dso_as2650[8]
  PIN dso_as2650[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 296.000 178.850 300.000 ;
    END
  END dso_as2650[9]
  PIN dso_as512512512[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END dso_as512512512[0]
  PIN dso_as512512512[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END dso_as512512512[10]
  PIN dso_as512512512[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END dso_as512512512[11]
  PIN dso_as512512512[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END dso_as512512512[12]
  PIN dso_as512512512[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END dso_as512512512[13]
  PIN dso_as512512512[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END dso_as512512512[14]
  PIN dso_as512512512[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END dso_as512512512[15]
  PIN dso_as512512512[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END dso_as512512512[16]
  PIN dso_as512512512[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END dso_as512512512[17]
  PIN dso_as512512512[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END dso_as512512512[18]
  PIN dso_as512512512[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END dso_as512512512[19]
  PIN dso_as512512512[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END dso_as512512512[1]
  PIN dso_as512512512[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END dso_as512512512[20]
  PIN dso_as512512512[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END dso_as512512512[21]
  PIN dso_as512512512[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END dso_as512512512[22]
  PIN dso_as512512512[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END dso_as512512512[23]
  PIN dso_as512512512[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END dso_as512512512[24]
  PIN dso_as512512512[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END dso_as512512512[25]
  PIN dso_as512512512[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END dso_as512512512[26]
  PIN dso_as512512512[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END dso_as512512512[27]
  PIN dso_as512512512[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END dso_as512512512[2]
  PIN dso_as512512512[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END dso_as512512512[3]
  PIN dso_as512512512[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END dso_as512512512[4]
  PIN dso_as512512512[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END dso_as512512512[5]
  PIN dso_as512512512[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END dso_as512512512[6]
  PIN dso_as512512512[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END dso_as512512512[7]
  PIN dso_as512512512[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END dso_as512512512[8]
  PIN dso_as512512512[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END dso_as512512512[9]
  PIN dso_as5401[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 238.040 300.000 238.640 ;
    END
  END dso_as5401[0]
  PIN dso_as5401[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.440 300.000 259.040 ;
    END
  END dso_as5401[10]
  PIN dso_as5401[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 260.480 300.000 261.080 ;
    END
  END dso_as5401[11]
  PIN dso_as5401[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 262.520 300.000 263.120 ;
    END
  END dso_as5401[12]
  PIN dso_as5401[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 264.560 300.000 265.160 ;
    END
  END dso_as5401[13]
  PIN dso_as5401[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 266.600 300.000 267.200 ;
    END
  END dso_as5401[14]
  PIN dso_as5401[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 268.640 300.000 269.240 ;
    END
  END dso_as5401[15]
  PIN dso_as5401[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 270.680 300.000 271.280 ;
    END
  END dso_as5401[16]
  PIN dso_as5401[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 272.720 300.000 273.320 ;
    END
  END dso_as5401[17]
  PIN dso_as5401[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 274.760 300.000 275.360 ;
    END
  END dso_as5401[18]
  PIN dso_as5401[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 276.800 300.000 277.400 ;
    END
  END dso_as5401[19]
  PIN dso_as5401[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 240.080 300.000 240.680 ;
    END
  END dso_as5401[1]
  PIN dso_as5401[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 278.840 300.000 279.440 ;
    END
  END dso_as5401[20]
  PIN dso_as5401[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 280.880 300.000 281.480 ;
    END
  END dso_as5401[21]
  PIN dso_as5401[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 282.920 300.000 283.520 ;
    END
  END dso_as5401[22]
  PIN dso_as5401[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 284.960 300.000 285.560 ;
    END
  END dso_as5401[23]
  PIN dso_as5401[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 287.000 300.000 287.600 ;
    END
  END dso_as5401[24]
  PIN dso_as5401[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 289.040 300.000 289.640 ;
    END
  END dso_as5401[25]
  PIN dso_as5401[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 291.080 300.000 291.680 ;
    END
  END dso_as5401[26]
  PIN dso_as5401[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 242.120 300.000 242.720 ;
    END
  END dso_as5401[2]
  PIN dso_as5401[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 244.160 300.000 244.760 ;
    END
  END dso_as5401[3]
  PIN dso_as5401[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 246.200 300.000 246.800 ;
    END
  END dso_as5401[4]
  PIN dso_as5401[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 248.240 300.000 248.840 ;
    END
  END dso_as5401[5]
  PIN dso_as5401[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 250.280 300.000 250.880 ;
    END
  END dso_as5401[6]
  PIN dso_as5401[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 252.320 300.000 252.920 ;
    END
  END dso_as5401[7]
  PIN dso_as5401[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 254.360 300.000 254.960 ;
    END
  END dso_as5401[8]
  PIN dso_as5401[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 256.400 300.000 257.000 ;
    END
  END dso_as5401[9]
  PIN dso_counter[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 213.560 300.000 214.160 ;
    END
  END dso_counter[0]
  PIN dso_counter[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 233.960 300.000 234.560 ;
    END
  END dso_counter[10]
  PIN dso_counter[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 236.000 300.000 236.600 ;
    END
  END dso_counter[11]
  PIN dso_counter[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 215.600 300.000 216.200 ;
    END
  END dso_counter[1]
  PIN dso_counter[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 217.640 300.000 218.240 ;
    END
  END dso_counter[2]
  PIN dso_counter[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 219.680 300.000 220.280 ;
    END
  END dso_counter[3]
  PIN dso_counter[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 221.720 300.000 222.320 ;
    END
  END dso_counter[4]
  PIN dso_counter[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 223.760 300.000 224.360 ;
    END
  END dso_counter[5]
  PIN dso_counter[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 225.800 300.000 226.400 ;
    END
  END dso_counter[6]
  PIN dso_counter[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 227.840 300.000 228.440 ;
    END
  END dso_counter[7]
  PIN dso_counter[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 229.880 300.000 230.480 ;
    END
  END dso_counter[8]
  PIN dso_counter[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 231.920 300.000 232.520 ;
    END
  END dso_counter[9]
  PIN dso_diceroll[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 296.000 62.930 300.000 ;
    END
  END dso_diceroll[0]
  PIN dso_diceroll[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 296.000 69.370 300.000 ;
    END
  END dso_diceroll[1]
  PIN dso_diceroll[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 296.000 75.810 300.000 ;
    END
  END dso_diceroll[2]
  PIN dso_diceroll[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 296.000 82.250 300.000 ;
    END
  END dso_diceroll[3]
  PIN dso_diceroll[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 296.000 88.690 300.000 ;
    END
  END dso_diceroll[4]
  PIN dso_diceroll[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 296.000 95.130 300.000 ;
    END
  END dso_diceroll[5]
  PIN dso_diceroll[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 296.000 101.570 300.000 ;
    END
  END dso_diceroll[6]
  PIN dso_diceroll[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 296.000 108.010 300.000 ;
    END
  END dso_diceroll[7]
  PIN dso_mc14500[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END dso_mc14500[0]
  PIN dso_mc14500[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END dso_mc14500[1]
  PIN dso_mc14500[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END dso_mc14500[2]
  PIN dso_mc14500[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END dso_mc14500[3]
  PIN dso_mc14500[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END dso_mc14500[4]
  PIN dso_mc14500[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END dso_mc14500[5]
  PIN dso_mc14500[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END dso_mc14500[6]
  PIN dso_mc14500[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END dso_mc14500[7]
  PIN dso_mc14500[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END dso_mc14500[8]
  PIN dso_multiplier[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 296.000 11.410 300.000 ;
    END
  END dso_multiplier[0]
  PIN dso_multiplier[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 296.000 17.850 300.000 ;
    END
  END dso_multiplier[1]
  PIN dso_multiplier[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 296.000 24.290 300.000 ;
    END
  END dso_multiplier[2]
  PIN dso_multiplier[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 296.000 30.730 300.000 ;
    END
  END dso_multiplier[3]
  PIN dso_multiplier[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 296.000 37.170 300.000 ;
    END
  END dso_multiplier[4]
  PIN dso_multiplier[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 296.000 43.610 300.000 ;
    END
  END dso_multiplier[5]
  PIN dso_multiplier[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 296.000 50.050 300.000 ;
    END
  END dso_multiplier[6]
  PIN dso_multiplier[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 296.000 56.490 300.000 ;
    END
  END dso_multiplier[7]
  PIN dso_posit[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END dso_posit[0]
  PIN dso_posit[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END dso_posit[1]
  PIN dso_posit[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END dso_posit[2]
  PIN dso_posit[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END dso_posit[3]
  PIN dso_tbb1143[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END dso_tbb1143[0]
  PIN dso_tbb1143[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END dso_tbb1143[1]
  PIN dso_tbb1143[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END dso_tbb1143[2]
  PIN dso_tbb1143[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END dso_tbb1143[3]
  PIN dso_tbb1143[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END dso_tbb1143[4]
  PIN dso_tbb1143[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END dso_tbb1143[5]
  PIN dso_tbb1143[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END dso_tbb1143[6]
  PIN dso_tbb1143[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END dso_tbb1143[7]
  PIN dso_tune
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END dso_tune
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END io_out[9]
  PIN oeb_6502
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END oeb_6502
  PIN oeb_as1802
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END oeb_as1802
  PIN oeb_as2650
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 296.000 114.450 300.000 ;
    END
  END oeb_as2650
  PIN oeb_as512512512
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END oeb_as512512512
  PIN oeb_as5401
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 293.120 300.000 293.720 ;
    END
  END oeb_as5401
  PIN oeb_mc14500
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END oeb_mc14500
  PIN rst_6502
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END rst_6502
  PIN rst_LCD
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END rst_LCD
  PIN rst_as1802
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END rst_as1802
  PIN rst_as2650
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END rst_as2650
  PIN rst_as512512512
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END rst_as512512512
  PIN rst_as5401
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END rst_as5401
  PIN rst_counter
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END rst_counter
  PIN rst_diceroll
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END rst_diceroll
  PIN rst_mc14500
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END rst_mc14500
  PIN rst_posit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END rst_posit
  PIN rst_tbb1143
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END rst_tbb1143
  PIN rst_tune
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END rst_tune
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 5.480 300.000 6.080 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 7.520 300.000 8.120 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 9.560 300.000 10.160 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 17.720 300.000 18.320 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 78.920 300.000 79.520 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 85.040 300.000 85.640 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 91.160 300.000 91.760 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 97.280 300.000 97.880 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 103.400 300.000 104.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 109.520 300.000 110.120 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 115.640 300.000 116.240 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 121.760 300.000 122.360 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 127.880 300.000 128.480 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 134.000 300.000 134.600 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 23.840 300.000 24.440 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 140.120 300.000 140.720 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 146.240 300.000 146.840 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 152.360 300.000 152.960 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 158.480 300.000 159.080 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 164.600 300.000 165.200 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 170.720 300.000 171.320 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 176.840 300.000 177.440 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 182.960 300.000 183.560 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 189.080 300.000 189.680 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 195.200 300.000 195.800 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 29.960 300.000 30.560 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.320 300.000 201.920 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 207.440 300.000 208.040 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 36.080 300.000 36.680 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 42.200 300.000 42.800 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 48.320 300.000 48.920 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 54.440 300.000 55.040 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 60.560 300.000 61.160 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 66.680 300.000 67.280 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 72.800 300.000 73.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 11.600 300.000 12.200 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 19.760 300.000 20.360 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 80.960 300.000 81.560 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 87.080 300.000 87.680 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 93.200 300.000 93.800 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 99.320 300.000 99.920 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 105.440 300.000 106.040 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 111.560 300.000 112.160 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 117.680 300.000 118.280 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 123.800 300.000 124.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 129.920 300.000 130.520 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 136.040 300.000 136.640 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 25.880 300.000 26.480 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 142.160 300.000 142.760 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 148.280 300.000 148.880 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 154.400 300.000 155.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 160.520 300.000 161.120 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 166.640 300.000 167.240 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 172.760 300.000 173.360 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 178.880 300.000 179.480 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 185.000 300.000 185.600 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 191.120 300.000 191.720 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 197.240 300.000 197.840 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 32.000 300.000 32.600 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 203.360 300.000 203.960 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 209.480 300.000 210.080 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 38.120 300.000 38.720 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 44.240 300.000 44.840 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 50.360 300.000 50.960 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 56.480 300.000 57.080 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 62.600 300.000 63.200 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 68.720 300.000 69.320 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 74.840 300.000 75.440 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 21.800 300.000 22.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 83.000 300.000 83.600 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 89.120 300.000 89.720 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 95.240 300.000 95.840 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 101.360 300.000 101.960 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 107.480 300.000 108.080 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 113.600 300.000 114.200 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 119.720 300.000 120.320 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 125.840 300.000 126.440 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 131.960 300.000 132.560 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 138.080 300.000 138.680 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 27.920 300.000 28.520 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 144.200 300.000 144.800 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 150.320 300.000 150.920 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 156.440 300.000 157.040 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 162.560 300.000 163.160 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 168.680 300.000 169.280 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 174.800 300.000 175.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 180.920 300.000 181.520 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 187.040 300.000 187.640 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 193.160 300.000 193.760 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 199.280 300.000 199.880 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 34.040 300.000 34.640 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 205.400 300.000 206.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 211.520 300.000 212.120 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 40.160 300.000 40.760 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 46.280 300.000 46.880 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 52.400 300.000 53.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 58.520 300.000 59.120 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 64.640 300.000 65.240 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 70.760 300.000 71.360 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 76.880 300.000 77.480 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 13.640 300.000 14.240 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 15.680 300.000 16.280 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 288.405 ;
      LAYER met1 ;
        RECT 4.670 0.380 298.930 295.760 ;
      LAYER met2 ;
        RECT 4.690 295.720 10.850 296.000 ;
        RECT 11.690 295.720 17.290 296.000 ;
        RECT 18.130 295.720 23.730 296.000 ;
        RECT 24.570 295.720 30.170 296.000 ;
        RECT 31.010 295.720 36.610 296.000 ;
        RECT 37.450 295.720 43.050 296.000 ;
        RECT 43.890 295.720 49.490 296.000 ;
        RECT 50.330 295.720 55.930 296.000 ;
        RECT 56.770 295.720 62.370 296.000 ;
        RECT 63.210 295.720 68.810 296.000 ;
        RECT 69.650 295.720 75.250 296.000 ;
        RECT 76.090 295.720 81.690 296.000 ;
        RECT 82.530 295.720 88.130 296.000 ;
        RECT 88.970 295.720 94.570 296.000 ;
        RECT 95.410 295.720 101.010 296.000 ;
        RECT 101.850 295.720 107.450 296.000 ;
        RECT 108.290 295.720 113.890 296.000 ;
        RECT 114.730 295.720 120.330 296.000 ;
        RECT 121.170 295.720 126.770 296.000 ;
        RECT 127.610 295.720 133.210 296.000 ;
        RECT 134.050 295.720 139.650 296.000 ;
        RECT 140.490 295.720 146.090 296.000 ;
        RECT 146.930 295.720 152.530 296.000 ;
        RECT 153.370 295.720 158.970 296.000 ;
        RECT 159.810 295.720 165.410 296.000 ;
        RECT 166.250 295.720 171.850 296.000 ;
        RECT 172.690 295.720 178.290 296.000 ;
        RECT 179.130 295.720 184.730 296.000 ;
        RECT 185.570 295.720 191.170 296.000 ;
        RECT 192.010 295.720 197.610 296.000 ;
        RECT 198.450 295.720 204.050 296.000 ;
        RECT 204.890 295.720 210.490 296.000 ;
        RECT 211.330 295.720 216.930 296.000 ;
        RECT 217.770 295.720 223.370 296.000 ;
        RECT 224.210 295.720 229.810 296.000 ;
        RECT 230.650 295.720 236.250 296.000 ;
        RECT 237.090 295.720 242.690 296.000 ;
        RECT 243.530 295.720 249.130 296.000 ;
        RECT 249.970 295.720 255.570 296.000 ;
        RECT 256.410 295.720 262.010 296.000 ;
        RECT 262.850 295.720 268.450 296.000 ;
        RECT 269.290 295.720 274.890 296.000 ;
        RECT 275.730 295.720 281.330 296.000 ;
        RECT 282.170 295.720 287.770 296.000 ;
        RECT 288.610 295.720 298.900 296.000 ;
        RECT 4.690 4.280 298.900 295.720 ;
        RECT 4.690 0.350 29.250 4.280 ;
        RECT 30.090 0.350 30.630 4.280 ;
        RECT 31.470 0.350 32.010 4.280 ;
        RECT 32.850 0.350 33.390 4.280 ;
        RECT 34.230 0.350 34.770 4.280 ;
        RECT 35.610 0.350 36.150 4.280 ;
        RECT 36.990 0.350 37.530 4.280 ;
        RECT 38.370 0.350 38.910 4.280 ;
        RECT 39.750 0.350 40.290 4.280 ;
        RECT 41.130 0.350 41.670 4.280 ;
        RECT 42.510 0.350 43.050 4.280 ;
        RECT 43.890 0.350 44.430 4.280 ;
        RECT 45.270 0.350 45.810 4.280 ;
        RECT 46.650 0.350 47.190 4.280 ;
        RECT 48.030 0.350 48.570 4.280 ;
        RECT 49.410 0.350 49.950 4.280 ;
        RECT 50.790 0.350 51.330 4.280 ;
        RECT 52.170 0.350 52.710 4.280 ;
        RECT 53.550 0.350 54.090 4.280 ;
        RECT 54.930 0.350 55.470 4.280 ;
        RECT 56.310 0.350 56.850 4.280 ;
        RECT 57.690 0.350 58.230 4.280 ;
        RECT 59.070 0.350 59.610 4.280 ;
        RECT 60.450 0.350 60.990 4.280 ;
        RECT 61.830 0.350 62.370 4.280 ;
        RECT 63.210 0.350 63.750 4.280 ;
        RECT 64.590 0.350 65.130 4.280 ;
        RECT 65.970 0.350 66.510 4.280 ;
        RECT 67.350 0.350 67.890 4.280 ;
        RECT 68.730 0.350 69.270 4.280 ;
        RECT 70.110 0.350 70.650 4.280 ;
        RECT 71.490 0.350 72.030 4.280 ;
        RECT 72.870 0.350 73.410 4.280 ;
        RECT 74.250 0.350 74.790 4.280 ;
        RECT 75.630 0.350 76.170 4.280 ;
        RECT 77.010 0.350 77.550 4.280 ;
        RECT 78.390 0.350 78.930 4.280 ;
        RECT 79.770 0.350 80.310 4.280 ;
        RECT 81.150 0.350 81.690 4.280 ;
        RECT 82.530 0.350 83.070 4.280 ;
        RECT 83.910 0.350 84.450 4.280 ;
        RECT 85.290 0.350 85.830 4.280 ;
        RECT 86.670 0.350 87.210 4.280 ;
        RECT 88.050 0.350 88.590 4.280 ;
        RECT 89.430 0.350 89.970 4.280 ;
        RECT 90.810 0.350 91.350 4.280 ;
        RECT 92.190 0.350 92.730 4.280 ;
        RECT 93.570 0.350 94.110 4.280 ;
        RECT 94.950 0.350 95.490 4.280 ;
        RECT 96.330 0.350 96.870 4.280 ;
        RECT 97.710 0.350 98.250 4.280 ;
        RECT 99.090 0.350 99.630 4.280 ;
        RECT 100.470 0.350 101.010 4.280 ;
        RECT 101.850 0.350 102.390 4.280 ;
        RECT 103.230 0.350 103.770 4.280 ;
        RECT 104.610 0.350 105.150 4.280 ;
        RECT 105.990 0.350 106.530 4.280 ;
        RECT 107.370 0.350 107.910 4.280 ;
        RECT 108.750 0.350 109.290 4.280 ;
        RECT 110.130 0.350 110.670 4.280 ;
        RECT 111.510 0.350 112.050 4.280 ;
        RECT 112.890 0.350 113.430 4.280 ;
        RECT 114.270 0.350 114.810 4.280 ;
        RECT 115.650 0.350 116.190 4.280 ;
        RECT 117.030 0.350 117.570 4.280 ;
        RECT 118.410 0.350 118.950 4.280 ;
        RECT 119.790 0.350 120.330 4.280 ;
        RECT 121.170 0.350 121.710 4.280 ;
        RECT 122.550 0.350 123.090 4.280 ;
        RECT 123.930 0.350 124.470 4.280 ;
        RECT 125.310 0.350 125.850 4.280 ;
        RECT 126.690 0.350 127.230 4.280 ;
        RECT 128.070 0.350 128.610 4.280 ;
        RECT 129.450 0.350 129.990 4.280 ;
        RECT 130.830 0.350 131.370 4.280 ;
        RECT 132.210 0.350 132.750 4.280 ;
        RECT 133.590 0.350 134.130 4.280 ;
        RECT 134.970 0.350 135.510 4.280 ;
        RECT 136.350 0.350 136.890 4.280 ;
        RECT 137.730 0.350 138.270 4.280 ;
        RECT 139.110 0.350 139.650 4.280 ;
        RECT 140.490 0.350 141.030 4.280 ;
        RECT 141.870 0.350 142.410 4.280 ;
        RECT 143.250 0.350 143.790 4.280 ;
        RECT 144.630 0.350 145.170 4.280 ;
        RECT 146.010 0.350 146.550 4.280 ;
        RECT 147.390 0.350 147.930 4.280 ;
        RECT 148.770 0.350 149.310 4.280 ;
        RECT 150.150 0.350 150.690 4.280 ;
        RECT 151.530 0.350 152.070 4.280 ;
        RECT 152.910 0.350 153.450 4.280 ;
        RECT 154.290 0.350 154.830 4.280 ;
        RECT 155.670 0.350 156.210 4.280 ;
        RECT 157.050 0.350 157.590 4.280 ;
        RECT 158.430 0.350 158.970 4.280 ;
        RECT 159.810 0.350 160.350 4.280 ;
        RECT 161.190 0.350 161.730 4.280 ;
        RECT 162.570 0.350 163.110 4.280 ;
        RECT 163.950 0.350 164.490 4.280 ;
        RECT 165.330 0.350 165.870 4.280 ;
        RECT 166.710 0.350 167.250 4.280 ;
        RECT 168.090 0.350 168.630 4.280 ;
        RECT 169.470 0.350 170.010 4.280 ;
        RECT 170.850 0.350 171.390 4.280 ;
        RECT 172.230 0.350 172.770 4.280 ;
        RECT 173.610 0.350 174.150 4.280 ;
        RECT 174.990 0.350 175.530 4.280 ;
        RECT 176.370 0.350 176.910 4.280 ;
        RECT 177.750 0.350 178.290 4.280 ;
        RECT 179.130 0.350 179.670 4.280 ;
        RECT 180.510 0.350 181.050 4.280 ;
        RECT 181.890 0.350 182.430 4.280 ;
        RECT 183.270 0.350 183.810 4.280 ;
        RECT 184.650 0.350 185.190 4.280 ;
        RECT 186.030 0.350 186.570 4.280 ;
        RECT 187.410 0.350 187.950 4.280 ;
        RECT 188.790 0.350 189.330 4.280 ;
        RECT 190.170 0.350 190.710 4.280 ;
        RECT 191.550 0.350 192.090 4.280 ;
        RECT 192.930 0.350 193.470 4.280 ;
        RECT 194.310 0.350 194.850 4.280 ;
        RECT 195.690 0.350 196.230 4.280 ;
        RECT 197.070 0.350 197.610 4.280 ;
        RECT 198.450 0.350 198.990 4.280 ;
        RECT 199.830 0.350 200.370 4.280 ;
        RECT 201.210 0.350 201.750 4.280 ;
        RECT 202.590 0.350 203.130 4.280 ;
        RECT 203.970 0.350 204.510 4.280 ;
        RECT 205.350 0.350 205.890 4.280 ;
        RECT 206.730 0.350 207.270 4.280 ;
        RECT 208.110 0.350 208.650 4.280 ;
        RECT 209.490 0.350 210.030 4.280 ;
        RECT 210.870 0.350 211.410 4.280 ;
        RECT 212.250 0.350 212.790 4.280 ;
        RECT 213.630 0.350 214.170 4.280 ;
        RECT 215.010 0.350 215.550 4.280 ;
        RECT 216.390 0.350 216.930 4.280 ;
        RECT 217.770 0.350 218.310 4.280 ;
        RECT 219.150 0.350 219.690 4.280 ;
        RECT 220.530 0.350 221.070 4.280 ;
        RECT 221.910 0.350 222.450 4.280 ;
        RECT 223.290 0.350 223.830 4.280 ;
        RECT 224.670 0.350 225.210 4.280 ;
        RECT 226.050 0.350 226.590 4.280 ;
        RECT 227.430 0.350 227.970 4.280 ;
        RECT 228.810 0.350 229.350 4.280 ;
        RECT 230.190 0.350 230.730 4.280 ;
        RECT 231.570 0.350 232.110 4.280 ;
        RECT 232.950 0.350 233.490 4.280 ;
        RECT 234.330 0.350 234.870 4.280 ;
        RECT 235.710 0.350 236.250 4.280 ;
        RECT 237.090 0.350 237.630 4.280 ;
        RECT 238.470 0.350 239.010 4.280 ;
        RECT 239.850 0.350 240.390 4.280 ;
        RECT 241.230 0.350 241.770 4.280 ;
        RECT 242.610 0.350 243.150 4.280 ;
        RECT 243.990 0.350 244.530 4.280 ;
        RECT 245.370 0.350 245.910 4.280 ;
        RECT 246.750 0.350 247.290 4.280 ;
        RECT 248.130 0.350 248.670 4.280 ;
        RECT 249.510 0.350 250.050 4.280 ;
        RECT 250.890 0.350 251.430 4.280 ;
        RECT 252.270 0.350 252.810 4.280 ;
        RECT 253.650 0.350 254.190 4.280 ;
        RECT 255.030 0.350 255.570 4.280 ;
        RECT 256.410 0.350 256.950 4.280 ;
        RECT 257.790 0.350 258.330 4.280 ;
        RECT 259.170 0.350 259.710 4.280 ;
        RECT 260.550 0.350 261.090 4.280 ;
        RECT 261.930 0.350 262.470 4.280 ;
        RECT 263.310 0.350 263.850 4.280 ;
        RECT 264.690 0.350 265.230 4.280 ;
        RECT 266.070 0.350 266.610 4.280 ;
        RECT 267.450 0.350 267.990 4.280 ;
        RECT 268.830 0.350 269.370 4.280 ;
        RECT 270.210 0.350 298.900 4.280 ;
      LAYER met3 ;
        RECT 4.000 292.720 295.600 293.585 ;
        RECT 4.000 292.080 296.000 292.720 ;
        RECT 4.000 290.680 295.600 292.080 ;
        RECT 4.000 290.040 296.000 290.680 ;
        RECT 4.000 288.640 295.600 290.040 ;
        RECT 4.000 288.000 296.000 288.640 ;
        RECT 4.000 286.600 295.600 288.000 ;
        RECT 4.000 285.960 296.000 286.600 ;
        RECT 4.000 284.560 295.600 285.960 ;
        RECT 4.000 283.920 296.000 284.560 ;
        RECT 4.000 282.520 295.600 283.920 ;
        RECT 4.000 281.880 296.000 282.520 ;
        RECT 4.000 280.480 295.600 281.880 ;
        RECT 4.000 279.840 296.000 280.480 ;
        RECT 4.400 278.440 295.600 279.840 ;
        RECT 4.000 277.800 296.000 278.440 ;
        RECT 4.000 277.120 295.600 277.800 ;
        RECT 4.400 276.400 295.600 277.120 ;
        RECT 4.400 275.760 296.000 276.400 ;
        RECT 4.400 275.720 295.600 275.760 ;
        RECT 4.000 274.400 295.600 275.720 ;
        RECT 4.400 274.360 295.600 274.400 ;
        RECT 4.400 273.720 296.000 274.360 ;
        RECT 4.400 273.000 295.600 273.720 ;
        RECT 4.000 272.320 295.600 273.000 ;
        RECT 4.000 271.680 296.000 272.320 ;
        RECT 4.400 270.280 295.600 271.680 ;
        RECT 4.000 269.640 296.000 270.280 ;
        RECT 4.000 268.960 295.600 269.640 ;
        RECT 4.400 268.240 295.600 268.960 ;
        RECT 4.400 267.600 296.000 268.240 ;
        RECT 4.400 267.560 295.600 267.600 ;
        RECT 4.000 266.240 295.600 267.560 ;
        RECT 4.400 266.200 295.600 266.240 ;
        RECT 4.400 265.560 296.000 266.200 ;
        RECT 4.400 264.840 295.600 265.560 ;
        RECT 4.000 264.160 295.600 264.840 ;
        RECT 4.000 263.520 296.000 264.160 ;
        RECT 4.400 262.120 295.600 263.520 ;
        RECT 4.000 261.480 296.000 262.120 ;
        RECT 4.000 260.800 295.600 261.480 ;
        RECT 4.400 260.080 295.600 260.800 ;
        RECT 4.400 259.440 296.000 260.080 ;
        RECT 4.400 259.400 295.600 259.440 ;
        RECT 4.000 258.080 295.600 259.400 ;
        RECT 4.400 258.040 295.600 258.080 ;
        RECT 4.400 257.400 296.000 258.040 ;
        RECT 4.400 256.680 295.600 257.400 ;
        RECT 4.000 256.000 295.600 256.680 ;
        RECT 4.000 255.360 296.000 256.000 ;
        RECT 4.400 253.960 295.600 255.360 ;
        RECT 4.000 253.320 296.000 253.960 ;
        RECT 4.000 252.640 295.600 253.320 ;
        RECT 4.400 251.920 295.600 252.640 ;
        RECT 4.400 251.280 296.000 251.920 ;
        RECT 4.400 251.240 295.600 251.280 ;
        RECT 4.000 249.920 295.600 251.240 ;
        RECT 4.400 249.880 295.600 249.920 ;
        RECT 4.400 249.240 296.000 249.880 ;
        RECT 4.400 248.520 295.600 249.240 ;
        RECT 4.000 247.840 295.600 248.520 ;
        RECT 4.000 247.200 296.000 247.840 ;
        RECT 4.400 245.800 295.600 247.200 ;
        RECT 4.000 245.160 296.000 245.800 ;
        RECT 4.000 244.480 295.600 245.160 ;
        RECT 4.400 243.760 295.600 244.480 ;
        RECT 4.400 243.120 296.000 243.760 ;
        RECT 4.400 243.080 295.600 243.120 ;
        RECT 4.000 241.760 295.600 243.080 ;
        RECT 4.400 241.720 295.600 241.760 ;
        RECT 4.400 241.080 296.000 241.720 ;
        RECT 4.400 240.360 295.600 241.080 ;
        RECT 4.000 239.680 295.600 240.360 ;
        RECT 4.000 239.040 296.000 239.680 ;
        RECT 4.400 237.640 295.600 239.040 ;
        RECT 4.000 237.000 296.000 237.640 ;
        RECT 4.000 236.320 295.600 237.000 ;
        RECT 4.400 235.600 295.600 236.320 ;
        RECT 4.400 234.960 296.000 235.600 ;
        RECT 4.400 234.920 295.600 234.960 ;
        RECT 4.000 233.600 295.600 234.920 ;
        RECT 4.400 233.560 295.600 233.600 ;
        RECT 4.400 232.920 296.000 233.560 ;
        RECT 4.400 232.200 295.600 232.920 ;
        RECT 4.000 231.520 295.600 232.200 ;
        RECT 4.000 230.880 296.000 231.520 ;
        RECT 4.400 229.480 295.600 230.880 ;
        RECT 4.000 228.840 296.000 229.480 ;
        RECT 4.000 228.160 295.600 228.840 ;
        RECT 4.400 227.440 295.600 228.160 ;
        RECT 4.400 226.800 296.000 227.440 ;
        RECT 4.400 226.760 295.600 226.800 ;
        RECT 4.000 225.440 295.600 226.760 ;
        RECT 4.400 225.400 295.600 225.440 ;
        RECT 4.400 224.760 296.000 225.400 ;
        RECT 4.400 224.040 295.600 224.760 ;
        RECT 4.000 223.360 295.600 224.040 ;
        RECT 4.000 222.720 296.000 223.360 ;
        RECT 4.400 221.320 295.600 222.720 ;
        RECT 4.000 220.680 296.000 221.320 ;
        RECT 4.000 220.000 295.600 220.680 ;
        RECT 4.400 219.280 295.600 220.000 ;
        RECT 4.400 218.640 296.000 219.280 ;
        RECT 4.400 218.600 295.600 218.640 ;
        RECT 4.000 217.280 295.600 218.600 ;
        RECT 4.400 217.240 295.600 217.280 ;
        RECT 4.400 216.600 296.000 217.240 ;
        RECT 4.400 215.880 295.600 216.600 ;
        RECT 4.000 215.200 295.600 215.880 ;
        RECT 4.000 214.560 296.000 215.200 ;
        RECT 4.400 213.160 295.600 214.560 ;
        RECT 4.000 212.520 296.000 213.160 ;
        RECT 4.000 211.840 295.600 212.520 ;
        RECT 4.400 211.120 295.600 211.840 ;
        RECT 4.400 210.480 296.000 211.120 ;
        RECT 4.400 210.440 295.600 210.480 ;
        RECT 4.000 209.120 295.600 210.440 ;
        RECT 4.400 209.080 295.600 209.120 ;
        RECT 4.400 208.440 296.000 209.080 ;
        RECT 4.400 207.720 295.600 208.440 ;
        RECT 4.000 207.040 295.600 207.720 ;
        RECT 4.000 206.400 296.000 207.040 ;
        RECT 4.400 205.000 295.600 206.400 ;
        RECT 4.000 204.360 296.000 205.000 ;
        RECT 4.000 203.680 295.600 204.360 ;
        RECT 4.400 202.960 295.600 203.680 ;
        RECT 4.400 202.320 296.000 202.960 ;
        RECT 4.400 202.280 295.600 202.320 ;
        RECT 4.000 200.960 295.600 202.280 ;
        RECT 4.400 200.920 295.600 200.960 ;
        RECT 4.400 200.280 296.000 200.920 ;
        RECT 4.400 199.560 295.600 200.280 ;
        RECT 4.000 198.880 295.600 199.560 ;
        RECT 4.000 198.240 296.000 198.880 ;
        RECT 4.400 196.840 295.600 198.240 ;
        RECT 4.000 196.200 296.000 196.840 ;
        RECT 4.000 195.520 295.600 196.200 ;
        RECT 4.400 194.800 295.600 195.520 ;
        RECT 4.400 194.160 296.000 194.800 ;
        RECT 4.400 194.120 295.600 194.160 ;
        RECT 4.000 192.800 295.600 194.120 ;
        RECT 4.400 192.760 295.600 192.800 ;
        RECT 4.400 192.120 296.000 192.760 ;
        RECT 4.400 191.400 295.600 192.120 ;
        RECT 4.000 190.720 295.600 191.400 ;
        RECT 4.000 190.080 296.000 190.720 ;
        RECT 4.400 188.680 295.600 190.080 ;
        RECT 4.000 188.040 296.000 188.680 ;
        RECT 4.000 187.360 295.600 188.040 ;
        RECT 4.400 186.640 295.600 187.360 ;
        RECT 4.400 186.000 296.000 186.640 ;
        RECT 4.400 185.960 295.600 186.000 ;
        RECT 4.000 184.640 295.600 185.960 ;
        RECT 4.400 184.600 295.600 184.640 ;
        RECT 4.400 183.960 296.000 184.600 ;
        RECT 4.400 183.240 295.600 183.960 ;
        RECT 4.000 182.560 295.600 183.240 ;
        RECT 4.000 181.920 296.000 182.560 ;
        RECT 4.400 180.520 295.600 181.920 ;
        RECT 4.000 179.880 296.000 180.520 ;
        RECT 4.000 179.200 295.600 179.880 ;
        RECT 4.400 178.480 295.600 179.200 ;
        RECT 4.400 177.840 296.000 178.480 ;
        RECT 4.400 177.800 295.600 177.840 ;
        RECT 4.000 176.480 295.600 177.800 ;
        RECT 4.400 176.440 295.600 176.480 ;
        RECT 4.400 175.800 296.000 176.440 ;
        RECT 4.400 175.080 295.600 175.800 ;
        RECT 4.000 174.400 295.600 175.080 ;
        RECT 4.000 173.760 296.000 174.400 ;
        RECT 4.400 172.360 295.600 173.760 ;
        RECT 4.000 171.720 296.000 172.360 ;
        RECT 4.000 171.040 295.600 171.720 ;
        RECT 4.400 170.320 295.600 171.040 ;
        RECT 4.400 169.680 296.000 170.320 ;
        RECT 4.400 169.640 295.600 169.680 ;
        RECT 4.000 168.320 295.600 169.640 ;
        RECT 4.400 168.280 295.600 168.320 ;
        RECT 4.400 167.640 296.000 168.280 ;
        RECT 4.400 166.920 295.600 167.640 ;
        RECT 4.000 166.240 295.600 166.920 ;
        RECT 4.000 165.600 296.000 166.240 ;
        RECT 4.400 164.200 295.600 165.600 ;
        RECT 4.000 163.560 296.000 164.200 ;
        RECT 4.000 162.880 295.600 163.560 ;
        RECT 4.400 162.160 295.600 162.880 ;
        RECT 4.400 161.520 296.000 162.160 ;
        RECT 4.400 161.480 295.600 161.520 ;
        RECT 4.000 160.160 295.600 161.480 ;
        RECT 4.400 160.120 295.600 160.160 ;
        RECT 4.400 159.480 296.000 160.120 ;
        RECT 4.400 158.760 295.600 159.480 ;
        RECT 4.000 158.080 295.600 158.760 ;
        RECT 4.000 157.440 296.000 158.080 ;
        RECT 4.400 156.040 295.600 157.440 ;
        RECT 4.000 155.400 296.000 156.040 ;
        RECT 4.000 154.720 295.600 155.400 ;
        RECT 4.400 154.000 295.600 154.720 ;
        RECT 4.400 153.360 296.000 154.000 ;
        RECT 4.400 153.320 295.600 153.360 ;
        RECT 4.000 152.000 295.600 153.320 ;
        RECT 4.400 151.960 295.600 152.000 ;
        RECT 4.400 151.320 296.000 151.960 ;
        RECT 4.400 150.600 295.600 151.320 ;
        RECT 4.000 149.920 295.600 150.600 ;
        RECT 4.000 149.280 296.000 149.920 ;
        RECT 4.400 147.880 295.600 149.280 ;
        RECT 4.000 147.240 296.000 147.880 ;
        RECT 4.000 146.560 295.600 147.240 ;
        RECT 4.400 145.840 295.600 146.560 ;
        RECT 4.400 145.200 296.000 145.840 ;
        RECT 4.400 145.160 295.600 145.200 ;
        RECT 4.000 143.840 295.600 145.160 ;
        RECT 4.400 143.800 295.600 143.840 ;
        RECT 4.400 143.160 296.000 143.800 ;
        RECT 4.400 142.440 295.600 143.160 ;
        RECT 4.000 141.760 295.600 142.440 ;
        RECT 4.000 141.120 296.000 141.760 ;
        RECT 4.400 139.720 295.600 141.120 ;
        RECT 4.000 139.080 296.000 139.720 ;
        RECT 4.000 138.400 295.600 139.080 ;
        RECT 4.400 137.680 295.600 138.400 ;
        RECT 4.400 137.040 296.000 137.680 ;
        RECT 4.400 137.000 295.600 137.040 ;
        RECT 4.000 135.680 295.600 137.000 ;
        RECT 4.400 135.640 295.600 135.680 ;
        RECT 4.400 135.000 296.000 135.640 ;
        RECT 4.400 134.280 295.600 135.000 ;
        RECT 4.000 133.600 295.600 134.280 ;
        RECT 4.000 132.960 296.000 133.600 ;
        RECT 4.400 131.560 295.600 132.960 ;
        RECT 4.000 130.920 296.000 131.560 ;
        RECT 4.000 130.240 295.600 130.920 ;
        RECT 4.400 129.520 295.600 130.240 ;
        RECT 4.400 128.880 296.000 129.520 ;
        RECT 4.400 128.840 295.600 128.880 ;
        RECT 4.000 127.520 295.600 128.840 ;
        RECT 4.400 127.480 295.600 127.520 ;
        RECT 4.400 126.840 296.000 127.480 ;
        RECT 4.400 126.120 295.600 126.840 ;
        RECT 4.000 125.440 295.600 126.120 ;
        RECT 4.000 124.800 296.000 125.440 ;
        RECT 4.400 123.400 295.600 124.800 ;
        RECT 4.000 122.760 296.000 123.400 ;
        RECT 4.000 122.080 295.600 122.760 ;
        RECT 4.400 121.360 295.600 122.080 ;
        RECT 4.400 120.720 296.000 121.360 ;
        RECT 4.400 120.680 295.600 120.720 ;
        RECT 4.000 119.360 295.600 120.680 ;
        RECT 4.400 119.320 295.600 119.360 ;
        RECT 4.400 118.680 296.000 119.320 ;
        RECT 4.400 117.960 295.600 118.680 ;
        RECT 4.000 117.280 295.600 117.960 ;
        RECT 4.000 116.640 296.000 117.280 ;
        RECT 4.400 115.240 295.600 116.640 ;
        RECT 4.000 114.600 296.000 115.240 ;
        RECT 4.000 113.920 295.600 114.600 ;
        RECT 4.400 113.200 295.600 113.920 ;
        RECT 4.400 112.560 296.000 113.200 ;
        RECT 4.400 112.520 295.600 112.560 ;
        RECT 4.000 111.200 295.600 112.520 ;
        RECT 4.400 111.160 295.600 111.200 ;
        RECT 4.400 110.520 296.000 111.160 ;
        RECT 4.400 109.800 295.600 110.520 ;
        RECT 4.000 109.120 295.600 109.800 ;
        RECT 4.000 108.480 296.000 109.120 ;
        RECT 4.400 107.080 295.600 108.480 ;
        RECT 4.000 106.440 296.000 107.080 ;
        RECT 4.000 105.760 295.600 106.440 ;
        RECT 4.400 105.040 295.600 105.760 ;
        RECT 4.400 104.400 296.000 105.040 ;
        RECT 4.400 104.360 295.600 104.400 ;
        RECT 4.000 103.040 295.600 104.360 ;
        RECT 4.400 103.000 295.600 103.040 ;
        RECT 4.400 102.360 296.000 103.000 ;
        RECT 4.400 101.640 295.600 102.360 ;
        RECT 4.000 100.960 295.600 101.640 ;
        RECT 4.000 100.320 296.000 100.960 ;
        RECT 4.400 98.920 295.600 100.320 ;
        RECT 4.000 98.280 296.000 98.920 ;
        RECT 4.000 97.600 295.600 98.280 ;
        RECT 4.400 96.880 295.600 97.600 ;
        RECT 4.400 96.240 296.000 96.880 ;
        RECT 4.400 96.200 295.600 96.240 ;
        RECT 4.000 94.880 295.600 96.200 ;
        RECT 4.400 94.840 295.600 94.880 ;
        RECT 4.400 94.200 296.000 94.840 ;
        RECT 4.400 93.480 295.600 94.200 ;
        RECT 4.000 92.800 295.600 93.480 ;
        RECT 4.000 92.160 296.000 92.800 ;
        RECT 4.400 90.760 295.600 92.160 ;
        RECT 4.000 90.120 296.000 90.760 ;
        RECT 4.000 89.440 295.600 90.120 ;
        RECT 4.400 88.720 295.600 89.440 ;
        RECT 4.400 88.080 296.000 88.720 ;
        RECT 4.400 88.040 295.600 88.080 ;
        RECT 4.000 86.720 295.600 88.040 ;
        RECT 4.400 86.680 295.600 86.720 ;
        RECT 4.400 86.040 296.000 86.680 ;
        RECT 4.400 85.320 295.600 86.040 ;
        RECT 4.000 84.640 295.600 85.320 ;
        RECT 4.000 84.000 296.000 84.640 ;
        RECT 4.400 82.600 295.600 84.000 ;
        RECT 4.000 81.960 296.000 82.600 ;
        RECT 4.000 81.280 295.600 81.960 ;
        RECT 4.400 80.560 295.600 81.280 ;
        RECT 4.400 79.920 296.000 80.560 ;
        RECT 4.400 79.880 295.600 79.920 ;
        RECT 4.000 78.560 295.600 79.880 ;
        RECT 4.400 78.520 295.600 78.560 ;
        RECT 4.400 77.880 296.000 78.520 ;
        RECT 4.400 77.160 295.600 77.880 ;
        RECT 4.000 76.480 295.600 77.160 ;
        RECT 4.000 75.840 296.000 76.480 ;
        RECT 4.400 74.440 295.600 75.840 ;
        RECT 4.000 73.800 296.000 74.440 ;
        RECT 4.000 73.120 295.600 73.800 ;
        RECT 4.400 72.400 295.600 73.120 ;
        RECT 4.400 71.760 296.000 72.400 ;
        RECT 4.400 71.720 295.600 71.760 ;
        RECT 4.000 70.400 295.600 71.720 ;
        RECT 4.400 70.360 295.600 70.400 ;
        RECT 4.400 69.720 296.000 70.360 ;
        RECT 4.400 69.000 295.600 69.720 ;
        RECT 4.000 68.320 295.600 69.000 ;
        RECT 4.000 67.680 296.000 68.320 ;
        RECT 4.400 66.280 295.600 67.680 ;
        RECT 4.000 65.640 296.000 66.280 ;
        RECT 4.000 64.960 295.600 65.640 ;
        RECT 4.400 64.240 295.600 64.960 ;
        RECT 4.400 63.600 296.000 64.240 ;
        RECT 4.400 63.560 295.600 63.600 ;
        RECT 4.000 62.240 295.600 63.560 ;
        RECT 4.400 62.200 295.600 62.240 ;
        RECT 4.400 61.560 296.000 62.200 ;
        RECT 4.400 60.840 295.600 61.560 ;
        RECT 4.000 60.160 295.600 60.840 ;
        RECT 4.000 59.520 296.000 60.160 ;
        RECT 4.400 58.120 295.600 59.520 ;
        RECT 4.000 57.480 296.000 58.120 ;
        RECT 4.000 56.800 295.600 57.480 ;
        RECT 4.400 56.080 295.600 56.800 ;
        RECT 4.400 55.440 296.000 56.080 ;
        RECT 4.400 55.400 295.600 55.440 ;
        RECT 4.000 54.080 295.600 55.400 ;
        RECT 4.400 54.040 295.600 54.080 ;
        RECT 4.400 53.400 296.000 54.040 ;
        RECT 4.400 52.680 295.600 53.400 ;
        RECT 4.000 52.000 295.600 52.680 ;
        RECT 4.000 51.360 296.000 52.000 ;
        RECT 4.400 49.960 295.600 51.360 ;
        RECT 4.000 49.320 296.000 49.960 ;
        RECT 4.000 48.640 295.600 49.320 ;
        RECT 4.400 47.920 295.600 48.640 ;
        RECT 4.400 47.280 296.000 47.920 ;
        RECT 4.400 47.240 295.600 47.280 ;
        RECT 4.000 45.920 295.600 47.240 ;
        RECT 4.400 45.880 295.600 45.920 ;
        RECT 4.400 45.240 296.000 45.880 ;
        RECT 4.400 44.520 295.600 45.240 ;
        RECT 4.000 43.840 295.600 44.520 ;
        RECT 4.000 43.200 296.000 43.840 ;
        RECT 4.400 41.800 295.600 43.200 ;
        RECT 4.000 41.160 296.000 41.800 ;
        RECT 4.000 40.480 295.600 41.160 ;
        RECT 4.400 39.760 295.600 40.480 ;
        RECT 4.400 39.120 296.000 39.760 ;
        RECT 4.400 39.080 295.600 39.120 ;
        RECT 4.000 37.760 295.600 39.080 ;
        RECT 4.400 37.720 295.600 37.760 ;
        RECT 4.400 37.080 296.000 37.720 ;
        RECT 4.400 36.360 295.600 37.080 ;
        RECT 4.000 35.680 295.600 36.360 ;
        RECT 4.000 35.040 296.000 35.680 ;
        RECT 4.400 33.640 295.600 35.040 ;
        RECT 4.000 33.000 296.000 33.640 ;
        RECT 4.000 32.320 295.600 33.000 ;
        RECT 4.400 31.600 295.600 32.320 ;
        RECT 4.400 30.960 296.000 31.600 ;
        RECT 4.400 30.920 295.600 30.960 ;
        RECT 4.000 29.600 295.600 30.920 ;
        RECT 4.400 29.560 295.600 29.600 ;
        RECT 4.400 28.920 296.000 29.560 ;
        RECT 4.400 28.200 295.600 28.920 ;
        RECT 4.000 27.520 295.600 28.200 ;
        RECT 4.000 26.880 296.000 27.520 ;
        RECT 4.400 25.480 295.600 26.880 ;
        RECT 4.000 24.840 296.000 25.480 ;
        RECT 4.000 24.160 295.600 24.840 ;
        RECT 4.400 23.440 295.600 24.160 ;
        RECT 4.400 22.800 296.000 23.440 ;
        RECT 4.400 22.760 295.600 22.800 ;
        RECT 4.000 21.440 295.600 22.760 ;
        RECT 4.400 21.400 295.600 21.440 ;
        RECT 4.400 20.760 296.000 21.400 ;
        RECT 4.400 20.040 295.600 20.760 ;
        RECT 4.000 19.360 295.600 20.040 ;
        RECT 4.000 18.720 296.000 19.360 ;
        RECT 4.000 17.320 295.600 18.720 ;
        RECT 4.000 16.680 296.000 17.320 ;
        RECT 4.000 15.280 295.600 16.680 ;
        RECT 4.000 14.640 296.000 15.280 ;
        RECT 4.000 13.240 295.600 14.640 ;
        RECT 4.000 12.600 296.000 13.240 ;
        RECT 4.000 11.200 295.600 12.600 ;
        RECT 4.000 10.560 296.000 11.200 ;
        RECT 4.000 9.160 295.600 10.560 ;
        RECT 4.000 8.520 296.000 9.160 ;
        RECT 4.000 7.120 295.600 8.520 ;
        RECT 4.000 6.480 296.000 7.120 ;
        RECT 4.000 5.615 295.600 6.480 ;
      LAYER met4 ;
        RECT 147.495 11.735 174.240 283.385 ;
        RECT 176.640 11.735 244.425 283.385 ;
  END
END multiplexer
END LIBRARY

