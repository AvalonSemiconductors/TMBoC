magic
tech sky130B
magscale 1 2
timestamp 1680007426
<< obsli1 >>
rect 1104 2159 18860 17425
<< obsm1 >>
rect 842 2128 19122 17456
<< metal2 >>
rect 4986 19200 5042 20000
rect 14922 19200 14978 20000
rect 846 0 902 800
rect 2502 0 2558 800
rect 4158 0 4214 800
rect 5814 0 5870 800
rect 7470 0 7526 800
rect 9126 0 9182 800
rect 10782 0 10838 800
rect 12438 0 12494 800
rect 14094 0 14150 800
rect 15750 0 15806 800
rect 17406 0 17462 800
rect 19062 0 19118 800
<< obsm2 >>
rect 848 19144 4930 19200
rect 5098 19144 14866 19200
rect 15034 19144 19116 19200
rect 848 856 19116 19144
rect 958 800 2446 856
rect 2614 800 4102 856
rect 4270 800 5758 856
rect 5926 800 7414 856
rect 7582 800 9070 856
rect 9238 800 10726 856
rect 10894 800 12382 856
rect 12550 800 14038 856
rect 14206 800 15694 856
rect 15862 800 17350 856
rect 17518 800 19006 856
<< obsm3 >>
rect 3165 2143 19017 17441
<< metal4 >>
rect 3163 2128 3483 17456
rect 5382 2128 5702 17456
rect 7602 2128 7922 17456
rect 9821 2128 10141 17456
rect 12041 2128 12361 17456
rect 14260 2128 14580 17456
rect 16480 2128 16800 17456
rect 18699 2128 19019 17456
<< labels >>
rlabel metal2 s 4986 19200 5042 20000 6 clk
port 1 nsew signal input
rlabel metal2 s 846 0 902 800 6 io_out[0]
port 2 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 io_out[10]
port 3 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 io_out[11]
port 4 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 io_out[1]
port 5 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 io_out[2]
port 6 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 io_out[3]
port 7 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 io_out[4]
port 8 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 io_out[5]
port 9 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 io_out[6]
port 10 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 io_out[7]
port 11 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 io_out[8]
port 12 nsew signal output
rlabel metal2 s 15750 0 15806 800 6 io_out[9]
port 13 nsew signal output
rlabel metal2 s 14922 19200 14978 20000 6 rst
port 14 nsew signal input
rlabel metal4 s 3163 2128 3483 17456 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 7602 2128 7922 17456 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 12041 2128 12361 17456 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 16480 2128 16800 17456 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 5382 2128 5702 17456 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 9821 2128 10141 17456 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 14260 2128 14580 17456 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 18699 2128 19019 17456 6 vssd1
port 16 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 741110
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/MultiplexedCounter/runs/23_03_28_14_42/results/signoff/tt2_tholin_multiplexed_counter.magic.gds
string GDS_START 270124
<< end >>

