magic
tech sky130B
magscale 1 2
timestamp 1676498274
<< obsli1 >>
rect 1104 2159 68816 67473
<< obsm1 >>
rect 1104 2128 68816 67504
<< metal2 >>
rect 8730 0 8842 800
rect 26210 0 26322 800
rect 43690 0 43802 800
rect 61170 0 61282 800
<< obsm2 >>
rect 1400 856 68336 67493
rect 1400 800 8674 856
rect 8898 800 26154 856
rect 26378 800 43634 856
rect 43858 800 61114 856
rect 61338 800 68336 856
<< metal3 >>
rect 0 62508 800 62748
rect 0 48636 800 48876
rect 0 34764 800 35004
rect 0 20892 800 21132
rect 0 7020 800 7260
<< obsm3 >>
rect 800 62828 65966 67489
rect 880 62428 65966 62828
rect 800 48956 65966 62428
rect 880 48556 65966 48956
rect 800 35084 65966 48556
rect 880 34684 65966 35084
rect 800 21212 65966 34684
rect 880 20812 65966 21212
rect 800 7340 65966 20812
rect 880 6940 65966 7340
rect 800 2143 65966 6940
<< metal4 >>
rect 4208 2128 4528 67504
rect 19568 2128 19888 67504
rect 34928 2128 35248 67504
rect 50288 2128 50608 67504
rect 65648 2128 65968 67504
<< obsm4 >>
rect 3187 3435 4128 58037
rect 4608 3435 19488 58037
rect 19968 3435 34848 58037
rect 35328 3435 50208 58037
rect 50688 3435 57901 58037
<< labels >>
rlabel metal3 s 0 48636 800 48876 6 clk
port 1 nsew signal input
rlabel metal3 s 0 7020 800 7260 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 0 20892 800 21132 6 io_in[1]
port 3 nsew signal input
rlabel metal3 s 0 34764 800 35004 6 io_in[2]
port 4 nsew signal input
rlabel metal2 s 8730 0 8842 800 6 io_out[0]
port 5 nsew signal output
rlabel metal2 s 26210 0 26322 800 6 io_out[1]
port 6 nsew signal output
rlabel metal2 s 43690 0 43802 800 6 io_out[2]
port 7 nsew signal output
rlabel metal2 s 61170 0 61282 800 6 io_out[3]
port 8 nsew signal output
rlabel metal3 s 0 62508 800 62748 6 rst
port 9 nsew signal input
rlabel metal4 s 4208 2128 4528 67504 6 vccd1
port 10 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 67504 6 vccd1
port 10 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 67504 6 vccd1
port 10 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 67504 6 vssd1
port 11 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 67504 6 vssd1
port 11 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 70000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 13871292
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/PositUnit/runs/23_02_15_22_39/results/signoff/posit_unit.magic.gds
string GDS_START 1199032
<< end >>

