VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_as1802
  CLASS BLOCK ;
  FOREIGN wrapped_as1802 ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 350.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 346.000 313.170 350.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 346.000 14.170 350.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 346.000 244.170 350.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 346.000 267.170 350.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 346.000 290.170 350.000 ;
    END
  END io_in[12]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 346.000 37.170 350.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 346.000 60.170 350.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 346.000 83.170 350.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 346.000 106.170 350.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 346.000 129.170 350.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 346.000 152.170 350.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 346.000 175.170 350.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 346.000 198.170 350.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 346.000 221.170 350.000 ;
    END
  END io_in[9]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 339.360 350.000 339.960 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 8.880 350.000 9.480 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 131.280 350.000 131.880 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 143.520 350.000 144.120 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 155.760 350.000 156.360 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 168.000 350.000 168.600 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 180.240 350.000 180.840 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 192.480 350.000 193.080 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 204.720 350.000 205.320 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 216.960 350.000 217.560 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 229.200 350.000 229.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 241.440 350.000 242.040 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 21.120 350.000 21.720 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 253.680 350.000 254.280 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 265.920 350.000 266.520 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 278.160 350.000 278.760 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 290.400 350.000 291.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 302.640 350.000 303.240 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 314.880 350.000 315.480 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 327.120 350.000 327.720 ;
    END
  END io_out[26]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 33.360 350.000 33.960 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 45.600 350.000 46.200 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 57.840 350.000 58.440 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 70.080 350.000 70.680 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 82.320 350.000 82.920 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 94.560 350.000 95.160 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 106.800 350.000 107.400 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 119.040 350.000 119.640 ;
    END
  END io_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 346.000 336.170 350.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 337.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 337.520 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 333.145 344.270 335.975 ;
        RECT 5.330 327.705 344.270 330.535 ;
        RECT 5.330 322.265 344.270 325.095 ;
        RECT 5.330 316.825 344.270 319.655 ;
        RECT 5.330 311.385 344.270 314.215 ;
        RECT 5.330 305.945 344.270 308.775 ;
        RECT 5.330 300.505 344.270 303.335 ;
        RECT 5.330 295.065 344.270 297.895 ;
        RECT 5.330 289.625 344.270 292.455 ;
        RECT 5.330 284.185 344.270 287.015 ;
        RECT 5.330 278.745 344.270 281.575 ;
        RECT 5.330 273.305 344.270 276.135 ;
        RECT 5.330 267.865 344.270 270.695 ;
        RECT 5.330 262.425 344.270 265.255 ;
        RECT 5.330 256.985 344.270 259.815 ;
        RECT 5.330 251.545 344.270 254.375 ;
        RECT 5.330 246.105 344.270 248.935 ;
        RECT 5.330 240.665 344.270 243.495 ;
        RECT 5.330 235.225 344.270 238.055 ;
        RECT 5.330 229.785 344.270 232.615 ;
        RECT 5.330 224.345 344.270 227.175 ;
        RECT 5.330 218.905 344.270 221.735 ;
        RECT 5.330 213.465 344.270 216.295 ;
        RECT 5.330 208.025 344.270 210.855 ;
        RECT 5.330 202.585 344.270 205.415 ;
        RECT 5.330 197.145 344.270 199.975 ;
        RECT 5.330 191.705 344.270 194.535 ;
        RECT 5.330 186.265 344.270 189.095 ;
        RECT 5.330 180.825 344.270 183.655 ;
        RECT 5.330 175.385 344.270 178.215 ;
        RECT 5.330 169.945 344.270 172.775 ;
        RECT 5.330 164.505 344.270 167.335 ;
        RECT 5.330 159.065 344.270 161.895 ;
        RECT 5.330 153.625 344.270 156.455 ;
        RECT 5.330 148.185 344.270 151.015 ;
        RECT 5.330 142.745 344.270 145.575 ;
        RECT 5.330 137.305 344.270 140.135 ;
        RECT 5.330 131.865 344.270 134.695 ;
        RECT 5.330 126.425 344.270 129.255 ;
        RECT 5.330 120.985 344.270 123.815 ;
        RECT 5.330 115.545 344.270 118.375 ;
        RECT 5.330 110.105 344.270 112.935 ;
        RECT 5.330 104.665 344.270 107.495 ;
        RECT 5.330 99.225 344.270 102.055 ;
        RECT 5.330 93.785 344.270 96.615 ;
        RECT 5.330 88.345 344.270 91.175 ;
        RECT 5.330 82.905 344.270 85.735 ;
        RECT 5.330 77.465 344.270 80.295 ;
        RECT 5.330 72.025 344.270 74.855 ;
        RECT 5.330 66.585 344.270 69.415 ;
        RECT 5.330 61.145 344.270 63.975 ;
        RECT 5.330 55.705 344.270 58.535 ;
        RECT 5.330 50.265 344.270 53.095 ;
        RECT 5.330 44.825 344.270 47.655 ;
        RECT 5.330 39.385 344.270 42.215 ;
        RECT 5.330 33.945 344.270 36.775 ;
        RECT 5.330 28.505 344.270 31.335 ;
        RECT 5.330 23.065 344.270 25.895 ;
        RECT 5.330 17.625 344.270 20.455 ;
        RECT 5.330 12.185 344.270 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 344.080 337.365 ;
      LAYER met1 ;
        RECT 5.520 10.640 345.390 345.740 ;
      LAYER met2 ;
        RECT 14.450 345.720 36.610 346.530 ;
        RECT 37.450 345.720 59.610 346.530 ;
        RECT 60.450 345.720 82.610 346.530 ;
        RECT 83.450 345.720 105.610 346.530 ;
        RECT 106.450 345.720 128.610 346.530 ;
        RECT 129.450 345.720 151.610 346.530 ;
        RECT 152.450 345.720 174.610 346.530 ;
        RECT 175.450 345.720 197.610 346.530 ;
        RECT 198.450 345.720 220.610 346.530 ;
        RECT 221.450 345.720 243.610 346.530 ;
        RECT 244.450 345.720 266.610 346.530 ;
        RECT 267.450 345.720 289.610 346.530 ;
        RECT 290.450 345.720 312.610 346.530 ;
        RECT 313.450 345.720 335.610 346.530 ;
        RECT 336.450 345.720 345.370 346.530 ;
        RECT 14.170 8.995 345.370 345.720 ;
      LAYER met3 ;
        RECT 21.050 338.960 345.600 339.825 ;
        RECT 21.050 328.120 346.000 338.960 ;
        RECT 21.050 326.720 345.600 328.120 ;
        RECT 21.050 315.880 346.000 326.720 ;
        RECT 21.050 314.480 345.600 315.880 ;
        RECT 21.050 303.640 346.000 314.480 ;
        RECT 21.050 302.240 345.600 303.640 ;
        RECT 21.050 291.400 346.000 302.240 ;
        RECT 21.050 290.000 345.600 291.400 ;
        RECT 21.050 279.160 346.000 290.000 ;
        RECT 21.050 277.760 345.600 279.160 ;
        RECT 21.050 266.920 346.000 277.760 ;
        RECT 21.050 265.520 345.600 266.920 ;
        RECT 21.050 254.680 346.000 265.520 ;
        RECT 21.050 253.280 345.600 254.680 ;
        RECT 21.050 242.440 346.000 253.280 ;
        RECT 21.050 241.040 345.600 242.440 ;
        RECT 21.050 230.200 346.000 241.040 ;
        RECT 21.050 228.800 345.600 230.200 ;
        RECT 21.050 217.960 346.000 228.800 ;
        RECT 21.050 216.560 345.600 217.960 ;
        RECT 21.050 205.720 346.000 216.560 ;
        RECT 21.050 204.320 345.600 205.720 ;
        RECT 21.050 193.480 346.000 204.320 ;
        RECT 21.050 192.080 345.600 193.480 ;
        RECT 21.050 181.240 346.000 192.080 ;
        RECT 21.050 179.840 345.600 181.240 ;
        RECT 21.050 169.000 346.000 179.840 ;
        RECT 21.050 167.600 345.600 169.000 ;
        RECT 21.050 156.760 346.000 167.600 ;
        RECT 21.050 155.360 345.600 156.760 ;
        RECT 21.050 144.520 346.000 155.360 ;
        RECT 21.050 143.120 345.600 144.520 ;
        RECT 21.050 132.280 346.000 143.120 ;
        RECT 21.050 130.880 345.600 132.280 ;
        RECT 21.050 120.040 346.000 130.880 ;
        RECT 21.050 118.640 345.600 120.040 ;
        RECT 21.050 107.800 346.000 118.640 ;
        RECT 21.050 106.400 345.600 107.800 ;
        RECT 21.050 95.560 346.000 106.400 ;
        RECT 21.050 94.160 345.600 95.560 ;
        RECT 21.050 83.320 346.000 94.160 ;
        RECT 21.050 81.920 345.600 83.320 ;
        RECT 21.050 71.080 346.000 81.920 ;
        RECT 21.050 69.680 345.600 71.080 ;
        RECT 21.050 58.840 346.000 69.680 ;
        RECT 21.050 57.440 345.600 58.840 ;
        RECT 21.050 46.600 346.000 57.440 ;
        RECT 21.050 45.200 345.600 46.600 ;
        RECT 21.050 34.360 346.000 45.200 ;
        RECT 21.050 32.960 345.600 34.360 ;
        RECT 21.050 22.120 346.000 32.960 ;
        RECT 21.050 20.720 345.600 22.120 ;
        RECT 21.050 9.880 346.000 20.720 ;
        RECT 21.050 9.015 345.600 9.880 ;
      LAYER met4 ;
        RECT 92.295 47.775 97.440 324.865 ;
        RECT 99.840 47.775 174.240 324.865 ;
        RECT 176.640 47.775 251.040 324.865 ;
        RECT 253.440 47.775 297.785 324.865 ;
  END
END wrapped_as1802
END LIBRARY

