magic
tech sky130B
magscale 1 2
timestamp 1680002326
<< viali >>
rect 32505 37417 32539 37451
rect 12081 37349 12115 37383
rect 28641 37349 28675 37383
rect 5457 37281 5491 37315
rect 9413 37281 9447 37315
rect 38301 37281 38335 37315
rect 5273 37213 5307 37247
rect 9229 37213 9263 37247
rect 11897 37213 11931 37247
rect 15209 37213 15243 37247
rect 18521 37213 18555 37247
rect 25145 37213 25179 37247
rect 28457 37213 28491 37247
rect 32413 37213 32447 37247
rect 35081 37213 35115 37247
rect 38117 37213 38151 37247
rect 22109 37145 22143 37179
rect 15301 37077 15335 37111
rect 18613 37077 18647 37111
rect 22201 37077 22235 37111
rect 25237 37077 25271 37111
rect 35173 37077 35207 37111
rect 14289 36873 14323 36907
rect 14197 36805 14231 36839
rect 18613 36737 18647 36771
rect 19073 36737 19107 36771
rect 25145 36737 25179 36771
rect 25973 36737 26007 36771
rect 26157 36737 26191 36771
rect 30113 36737 30147 36771
rect 30297 36737 30331 36771
rect 14473 36669 14507 36703
rect 25053 36669 25087 36703
rect 25513 36601 25547 36635
rect 13829 36533 13863 36567
rect 25973 36533 26007 36567
rect 30113 36533 30147 36567
rect 24869 36329 24903 36363
rect 30849 36329 30883 36363
rect 31033 36329 31067 36363
rect 14565 36261 14599 36295
rect 37013 36261 37047 36295
rect 14933 36193 14967 36227
rect 17233 36193 17267 36227
rect 25881 36193 25915 36227
rect 26065 36193 26099 36227
rect 29745 36193 29779 36227
rect 33241 36193 33275 36227
rect 17325 36125 17359 36159
rect 17509 36125 17543 36159
rect 24777 36125 24811 36159
rect 29009 36125 29043 36159
rect 29193 36125 29227 36159
rect 30021 36125 30055 36159
rect 30205 36125 30239 36159
rect 33333 36125 33367 36159
rect 34161 36125 34195 36159
rect 37197 36125 37231 36159
rect 15117 36057 15151 36091
rect 17969 36057 18003 36091
rect 25789 36057 25823 36091
rect 30665 36057 30699 36091
rect 15025 35989 15059 36023
rect 25421 35989 25455 36023
rect 29193 35989 29227 36023
rect 29929 35989 29963 36023
rect 30865 35989 30899 36023
rect 33701 35989 33735 36023
rect 34253 35989 34287 36023
rect 14289 35785 14323 35819
rect 21465 35785 21499 35819
rect 22569 35785 22603 35819
rect 34805 35785 34839 35819
rect 14197 35717 14231 35751
rect 29009 35717 29043 35751
rect 30297 35717 30331 35751
rect 31401 35717 31435 35751
rect 18797 35649 18831 35683
rect 19441 35649 19475 35683
rect 21281 35649 21315 35683
rect 21465 35649 21499 35683
rect 22385 35649 22419 35683
rect 23213 35649 23247 35683
rect 23397 35649 23431 35683
rect 25789 35649 25823 35683
rect 28917 35649 28951 35683
rect 29101 35649 29135 35683
rect 29837 35649 29871 35683
rect 29929 35649 29963 35683
rect 31217 35649 31251 35683
rect 31493 35649 31527 35683
rect 32965 35649 32999 35683
rect 33517 35649 33551 35683
rect 33793 35649 33827 35683
rect 34713 35649 34747 35683
rect 14473 35581 14507 35615
rect 22661 35581 22695 35615
rect 24961 35581 24995 35615
rect 25513 35581 25547 35615
rect 25973 35581 26007 35615
rect 30021 35581 30055 35615
rect 20269 35513 20303 35547
rect 23489 35513 23523 35547
rect 30757 35513 30791 35547
rect 13829 35445 13863 35479
rect 22109 35445 22143 35479
rect 31217 35445 31251 35479
rect 33149 35445 33183 35479
rect 20085 35241 20119 35275
rect 21281 35241 21315 35275
rect 21741 35241 21775 35275
rect 23213 35241 23247 35275
rect 24777 35241 24811 35275
rect 31953 35241 31987 35275
rect 20361 35173 20395 35207
rect 20453 35173 20487 35207
rect 18889 35105 18923 35139
rect 22753 35105 22787 35139
rect 27261 35105 27295 35139
rect 30297 35105 30331 35139
rect 33057 35105 33091 35139
rect 34253 35105 34287 35139
rect 35081 35105 35115 35139
rect 18429 35037 18463 35071
rect 18705 35037 18739 35071
rect 20269 35037 20303 35071
rect 20567 35037 20601 35071
rect 20729 35031 20763 35065
rect 21189 35037 21223 35071
rect 21557 35037 21591 35071
rect 22477 35037 22511 35071
rect 22661 35037 22695 35071
rect 23213 35037 23247 35071
rect 23305 35037 23339 35071
rect 24961 35037 24995 35071
rect 25053 35037 25087 35071
rect 26433 35037 26467 35071
rect 26801 35037 26835 35071
rect 30205 35037 30239 35071
rect 32137 35037 32171 35071
rect 32413 35037 32447 35071
rect 32781 35037 32815 35071
rect 33241 35037 33275 35071
rect 34161 35037 34195 35071
rect 34345 35037 34379 35071
rect 35173 35037 35207 35071
rect 22293 34969 22327 35003
rect 24777 34969 24811 35003
rect 23581 34901 23615 34935
rect 29745 34901 29779 34935
rect 30113 34901 30147 34935
rect 36001 34901 36035 34935
rect 18797 34697 18831 34731
rect 30021 34697 30055 34731
rect 32597 34697 32631 34731
rect 17417 34561 17451 34595
rect 18153 34561 18187 34595
rect 18245 34561 18279 34595
rect 18797 34561 18831 34595
rect 20269 34561 20303 34595
rect 20361 34561 20395 34595
rect 20729 34561 20763 34595
rect 21373 34561 21407 34595
rect 22017 34561 22051 34595
rect 22201 34561 22235 34595
rect 23962 34563 23996 34597
rect 24225 34561 24259 34595
rect 24317 34561 24351 34595
rect 24593 34561 24627 34595
rect 24777 34561 24811 34595
rect 25605 34561 25639 34595
rect 29837 34561 29871 34595
rect 30021 34561 30055 34595
rect 32321 34561 32355 34595
rect 33149 34561 33183 34595
rect 33517 34561 33551 34595
rect 25421 34493 25455 34527
rect 25789 34493 25823 34527
rect 32597 34493 32631 34527
rect 22385 34425 22419 34459
rect 34345 34425 34379 34459
rect 21465 34357 21499 34391
rect 23581 34357 23615 34391
rect 32413 34357 32447 34391
rect 16957 34153 16991 34187
rect 32781 34153 32815 34187
rect 26801 34085 26835 34119
rect 17325 34017 17359 34051
rect 18705 34017 18739 34051
rect 17141 33949 17175 33983
rect 17233 33949 17267 33983
rect 17417 33949 17451 33983
rect 17969 33949 18003 33983
rect 18061 33949 18095 33983
rect 18245 33949 18279 33983
rect 21189 33949 21223 33983
rect 21373 33949 21407 33983
rect 21649 33949 21683 33983
rect 21925 33949 21959 33983
rect 22201 33949 22235 33983
rect 25421 33949 25455 33983
rect 25789 33949 25823 33983
rect 26433 33949 26467 33983
rect 32689 33949 32723 33983
rect 20821 33881 20855 33915
rect 32505 33881 32539 33915
rect 25053 33609 25087 33643
rect 32781 33609 32815 33643
rect 16313 33541 16347 33575
rect 19441 33541 19475 33575
rect 31585 33541 31619 33575
rect 16037 33473 16071 33507
rect 16221 33473 16255 33507
rect 17233 33473 17267 33507
rect 17509 33473 17543 33507
rect 17693 33473 17727 33507
rect 18337 33473 18371 33507
rect 18889 33473 18923 33507
rect 19073 33473 19107 33507
rect 25053 33473 25087 33507
rect 26433 33473 26467 33507
rect 27353 33473 27387 33507
rect 27905 33473 27939 33507
rect 29745 33473 29779 33507
rect 30113 33473 30147 33507
rect 32597 33473 32631 33507
rect 17049 33405 17083 33439
rect 18153 33405 18187 33439
rect 24869 33405 24903 33439
rect 25421 33405 25455 33439
rect 32413 33405 32447 33439
rect 26525 33269 26559 33303
rect 16957 33065 16991 33099
rect 24685 33065 24719 33099
rect 25789 33065 25823 33099
rect 26985 33065 27019 33099
rect 23397 32997 23431 33031
rect 24961 32997 24995 33031
rect 28365 32997 28399 33031
rect 16589 32929 16623 32963
rect 18153 32929 18187 32963
rect 23581 32929 23615 32963
rect 25053 32929 25087 32963
rect 16773 32861 16807 32895
rect 17785 32861 17819 32895
rect 17969 32861 18003 32895
rect 23121 32861 23155 32895
rect 24869 32861 24903 32895
rect 25145 32861 25179 32895
rect 25329 32861 25363 32895
rect 25973 32861 26007 32895
rect 26065 32861 26099 32895
rect 26249 32861 26283 32895
rect 26341 32861 26375 32895
rect 27169 32861 27203 32895
rect 27261 32861 27295 32895
rect 27445 32861 27479 32895
rect 27537 32861 27571 32895
rect 28089 32861 28123 32895
rect 28641 32861 28675 32895
rect 28917 32861 28951 32895
rect 17509 32521 17543 32555
rect 18705 32521 18739 32555
rect 28089 32521 28123 32555
rect 18337 32453 18371 32487
rect 18553 32453 18587 32487
rect 21097 32453 21131 32487
rect 28917 32453 28951 32487
rect 34161 32453 34195 32487
rect 17509 32385 17543 32419
rect 20821 32385 20855 32419
rect 21005 32385 21039 32419
rect 23121 32385 23155 32419
rect 23489 32385 23523 32419
rect 27261 32385 27295 32419
rect 27353 32385 27387 32419
rect 27997 32385 28031 32419
rect 28273 32385 28307 32419
rect 28825 32385 28859 32419
rect 29009 32385 29043 32419
rect 33885 32385 33919 32419
rect 34621 32385 34655 32419
rect 34805 32385 34839 32419
rect 35265 32385 35299 32419
rect 17325 32317 17359 32351
rect 17877 32317 17911 32351
rect 34161 32317 34195 32351
rect 35357 32317 35391 32351
rect 27261 32249 27295 32283
rect 18521 32181 18555 32215
rect 33977 32181 34011 32215
rect 34621 32181 34655 32215
rect 23581 31977 23615 32011
rect 17693 31909 17727 31943
rect 23397 31909 23431 31943
rect 23121 31841 23155 31875
rect 27721 31841 27755 31875
rect 34253 31841 34287 31875
rect 35449 31841 35483 31875
rect 14381 31773 14415 31807
rect 17509 31773 17543 31807
rect 17693 31773 17727 31807
rect 27629 31773 27663 31807
rect 27813 31773 27847 31807
rect 33517 31773 33551 31807
rect 33701 31773 33735 31807
rect 34161 31773 34195 31807
rect 34345 31773 34379 31807
rect 35357 31773 35391 31807
rect 14933 31705 14967 31739
rect 33701 31637 33735 31671
rect 34897 31637 34931 31671
rect 35265 31637 35299 31671
rect 17233 31433 17267 31467
rect 12909 31365 12943 31399
rect 15301 31365 15335 31399
rect 30573 31365 30607 31399
rect 34529 31365 34563 31399
rect 5273 31297 5307 31331
rect 12633 31297 12667 31331
rect 15025 31297 15059 31331
rect 15117 31297 15151 31331
rect 17141 31297 17175 31331
rect 19717 31297 19751 31331
rect 19809 31297 19843 31331
rect 19993 31297 20027 31331
rect 20545 31297 20579 31331
rect 22385 31297 22419 31331
rect 23397 31297 23431 31331
rect 30389 31297 30423 31331
rect 30665 31297 30699 31331
rect 34069 31297 34103 31331
rect 34161 31297 34195 31331
rect 5549 31229 5583 31263
rect 19165 31229 19199 31263
rect 20269 31229 20303 31263
rect 33793 31229 33827 31263
rect 5365 31161 5399 31195
rect 23213 31161 23247 31195
rect 34713 31161 34747 31195
rect 5457 31093 5491 31127
rect 14381 31093 14415 31127
rect 22385 31093 22419 31127
rect 30205 31093 30239 31127
rect 33885 30889 33919 30923
rect 14381 30821 14415 30855
rect 21097 30821 21131 30855
rect 29101 30821 29135 30855
rect 35449 30821 35483 30855
rect 4353 30753 4387 30787
rect 11069 30753 11103 30787
rect 30021 30753 30055 30787
rect 30113 30753 30147 30787
rect 31125 30753 31159 30787
rect 31217 30753 31251 30787
rect 34989 30753 35023 30787
rect 4629 30685 4663 30719
rect 9873 30685 9907 30719
rect 10885 30685 10919 30719
rect 14381 30685 14415 30719
rect 14565 30685 14599 30719
rect 18153 30685 18187 30719
rect 18429 30685 18463 30719
rect 19901 30685 19935 30719
rect 19993 30685 20027 30719
rect 20361 30685 20395 30719
rect 20913 30685 20947 30719
rect 21189 30685 21223 30719
rect 29929 30685 29963 30719
rect 30205 30685 30239 30719
rect 30941 30685 30975 30719
rect 31033 30685 31067 30719
rect 33793 30685 33827 30719
rect 33977 30685 34011 30719
rect 35081 30685 35115 30719
rect 6009 30617 6043 30651
rect 9689 30617 9723 30651
rect 28733 30617 28767 30651
rect 10057 30549 10091 30583
rect 17969 30549 18003 30583
rect 18337 30549 18371 30583
rect 29193 30549 29227 30583
rect 29745 30549 29779 30583
rect 30757 30549 30791 30583
rect 4813 30345 4847 30379
rect 18889 30345 18923 30379
rect 20846 30345 20880 30379
rect 5457 30277 5491 30311
rect 6745 30277 6779 30311
rect 10241 30277 10275 30311
rect 17233 30277 17267 30311
rect 28365 30277 28399 30311
rect 32413 30277 32447 30311
rect 33793 30277 33827 30311
rect 5089 30209 5123 30243
rect 6561 30209 6595 30243
rect 6837 30209 6871 30243
rect 8769 30209 8803 30243
rect 8953 30209 8987 30243
rect 10977 30209 11011 30243
rect 15117 30209 15151 30243
rect 15301 30209 15335 30243
rect 17141 30209 17175 30243
rect 17325 30209 17359 30243
rect 20545 30209 20579 30243
rect 20729 30209 20763 30243
rect 21281 30209 21315 30243
rect 24317 30209 24351 30243
rect 24501 30209 24535 30243
rect 28181 30209 28215 30243
rect 28457 30209 28491 30243
rect 29469 30209 29503 30243
rect 29653 30209 29687 30243
rect 29837 30209 29871 30243
rect 30573 30209 30607 30243
rect 30757 30209 30791 30243
rect 32321 30209 32355 30243
rect 32689 30209 32723 30243
rect 32965 30209 32999 30243
rect 33609 30209 33643 30243
rect 33885 30209 33919 30243
rect 4997 30141 5031 30175
rect 5365 30141 5399 30175
rect 9689 30141 9723 30175
rect 12817 30141 12851 30175
rect 13093 30141 13127 30175
rect 17877 30141 17911 30175
rect 33425 30141 33459 30175
rect 6561 30073 6595 30107
rect 29285 30073 29319 30107
rect 8861 30005 8895 30039
rect 11069 30005 11103 30039
rect 14565 30005 14599 30039
rect 15209 30005 15243 30039
rect 24317 30005 24351 30039
rect 28181 30005 28215 30039
rect 30665 30005 30699 30039
rect 6469 29801 6503 29835
rect 7573 29801 7607 29835
rect 18521 29801 18555 29835
rect 24777 29801 24811 29835
rect 24961 29801 24995 29835
rect 28457 29801 28491 29835
rect 29745 29801 29779 29835
rect 32045 29801 32079 29835
rect 8309 29733 8343 29767
rect 9137 29733 9171 29767
rect 11161 29733 11195 29767
rect 20729 29733 20763 29767
rect 33057 29733 33091 29767
rect 5181 29665 5215 29699
rect 6745 29665 6779 29699
rect 6929 29665 6963 29699
rect 20913 29665 20947 29699
rect 23765 29665 23799 29699
rect 23949 29665 23983 29699
rect 26065 29665 26099 29699
rect 28549 29665 28583 29699
rect 4169 29597 4203 29631
rect 4353 29597 4387 29631
rect 6653 29597 6687 29631
rect 6837 29597 6871 29631
rect 7481 29597 7515 29631
rect 8309 29597 8343 29631
rect 8493 29597 8527 29631
rect 9321 29597 9355 29631
rect 9413 29597 9447 29631
rect 10333 29597 10367 29631
rect 11253 29597 11287 29631
rect 13553 29597 13587 29631
rect 13737 29597 13771 29631
rect 14841 29597 14875 29631
rect 15117 29597 15151 29631
rect 15209 29597 15243 29631
rect 15485 29597 15519 29631
rect 15761 29597 15795 29631
rect 17693 29597 17727 29631
rect 17877 29597 17911 29631
rect 17969 29597 18003 29631
rect 18521 29597 18555 29631
rect 18705 29597 18739 29631
rect 19625 29597 19659 29631
rect 19717 29597 19751 29631
rect 19901 29597 19935 29631
rect 19993 29597 20027 29631
rect 21373 29597 21407 29631
rect 21557 29597 21591 29631
rect 23673 29597 23707 29631
rect 23857 29597 23891 29631
rect 25973 29597 26007 29631
rect 28273 29597 28307 29631
rect 29745 29597 29779 29631
rect 30021 29597 30055 29631
rect 32229 29597 32263 29631
rect 32413 29597 32447 29631
rect 32505 29597 32539 29631
rect 33149 29597 33183 29631
rect 33241 29597 33275 29631
rect 4445 29529 4479 29563
rect 6009 29529 6043 29563
rect 9137 29529 9171 29563
rect 14381 29529 14415 29563
rect 20453 29529 20487 29563
rect 21465 29529 21499 29563
rect 24593 29529 24627 29563
rect 32965 29529 32999 29563
rect 13737 29461 13771 29495
rect 19441 29461 19475 29495
rect 23489 29461 23523 29495
rect 24793 29461 24827 29495
rect 26341 29461 26375 29495
rect 28089 29461 28123 29495
rect 29929 29461 29963 29495
rect 6561 29257 6595 29291
rect 8401 29257 8435 29291
rect 18797 29257 18831 29291
rect 20085 29257 20119 29291
rect 23765 29257 23799 29291
rect 23949 29257 23983 29291
rect 25789 29257 25823 29291
rect 28089 29257 28123 29291
rect 25605 29189 25639 29223
rect 4997 29121 5031 29155
rect 5457 29121 5491 29155
rect 6837 29121 6871 29155
rect 6929 29121 6963 29155
rect 8217 29121 8251 29155
rect 14105 29121 14139 29155
rect 14197 29121 14231 29155
rect 14381 29121 14415 29155
rect 18981 29121 19015 29155
rect 19165 29121 19199 29155
rect 20269 29121 20303 29155
rect 20361 29121 20395 29155
rect 20545 29121 20579 29155
rect 20729 29121 20763 29155
rect 24777 29121 24811 29155
rect 24869 29121 24903 29155
rect 25053 29121 25087 29155
rect 25881 29121 25915 29155
rect 27813 29121 27847 29155
rect 28733 29121 28767 29155
rect 6745 29053 6779 29087
rect 7021 29053 7055 29087
rect 8033 29053 8067 29087
rect 8953 29053 8987 29087
rect 9229 29053 9263 29087
rect 19073 29053 19107 29087
rect 19257 29053 19291 29087
rect 22477 29053 22511 29087
rect 23397 29053 23431 29087
rect 23581 29053 23615 29087
rect 23673 29053 23707 29087
rect 24041 29053 24075 29087
rect 24593 29053 24627 29087
rect 27629 29053 27663 29087
rect 28181 29053 28215 29087
rect 29285 29053 29319 29087
rect 5365 28985 5399 29019
rect 13921 28985 13955 29019
rect 14289 28985 14323 29019
rect 20453 28985 20487 29019
rect 22845 28985 22879 29019
rect 24961 28985 24995 29019
rect 25605 28985 25639 29019
rect 10517 28917 10551 28951
rect 22937 28917 22971 28951
rect 9229 28713 9263 28747
rect 10333 28713 10367 28747
rect 14933 28713 14967 28747
rect 18797 28713 18831 28747
rect 19901 28713 19935 28747
rect 20085 28713 20119 28747
rect 23949 28713 23983 28747
rect 29929 28713 29963 28747
rect 28273 28645 28307 28679
rect 30113 28645 30147 28679
rect 33517 28645 33551 28679
rect 5549 28577 5583 28611
rect 6101 28577 6135 28611
rect 10701 28577 10735 28611
rect 24593 28577 24627 28611
rect 32965 28577 32999 28611
rect 5733 28509 5767 28543
rect 9413 28509 9447 28543
rect 9597 28509 9631 28543
rect 9715 28509 9749 28543
rect 9873 28509 9907 28543
rect 10517 28509 10551 28543
rect 10609 28509 10643 28543
rect 10793 28509 10827 28543
rect 14841 28509 14875 28543
rect 18705 28509 18739 28543
rect 19533 28509 19567 28543
rect 22753 28509 22787 28543
rect 23857 28509 23891 28543
rect 24777 28509 24811 28543
rect 28641 28509 28675 28543
rect 33149 28509 33183 28543
rect 33517 28509 33551 28543
rect 33885 28509 33919 28543
rect 9505 28441 9539 28475
rect 19901 28441 19935 28475
rect 23305 28441 23339 28475
rect 24961 28441 24995 28475
rect 28457 28441 28491 28475
rect 29745 28441 29779 28475
rect 5733 28373 5767 28407
rect 28549 28373 28583 28407
rect 28825 28373 28859 28407
rect 29945 28373 29979 28407
rect 5289 28169 5323 28203
rect 9321 28169 9355 28203
rect 24777 28169 24811 28203
rect 29101 28169 29135 28203
rect 29469 28169 29503 28203
rect 31217 28169 31251 28203
rect 5089 28101 5123 28135
rect 9689 28101 9723 28135
rect 16037 28101 16071 28135
rect 22569 28101 22603 28135
rect 24593 28101 24627 28135
rect 7573 28033 7607 28067
rect 9505 28033 9539 28067
rect 9781 28033 9815 28067
rect 15853 28033 15887 28067
rect 16129 28033 16163 28067
rect 16957 28033 16991 28067
rect 22201 28033 22235 28067
rect 22385 28033 22419 28067
rect 24409 28033 24443 28067
rect 28181 28033 28215 28067
rect 28457 28033 28491 28067
rect 28641 28033 28675 28067
rect 29285 28033 29319 28067
rect 29561 28033 29595 28067
rect 31401 28033 31435 28067
rect 31493 28033 31527 28067
rect 31677 28033 31711 28067
rect 32321 28033 32355 28067
rect 32505 28033 32539 28067
rect 33425 28033 33459 28067
rect 33609 28033 33643 28067
rect 34069 28033 34103 28067
rect 34345 28033 34379 28067
rect 34437 28033 34471 28067
rect 31585 27965 31619 27999
rect 33793 27965 33827 27999
rect 22201 27897 22235 27931
rect 5273 27829 5307 27863
rect 5457 27829 5491 27863
rect 7757 27829 7791 27863
rect 15669 27829 15703 27863
rect 17049 27829 17083 27863
rect 27997 27829 28031 27863
rect 32321 27829 32355 27863
rect 32137 27625 32171 27659
rect 4353 27557 4387 27591
rect 7205 27557 7239 27591
rect 19809 27557 19843 27591
rect 34069 27557 34103 27591
rect 4537 27489 4571 27523
rect 14841 27489 14875 27523
rect 25421 27489 25455 27523
rect 28457 27489 28491 27523
rect 31585 27489 31619 27523
rect 4261 27421 4295 27455
rect 7113 27421 7147 27455
rect 14473 27421 14507 27455
rect 14749 27421 14783 27455
rect 15945 27421 15979 27455
rect 16221 27421 16255 27455
rect 18245 27421 18279 27455
rect 18521 27421 18555 27455
rect 19441 27421 19475 27455
rect 19595 27421 19629 27455
rect 24593 27421 24627 27455
rect 24777 27421 24811 27455
rect 25329 27421 25363 27455
rect 25513 27421 25547 27455
rect 28181 27421 28215 27455
rect 28585 27421 28619 27455
rect 31217 27421 31251 27455
rect 32045 27421 32079 27455
rect 32689 27421 32723 27455
rect 32965 27421 32999 27455
rect 33333 27421 33367 27455
rect 34069 27421 34103 27455
rect 34161 27421 34195 27455
rect 28365 27353 28399 27387
rect 28457 27353 28491 27387
rect 31033 27353 31067 27387
rect 4537 27285 4571 27319
rect 17325 27285 17359 27319
rect 18061 27285 18095 27319
rect 18429 27285 18463 27319
rect 24777 27285 24811 27319
rect 18245 27081 18279 27115
rect 22017 27081 22051 27115
rect 22385 27081 22419 27115
rect 25605 27081 25639 27115
rect 32689 27081 32723 27115
rect 15853 27013 15887 27047
rect 16037 27013 16071 27047
rect 17132 27013 17166 27047
rect 26249 27013 26283 27047
rect 31769 27013 31803 27047
rect 3157 26945 3191 26979
rect 4629 26945 4663 26979
rect 4905 26945 4939 26979
rect 12449 26945 12483 26979
rect 13921 26945 13955 26979
rect 14289 26945 14323 26979
rect 16865 26945 16899 26979
rect 19441 26945 19475 26979
rect 22201 26945 22235 26979
rect 22477 26945 22511 26979
rect 24593 26945 24627 26979
rect 24777 26945 24811 26979
rect 25145 26945 25179 26979
rect 26065 26945 26099 26979
rect 27905 26945 27939 26979
rect 27997 26945 28031 26979
rect 28181 26945 28215 26979
rect 28273 26945 28307 26979
rect 31401 26945 31435 26979
rect 31677 26945 31711 26979
rect 32597 26945 32631 26979
rect 33149 26945 33183 26979
rect 3065 26877 3099 26911
rect 3525 26877 3559 26911
rect 4813 26877 4847 26911
rect 12265 26877 12299 26911
rect 13369 26877 13403 26911
rect 14013 26877 14047 26911
rect 14197 26877 14231 26911
rect 19717 26877 19751 26911
rect 25973 26877 26007 26911
rect 33425 26877 33459 26911
rect 4721 26809 4755 26843
rect 19257 26809 19291 26843
rect 25053 26809 25087 26843
rect 4445 26741 4479 26775
rect 12633 26741 12667 26775
rect 16037 26741 16071 26775
rect 16221 26741 16255 26775
rect 19625 26741 19659 26775
rect 27721 26741 27755 26775
rect 9137 26537 9171 26571
rect 26065 26537 26099 26571
rect 33885 26537 33919 26571
rect 5089 26469 5123 26503
rect 10057 26469 10091 26503
rect 20361 26469 20395 26503
rect 22201 26469 22235 26503
rect 32597 26469 32631 26503
rect 2789 26401 2823 26435
rect 4629 26401 4663 26435
rect 12173 26401 12207 26435
rect 14933 26401 14967 26435
rect 21465 26401 21499 26435
rect 23673 26401 23707 26435
rect 32965 26401 32999 26435
rect 2697 26333 2731 26367
rect 4169 26333 4203 26367
rect 4261 26333 4295 26367
rect 4537 26333 4571 26367
rect 5365 26333 5399 26367
rect 9321 26333 9355 26367
rect 9597 26333 9631 26367
rect 10333 26333 10367 26367
rect 12081 26333 12115 26367
rect 12357 26333 12391 26367
rect 12725 26333 12759 26367
rect 14381 26333 14415 26367
rect 16313 26333 16347 26367
rect 20545 26333 20579 26367
rect 21373 26333 21407 26367
rect 21557 26333 21591 26367
rect 22385 26333 22419 26367
rect 22477 26333 22511 26367
rect 22661 26333 22695 26367
rect 22753 26333 22787 26367
rect 23397 26333 23431 26367
rect 24869 26333 24903 26367
rect 25237 26333 25271 26367
rect 25329 26333 25363 26367
rect 26065 26333 26099 26367
rect 31493 26333 31527 26367
rect 31769 26333 31803 26367
rect 32873 26333 32907 26367
rect 33517 26333 33551 26367
rect 33701 26333 33735 26367
rect 3341 26265 3375 26299
rect 5089 26265 5123 26299
rect 5273 26265 5307 26299
rect 10057 26265 10091 26299
rect 31677 26265 31711 26299
rect 32321 26265 32355 26299
rect 3985 26197 4019 26231
rect 9505 26197 9539 26231
rect 10241 26197 10275 26231
rect 17601 26197 17635 26231
rect 31309 26197 31343 26231
rect 5181 25993 5215 26027
rect 12449 25993 12483 26027
rect 18429 25993 18463 26027
rect 4721 25925 4755 25959
rect 5457 25925 5491 25959
rect 5549 25925 5583 25959
rect 8953 25925 8987 25959
rect 16221 25925 16255 25959
rect 2421 25857 2455 25891
rect 2605 25857 2639 25891
rect 3341 25857 3375 25891
rect 5365 25857 5399 25891
rect 5733 25857 5767 25891
rect 5825 25857 5859 25891
rect 9873 25857 9907 25891
rect 10057 25857 10091 25891
rect 10149 25857 10183 25891
rect 10609 25857 10643 25891
rect 10793 25857 10827 25891
rect 12081 25857 12115 25891
rect 12265 25857 12299 25891
rect 12541 25857 12575 25891
rect 15669 25857 15703 25891
rect 17316 25857 17350 25891
rect 23857 25857 23891 25891
rect 28641 25857 28675 25891
rect 31033 25857 31067 25891
rect 31217 25857 31251 25891
rect 31309 25857 31343 25891
rect 3065 25789 3099 25823
rect 17049 25789 17083 25823
rect 24041 25789 24075 25823
rect 9321 25721 9355 25755
rect 9965 25721 9999 25755
rect 2513 25653 2547 25687
rect 9413 25653 9447 25687
rect 10701 25653 10735 25687
rect 29929 25653 29963 25687
rect 30849 25653 30883 25687
rect 3249 25449 3283 25483
rect 5365 25449 5399 25483
rect 8401 25449 8435 25483
rect 10701 25449 10735 25483
rect 16957 25449 16991 25483
rect 17877 25449 17911 25483
rect 31953 25449 31987 25483
rect 3985 25381 4019 25415
rect 7573 25381 7607 25415
rect 10885 25381 10919 25415
rect 13461 25381 13495 25415
rect 8585 25313 8619 25347
rect 9321 25313 9355 25347
rect 9689 25313 9723 25347
rect 9781 25313 9815 25347
rect 20453 25313 20487 25347
rect 3249 25245 3283 25279
rect 3433 25245 3467 25279
rect 4169 25245 4203 25279
rect 4261 25245 4295 25279
rect 5089 25245 5123 25279
rect 5181 25245 5215 25279
rect 7757 25245 7791 25279
rect 7849 25245 7883 25279
rect 8309 25245 8343 25279
rect 9413 25245 9447 25279
rect 10333 25245 10367 25279
rect 10609 25245 10643 25279
rect 11713 25245 11747 25279
rect 12357 25245 12391 25279
rect 12541 25245 12575 25279
rect 13185 25245 13219 25279
rect 13461 25245 13495 25279
rect 18061 25245 18095 25279
rect 18337 25245 18371 25279
rect 19441 25245 19475 25279
rect 19625 25245 19659 25279
rect 20085 25245 20119 25279
rect 20361 25245 20395 25279
rect 23213 25245 23247 25279
rect 27353 25245 27387 25279
rect 30573 25245 30607 25279
rect 30840 25245 30874 25279
rect 32505 25245 32539 25279
rect 3985 25177 4019 25211
rect 7573 25177 7607 25211
rect 8585 25177 8619 25211
rect 11805 25177 11839 25211
rect 15669 25177 15703 25211
rect 18245 25177 18279 25211
rect 23581 25177 23615 25211
rect 27620 25177 27654 25211
rect 9137 25109 9171 25143
rect 9505 25109 9539 25143
rect 12633 25109 12667 25143
rect 19625 25109 19659 25143
rect 28733 25109 28767 25143
rect 32597 25109 32631 25143
rect 9873 24905 9907 24939
rect 10517 24905 10551 24939
rect 24777 24905 24811 24939
rect 13277 24837 13311 24871
rect 7849 24769 7883 24803
rect 8116 24769 8150 24803
rect 9781 24769 9815 24803
rect 9965 24769 9999 24803
rect 10425 24769 10459 24803
rect 12265 24769 12299 24803
rect 12357 24769 12391 24803
rect 12909 24769 12943 24803
rect 13185 24769 13219 24803
rect 16865 24769 16899 24803
rect 17049 24769 17083 24803
rect 17233 24769 17267 24803
rect 17325 24769 17359 24803
rect 22661 24769 22695 24803
rect 22845 24769 22879 24803
rect 22937 24769 22971 24803
rect 23397 24769 23431 24803
rect 29745 24769 29779 24803
rect 32505 24769 32539 24803
rect 32689 24769 32723 24803
rect 32781 24769 32815 24803
rect 23673 24701 23707 24735
rect 27629 24701 27663 24735
rect 27905 24701 27939 24735
rect 32321 24701 32355 24735
rect 31033 24633 31067 24667
rect 9229 24565 9263 24599
rect 22477 24565 22511 24599
rect 29193 24565 29227 24599
rect 16865 24361 16899 24395
rect 24041 24361 24075 24395
rect 27261 24361 27295 24395
rect 31401 24361 31435 24395
rect 24961 24225 24995 24259
rect 26433 24225 26467 24259
rect 15485 24157 15519 24191
rect 15752 24157 15786 24191
rect 22661 24157 22695 24191
rect 24685 24157 24719 24191
rect 25881 24157 25915 24191
rect 27445 24157 27479 24191
rect 27721 24157 27755 24191
rect 30021 24157 30055 24191
rect 21833 24089 21867 24123
rect 22201 24089 22235 24123
rect 22906 24089 22940 24123
rect 27629 24089 27663 24123
rect 30288 24089 30322 24123
rect 22477 23817 22511 23851
rect 22845 23817 22879 23851
rect 27813 23817 27847 23851
rect 25145 23749 25179 23783
rect 12725 23681 12759 23715
rect 19717 23681 19751 23715
rect 20361 23681 20395 23715
rect 22661 23681 22695 23715
rect 22934 23681 22968 23715
rect 23397 23681 23431 23715
rect 25697 23681 25731 23715
rect 27537 23681 27571 23715
rect 27721 23681 27755 23715
rect 34805 23681 34839 23715
rect 36001 23681 36035 23715
rect 36093 23681 36127 23715
rect 13001 23613 13035 23647
rect 20453 23613 20487 23647
rect 25973 23613 26007 23647
rect 34529 23613 34563 23647
rect 35357 23613 35391 23647
rect 14473 23477 14507 23511
rect 19809 23477 19843 23511
rect 36277 23477 36311 23511
rect 7389 23273 7423 23307
rect 14381 23273 14415 23307
rect 19441 23273 19475 23307
rect 23213 23273 23247 23307
rect 27813 23273 27847 23307
rect 32505 23273 32539 23307
rect 3985 23205 4019 23239
rect 25973 23205 26007 23239
rect 13461 23137 13495 23171
rect 19717 23137 19751 23171
rect 20085 23137 20119 23171
rect 20821 23137 20855 23171
rect 20913 23137 20947 23171
rect 35817 23137 35851 23171
rect 36461 23137 36495 23171
rect 4537 23069 4571 23103
rect 12541 23069 12575 23103
rect 13001 23069 13035 23103
rect 13185 23069 13219 23103
rect 13553 23069 13587 23103
rect 14289 23069 14323 23103
rect 14473 23069 14507 23103
rect 19625 23069 19659 23103
rect 20729 23069 20763 23103
rect 21005 23069 21039 23103
rect 23397 23069 23431 23103
rect 23581 23069 23615 23103
rect 23673 23069 23707 23103
rect 24593 23069 24627 23103
rect 31217 23069 31251 23103
rect 35909 23069 35943 23103
rect 4169 23001 4203 23035
rect 7665 23001 7699 23035
rect 7941 23001 7975 23035
rect 24860 23001 24894 23035
rect 26525 23001 26559 23035
rect 4261 22933 4295 22967
rect 4353 22933 4387 22967
rect 7849 22933 7883 22967
rect 19809 22933 19843 22967
rect 19993 22933 20027 22967
rect 20545 22933 20579 22967
rect 4997 22729 5031 22763
rect 8677 22729 8711 22763
rect 17785 22729 17819 22763
rect 25881 22729 25915 22763
rect 26249 22729 26283 22763
rect 29837 22729 29871 22763
rect 36369 22729 36403 22763
rect 3525 22661 3559 22695
rect 8033 22661 8067 22695
rect 14749 22661 14783 22695
rect 17601 22661 17635 22695
rect 19349 22661 19383 22695
rect 19441 22661 19475 22695
rect 20361 22661 20395 22695
rect 6561 22593 6595 22627
rect 7021 22593 7055 22627
rect 7389 22593 7423 22627
rect 8180 22593 8214 22627
rect 9689 22593 9723 22627
rect 11805 22593 11839 22627
rect 11897 22593 11931 22627
rect 13001 22593 13035 22627
rect 18521 22593 18555 22627
rect 19073 22593 19107 22627
rect 20177 22593 20211 22627
rect 20453 22593 20487 22627
rect 23673 22593 23707 22627
rect 26065 22593 26099 22627
rect 26341 22593 26375 22627
rect 27813 22593 27847 22627
rect 28089 22593 28123 22627
rect 28181 22593 28215 22627
rect 29929 22593 29963 22627
rect 30481 22593 30515 22627
rect 33333 22593 33367 22627
rect 33425 22593 33459 22627
rect 35541 22593 35575 22627
rect 35633 22593 35667 22627
rect 35725 22593 35759 22627
rect 36277 22593 36311 22627
rect 36461 22593 36495 22627
rect 3249 22525 3283 22559
rect 7481 22525 7515 22559
rect 8401 22525 8435 22559
rect 12081 22525 12115 22559
rect 18981 22525 19015 22559
rect 27721 22525 27755 22559
rect 30665 22525 30699 22559
rect 35449 22525 35483 22559
rect 33609 22457 33643 22491
rect 8309 22389 8343 22423
rect 9781 22389 9815 22423
rect 17785 22389 17819 22423
rect 17969 22389 18003 22423
rect 18797 22389 18831 22423
rect 19993 22389 20027 22423
rect 24961 22389 24995 22423
rect 27537 22389 27571 22423
rect 35265 22389 35299 22423
rect 3249 22185 3283 22219
rect 3433 22185 3467 22219
rect 7205 22185 7239 22219
rect 26341 22185 26375 22219
rect 27813 22185 27847 22219
rect 30205 22185 30239 22219
rect 33793 22185 33827 22219
rect 37105 22185 37139 22219
rect 6561 22117 6595 22151
rect 24869 22117 24903 22151
rect 34897 22117 34931 22151
rect 4353 22049 4387 22083
rect 9597 22049 9631 22083
rect 10701 22049 10735 22083
rect 10977 22049 11011 22083
rect 27721 22049 27755 22083
rect 32965 22049 32999 22083
rect 36001 22049 36035 22083
rect 2421 21981 2455 22015
rect 4077 21981 4111 22015
rect 4169 21981 4203 22015
rect 7113 21981 7147 22015
rect 7297 21981 7331 22015
rect 8309 21981 8343 22015
rect 8493 21981 8527 22015
rect 9321 21981 9355 22015
rect 9413 21981 9447 22015
rect 9689 21981 9723 22015
rect 14381 21981 14415 22015
rect 15853 21981 15887 22015
rect 16037 21981 16071 22015
rect 16221 21981 16255 22015
rect 16865 21981 16899 22015
rect 19441 21981 19475 22015
rect 19708 21981 19742 22015
rect 24593 21981 24627 22015
rect 24777 21981 24811 22015
rect 26249 21981 26283 22015
rect 26433 21981 26467 22015
rect 27629 21981 27663 22015
rect 29929 21981 29963 22015
rect 30757 21981 30791 22015
rect 30941 21981 30975 22015
rect 32505 21981 32539 22015
rect 33333 21981 33367 22015
rect 35173 21981 35207 22015
rect 36185 21981 36219 22015
rect 36369 21981 36403 22015
rect 37013 21981 37047 22015
rect 37841 21981 37875 22015
rect 38025 21981 38059 22015
rect 3065 21913 3099 21947
rect 6193 21913 6227 21947
rect 8401 21913 8435 21947
rect 14841 21913 14875 21947
rect 16129 21913 16163 21947
rect 17110 21913 17144 21947
rect 30113 21913 30147 21947
rect 30849 21913 30883 21947
rect 34897 21913 34931 21947
rect 36829 21913 36863 21947
rect 37933 21913 37967 21947
rect 2513 21845 2547 21879
rect 3275 21845 3309 21879
rect 6653 21845 6687 21879
rect 9137 21845 9171 21879
rect 12449 21845 12483 21879
rect 16405 21845 16439 21879
rect 18245 21845 18279 21879
rect 20821 21845 20855 21879
rect 27997 21845 28031 21879
rect 35081 21845 35115 21879
rect 6929 21641 6963 21675
rect 7573 21641 7607 21675
rect 9689 21641 9723 21675
rect 11069 21641 11103 21675
rect 24501 21641 24535 21675
rect 34621 21641 34655 21675
rect 4537 21573 4571 21607
rect 16221 21573 16255 21607
rect 18245 21573 18279 21607
rect 23388 21573 23422 21607
rect 36921 21573 36955 21607
rect 1869 21505 1903 21539
rect 4261 21505 4295 21539
rect 4445 21505 4479 21539
rect 6745 21505 6779 21539
rect 7481 21505 7515 21539
rect 7665 21505 7699 21539
rect 9229 21505 9263 21539
rect 9505 21505 9539 21539
rect 10885 21505 10919 21539
rect 10977 21505 11011 21539
rect 12081 21505 12115 21539
rect 13001 21505 13035 21539
rect 16037 21505 16071 21539
rect 16313 21505 16347 21539
rect 21097 21505 21131 21539
rect 21281 21505 21315 21539
rect 21373 21505 21407 21539
rect 27997 21505 28031 21539
rect 28181 21505 28215 21539
rect 33241 21505 33275 21539
rect 34621 21505 34655 21539
rect 2145 21437 2179 21471
rect 6561 21437 6595 21471
rect 9413 21437 9447 21471
rect 23121 21437 23155 21471
rect 28365 21437 28399 21471
rect 33333 21437 33367 21471
rect 34759 21437 34793 21471
rect 34989 21437 35023 21471
rect 36093 21437 36127 21471
rect 3617 21301 3651 21335
rect 9229 21301 9263 21335
rect 12173 21301 12207 21335
rect 14289 21301 14323 21335
rect 15853 21301 15887 21335
rect 19533 21301 19567 21335
rect 20913 21301 20947 21335
rect 33517 21301 33551 21335
rect 5549 21097 5583 21131
rect 10977 21097 11011 21131
rect 27353 21097 27387 21131
rect 36001 21097 36035 21131
rect 5733 21029 5767 21063
rect 35357 21029 35391 21063
rect 3065 20961 3099 20995
rect 12265 20961 12299 20995
rect 14933 20961 14967 20995
rect 17417 20961 17451 20995
rect 22569 20961 22603 20995
rect 35449 20961 35483 20995
rect 36645 20961 36679 20995
rect 2789 20893 2823 20927
rect 3249 20893 3283 20927
rect 7389 20893 7423 20927
rect 7573 20893 7607 20927
rect 9137 20893 9171 20927
rect 9597 20893 9631 20927
rect 9781 20893 9815 20927
rect 10885 20893 10919 20927
rect 11989 20893 12023 20927
rect 14381 20893 14415 20927
rect 20821 20893 20855 20927
rect 26065 20893 26099 20927
rect 29745 20893 29779 20927
rect 29929 20893 29963 20927
rect 34897 20893 34931 20927
rect 35081 20893 35115 20927
rect 36165 20893 36199 20927
rect 36277 20893 36311 20927
rect 5365 20825 5399 20859
rect 5581 20825 5615 20859
rect 7481 20825 7515 20859
rect 15669 20825 15703 20859
rect 36553 20825 36587 20859
rect 10425 20757 10459 20791
rect 29837 20757 29871 20791
rect 2789 20553 2823 20587
rect 6938 20553 6972 20587
rect 9229 20553 9263 20587
rect 16865 20553 16899 20587
rect 17233 20553 17267 20587
rect 19533 20553 19567 20587
rect 21097 20553 21131 20587
rect 6561 20485 6595 20519
rect 13001 20485 13035 20519
rect 18245 20485 18279 20519
rect 20821 20485 20855 20519
rect 26249 20485 26283 20519
rect 2697 20417 2731 20451
rect 7205 20417 7239 20451
rect 7665 20417 7699 20451
rect 9045 20417 9079 20451
rect 11897 20417 11931 20451
rect 15393 20417 15427 20451
rect 15577 20417 15611 20451
rect 15669 20417 15703 20451
rect 17049 20417 17083 20451
rect 17325 20417 17359 20451
rect 20453 20417 20487 20451
rect 20546 20417 20580 20451
rect 20729 20417 20763 20451
rect 20918 20417 20952 20451
rect 23765 20417 23799 20451
rect 26065 20417 26099 20451
rect 26341 20417 26375 20451
rect 30573 20417 30607 20451
rect 30757 20417 30791 20451
rect 30849 20417 30883 20451
rect 9505 20349 9539 20383
rect 9597 20349 9631 20383
rect 12173 20349 12207 20383
rect 14749 20349 14783 20383
rect 24041 20349 24075 20383
rect 38117 20349 38151 20383
rect 6929 20213 6963 20247
rect 7757 20213 7791 20247
rect 15209 20213 15243 20247
rect 25881 20213 25915 20247
rect 30389 20213 30423 20247
rect 17233 20009 17267 20043
rect 20821 20009 20855 20043
rect 21925 20009 21959 20043
rect 27537 20009 27571 20043
rect 28365 20009 28399 20043
rect 28641 20009 28675 20043
rect 31125 20009 31159 20043
rect 34989 20009 35023 20043
rect 36737 20009 36771 20043
rect 13737 19941 13771 19975
rect 19441 19873 19475 19907
rect 30021 19873 30055 19907
rect 36093 19873 36127 19907
rect 12357 19805 12391 19839
rect 14473 19805 14507 19839
rect 14657 19805 14691 19839
rect 14749 19805 14783 19839
rect 15853 19805 15887 19839
rect 16120 19805 16154 19839
rect 19708 19805 19742 19839
rect 21281 19805 21315 19839
rect 21374 19805 21408 19839
rect 21649 19805 21683 19839
rect 21787 19805 21821 19839
rect 23673 19805 23707 19839
rect 24777 19805 24811 19839
rect 24870 19805 24904 19839
rect 25053 19805 25087 19839
rect 25242 19805 25276 19839
rect 26065 19805 26099 19839
rect 28273 19805 28307 19839
rect 28457 19805 28491 19839
rect 29745 19805 29779 19839
rect 32045 19805 32079 19839
rect 32321 19805 32355 19839
rect 34989 19805 35023 19839
rect 35081 19805 35115 19839
rect 35725 19805 35759 19839
rect 36001 19805 36035 19839
rect 36553 19805 36587 19839
rect 36707 19805 36741 19839
rect 12624 19737 12658 19771
rect 14289 19737 14323 19771
rect 21557 19737 21591 19771
rect 25145 19737 25179 19771
rect 23765 19669 23799 19703
rect 25421 19669 25455 19703
rect 31861 19669 31895 19703
rect 32229 19669 32263 19703
rect 7665 19465 7699 19499
rect 14013 19465 14047 19499
rect 18337 19465 18371 19499
rect 23857 19465 23891 19499
rect 26617 19465 26651 19499
rect 36645 19465 36679 19499
rect 7481 19397 7515 19431
rect 25504 19397 25538 19431
rect 27537 19397 27571 19431
rect 31309 19397 31343 19431
rect 4813 19329 4847 19363
rect 5089 19329 5123 19363
rect 6745 19329 6779 19363
rect 7941 19329 7975 19363
rect 12725 19329 12759 19363
rect 17969 19329 18003 19363
rect 22477 19329 22511 19363
rect 22744 19329 22778 19363
rect 27353 19329 27387 19363
rect 27629 19329 27663 19363
rect 35541 19329 35575 19363
rect 35725 19329 35759 19363
rect 36185 19329 36219 19363
rect 36461 19329 36495 19363
rect 7021 19261 7055 19295
rect 18061 19261 18095 19295
rect 25237 19261 25271 19295
rect 29653 19261 29687 19295
rect 29929 19261 29963 19295
rect 36277 19261 36311 19295
rect 35541 19193 35575 19227
rect 4905 19125 4939 19159
rect 6561 19125 6595 19159
rect 6929 19125 6963 19159
rect 7665 19125 7699 19159
rect 18153 19125 18187 19159
rect 27169 19125 27203 19159
rect 6929 18921 6963 18955
rect 13277 18921 13311 18955
rect 13461 18921 13495 18955
rect 22201 18921 22235 18955
rect 23213 18921 23247 18955
rect 26893 18921 26927 18955
rect 28457 18921 28491 18955
rect 16773 18853 16807 18887
rect 36093 18853 36127 18887
rect 4261 18785 4295 18819
rect 18889 18785 18923 18819
rect 28633 18785 28667 18819
rect 28917 18785 28951 18819
rect 30389 18785 30423 18819
rect 32965 18785 32999 18819
rect 2145 18717 2179 18751
rect 2329 18717 2363 18751
rect 2789 18717 2823 18751
rect 2973 18717 3007 18751
rect 3985 18717 4019 18751
rect 10057 18717 10091 18751
rect 16589 18717 16623 18751
rect 16773 18717 16807 18751
rect 17417 18717 17451 18751
rect 17601 18717 17635 18751
rect 18521 18717 18555 18751
rect 23397 18717 23431 18751
rect 23673 18717 23707 18751
rect 25513 18717 25547 18751
rect 28711 18717 28745 18751
rect 28826 18717 28860 18751
rect 30113 18717 30147 18751
rect 35725 18717 35759 18751
rect 35909 18717 35943 18751
rect 36185 18717 36219 18751
rect 36461 18717 36495 18751
rect 6745 18649 6779 18683
rect 6929 18649 6963 18683
rect 13093 18649 13127 18683
rect 18337 18649 18371 18683
rect 22017 18649 22051 18683
rect 22201 18649 22235 18683
rect 23581 18649 23615 18683
rect 25780 18649 25814 18683
rect 29929 18649 29963 18683
rect 33517 18649 33551 18683
rect 2237 18581 2271 18615
rect 2973 18581 3007 18615
rect 5733 18581 5767 18615
rect 7113 18581 7147 18615
rect 10149 18581 10183 18615
rect 13277 18581 13311 18615
rect 17417 18581 17451 18615
rect 22385 18581 22419 18615
rect 3617 18377 3651 18411
rect 4077 18377 4111 18411
rect 14289 18377 14323 18411
rect 17233 18377 17267 18411
rect 26065 18377 26099 18411
rect 29929 18377 29963 18411
rect 35817 18377 35851 18411
rect 36185 18377 36219 18411
rect 2145 18309 2179 18343
rect 13176 18309 13210 18343
rect 18337 18309 18371 18343
rect 18889 18309 18923 18343
rect 22569 18309 22603 18343
rect 35633 18309 35667 18343
rect 35909 18309 35943 18343
rect 4261 18241 4295 18275
rect 7849 18241 7883 18275
rect 10324 18241 10358 18275
rect 10425 18241 10459 18275
rect 10609 18241 10643 18275
rect 12909 18241 12943 18275
rect 17233 18241 17267 18275
rect 17601 18241 17635 18275
rect 18521 18241 18555 18275
rect 19349 18241 19383 18275
rect 19533 18241 19567 18275
rect 24777 18241 24811 18275
rect 28641 18241 28675 18275
rect 30849 18241 30883 18275
rect 31033 18241 31067 18275
rect 32781 18241 32815 18275
rect 33149 18241 33183 18275
rect 33333 18241 33367 18275
rect 33701 18241 33735 18275
rect 34529 18241 34563 18275
rect 34989 18241 35023 18275
rect 36001 18241 36035 18275
rect 1869 18173 1903 18207
rect 4537 18173 4571 18207
rect 11069 18173 11103 18207
rect 19901 18173 19935 18207
rect 32965 18173 32999 18207
rect 34805 18173 34839 18207
rect 4445 18105 4479 18139
rect 9137 18037 9171 18071
rect 23857 18037 23891 18071
rect 30941 18037 30975 18071
rect 2789 17833 2823 17867
rect 22109 17833 22143 17867
rect 24869 17833 24903 17867
rect 28273 17833 28307 17867
rect 33425 17833 33459 17867
rect 28457 17697 28491 17731
rect 28549 17697 28583 17731
rect 33609 17697 33643 17731
rect 2789 17629 2823 17663
rect 2973 17629 3007 17663
rect 8493 17629 8527 17663
rect 9137 17629 9171 17663
rect 12357 17629 12391 17663
rect 15393 17629 15427 17663
rect 18153 17629 18187 17663
rect 18705 17629 18739 17663
rect 23213 17629 23247 17663
rect 23489 17629 23523 17663
rect 25145 17629 25179 17663
rect 25605 17629 25639 17663
rect 28641 17629 28675 17663
rect 28733 17629 28767 17663
rect 29745 17629 29779 17663
rect 32321 17629 32355 17663
rect 32597 17629 32631 17663
rect 33793 17629 33827 17663
rect 34161 17629 34195 17663
rect 34345 17629 34379 17663
rect 8217 17561 8251 17595
rect 9413 17561 9447 17595
rect 12624 17561 12658 17595
rect 18889 17561 18923 17595
rect 20821 17561 20855 17595
rect 24685 17561 24719 17595
rect 24869 17561 24903 17595
rect 32689 17561 32723 17595
rect 7923 17493 7957 17527
rect 8401 17493 8435 17527
rect 10885 17493 10919 17527
rect 13737 17493 13771 17527
rect 16681 17493 16715 17527
rect 23029 17493 23063 17527
rect 23397 17493 23431 17527
rect 26893 17493 26927 17527
rect 31033 17493 31067 17527
rect 10057 17289 10091 17323
rect 18889 17289 18923 17323
rect 21373 17289 21407 17323
rect 32505 17289 32539 17323
rect 33149 17289 33183 17323
rect 7389 17221 7423 17255
rect 18613 17221 18647 17255
rect 32597 17221 32631 17255
rect 5365 17153 5399 17187
rect 5549 17153 5583 17187
rect 6745 17153 6779 17187
rect 10701 17153 10735 17187
rect 10885 17153 10919 17187
rect 12992 17153 13026 17187
rect 14657 17153 14691 17187
rect 16865 17153 16899 17187
rect 17509 17153 17543 17187
rect 18245 17153 18279 17187
rect 18338 17153 18372 17187
rect 18521 17153 18555 17187
rect 18710 17153 18744 17187
rect 21189 17153 21223 17187
rect 21465 17153 21499 17187
rect 22017 17153 22051 17187
rect 22284 17153 22318 17187
rect 23857 17153 23891 17187
rect 24113 17153 24147 17187
rect 32413 17153 32447 17187
rect 32689 17153 32723 17187
rect 33333 17153 33367 17187
rect 33609 17153 33643 17187
rect 33793 17153 33827 17187
rect 5273 17085 5307 17119
rect 6009 17085 6043 17119
rect 10057 17085 10091 17119
rect 10149 17085 10183 17119
rect 12725 17085 12759 17119
rect 15025 17085 15059 17119
rect 10793 17017 10827 17051
rect 9597 16949 9631 16983
rect 14105 16949 14139 16983
rect 17325 16949 17359 16983
rect 21005 16949 21039 16983
rect 23397 16949 23431 16983
rect 25237 16949 25271 16983
rect 3249 16745 3283 16779
rect 13277 16745 13311 16779
rect 23397 16745 23431 16779
rect 33057 16745 33091 16779
rect 36185 16745 36219 16779
rect 36737 16745 36771 16779
rect 3433 16677 3467 16711
rect 5089 16609 5123 16643
rect 5365 16609 5399 16643
rect 21005 16609 21039 16643
rect 7389 16541 7423 16575
rect 13461 16541 13495 16575
rect 13737 16541 13771 16575
rect 17233 16541 17267 16575
rect 17417 16541 17451 16575
rect 17693 16541 17727 16575
rect 21261 16541 21295 16575
rect 23581 16541 23615 16575
rect 23857 16541 23891 16575
rect 25973 16541 26007 16575
rect 26249 16541 26283 16575
rect 29745 16541 29779 16575
rect 33241 16541 33275 16575
rect 33517 16541 33551 16575
rect 36093 16541 36127 16575
rect 36921 16541 36955 16575
rect 37105 16541 37139 16575
rect 37197 16541 37231 16575
rect 3065 16473 3099 16507
rect 3281 16473 3315 16507
rect 7665 16473 7699 16507
rect 23765 16473 23799 16507
rect 29990 16473 30024 16507
rect 35909 16473 35943 16507
rect 6837 16405 6871 16439
rect 13645 16405 13679 16439
rect 22385 16405 22419 16439
rect 25789 16405 25823 16439
rect 26157 16405 26191 16439
rect 31125 16405 31159 16439
rect 33425 16405 33459 16439
rect 13369 16201 13403 16235
rect 15209 16201 15243 16235
rect 20821 16201 20855 16235
rect 28549 16201 28583 16235
rect 35909 16201 35943 16235
rect 36829 16201 36863 16235
rect 37841 16201 37875 16235
rect 6009 16133 6043 16167
rect 6837 16133 6871 16167
rect 14841 16133 14875 16167
rect 25504 16133 25538 16167
rect 28917 16133 28951 16167
rect 5641 16065 5675 16099
rect 5917 16065 5951 16099
rect 6561 16065 6595 16099
rect 9229 16065 9263 16099
rect 13553 16065 13587 16099
rect 13737 16065 13771 16099
rect 13829 16065 13863 16099
rect 14565 16065 14599 16099
rect 14658 16065 14692 16099
rect 14933 16065 14967 16099
rect 15071 16065 15105 16099
rect 16865 16065 16899 16099
rect 17233 16065 17267 16099
rect 17417 16065 17451 16099
rect 18061 16065 18095 16099
rect 18429 16065 18463 16099
rect 18613 16065 18647 16099
rect 21005 16065 21039 16099
rect 21097 16065 21131 16099
rect 21281 16065 21315 16099
rect 21373 16065 21407 16099
rect 28733 16065 28767 16099
rect 29009 16065 29043 16099
rect 29736 16065 29770 16099
rect 35817 16065 35851 16099
rect 36001 16065 36035 16099
rect 36645 16065 36679 16099
rect 37657 16065 37691 16099
rect 9505 15997 9539 16031
rect 25237 15997 25271 16031
rect 29469 15997 29503 16031
rect 36461 15997 36495 16031
rect 37473 15997 37507 16031
rect 8309 15861 8343 15895
rect 10977 15861 11011 15895
rect 26617 15861 26651 15895
rect 30849 15861 30883 15895
rect 30665 15657 30699 15691
rect 34253 15657 34287 15691
rect 35265 15657 35299 15691
rect 37381 15657 37415 15691
rect 36829 15589 36863 15623
rect 7205 15521 7239 15555
rect 9965 15521 9999 15555
rect 12173 15521 12207 15555
rect 16681 15521 16715 15555
rect 18153 15521 18187 15555
rect 25789 15521 25823 15555
rect 29929 15521 29963 15555
rect 36369 15521 36403 15555
rect 6837 15453 6871 15487
rect 7113 15453 7147 15487
rect 9689 15453 9723 15487
rect 9781 15453 9815 15487
rect 10425 15453 10459 15487
rect 16405 15453 16439 15487
rect 17049 15453 17083 15487
rect 17785 15453 17819 15487
rect 18061 15453 18095 15487
rect 19441 15453 19475 15487
rect 19625 15453 19659 15487
rect 24777 15453 24811 15487
rect 25053 15453 25087 15487
rect 25145 15453 25179 15487
rect 29745 15453 29779 15487
rect 30849 15453 30883 15487
rect 31125 15453 31159 15487
rect 34161 15453 34195 15487
rect 34345 15453 34379 15487
rect 35081 15453 35115 15487
rect 36553 15453 36587 15487
rect 36921 15453 36955 15487
rect 37381 15453 37415 15487
rect 37565 15453 37599 15487
rect 19809 15385 19843 15419
rect 24961 15385 24995 15419
rect 26056 15385 26090 15419
rect 34897 15385 34931 15419
rect 25329 15317 25363 15351
rect 27169 15317 27203 15351
rect 31033 15317 31067 15351
rect 2605 15113 2639 15147
rect 2973 15113 3007 15147
rect 3157 15113 3191 15147
rect 21281 15113 21315 15147
rect 26157 15113 26191 15147
rect 26525 15113 26559 15147
rect 28181 15113 28215 15147
rect 33517 15113 33551 15147
rect 34897 15113 34931 15147
rect 34989 15113 35023 15147
rect 36829 15113 36863 15147
rect 20913 15045 20947 15079
rect 21005 15045 21039 15079
rect 30849 15045 30883 15079
rect 35173 15045 35207 15079
rect 36461 15045 36495 15079
rect 36661 15045 36695 15079
rect 3249 14977 3283 15011
rect 3709 14977 3743 15011
rect 3893 14977 3927 15011
rect 13921 14977 13955 15011
rect 16865 14977 16899 15011
rect 17509 14977 17543 15011
rect 18797 14977 18831 15011
rect 19257 14977 19291 15011
rect 20644 14977 20678 15011
rect 20730 14977 20764 15011
rect 21143 14977 21177 15011
rect 26341 14977 26375 15011
rect 26617 14977 26651 15011
rect 28457 14977 28491 15011
rect 28641 14977 28675 15011
rect 30573 14977 30607 15011
rect 30757 14977 30791 15011
rect 30941 14977 30975 15011
rect 32689 14977 32723 15011
rect 33333 14977 33367 15011
rect 33609 14977 33643 15011
rect 33701 14977 33735 15011
rect 34805 14977 34839 15011
rect 35817 14977 35851 15011
rect 2789 14909 2823 14943
rect 2881 14909 2915 14943
rect 14197 14909 14231 14943
rect 17601 14909 17635 14943
rect 19533 14909 19567 14943
rect 28365 14909 28399 14943
rect 28549 14909 28583 14943
rect 34621 14909 34655 14943
rect 35633 14909 35667 14943
rect 32781 14841 32815 14875
rect 3801 14773 3835 14807
rect 31125 14773 31159 14807
rect 33885 14773 33919 14807
rect 36001 14773 36035 14807
rect 36645 14773 36679 14807
rect 20637 14569 20671 14603
rect 26893 14569 26927 14603
rect 34897 14569 34931 14603
rect 35909 14569 35943 14603
rect 3065 14433 3099 14467
rect 3157 14433 3191 14467
rect 17325 14433 17359 14467
rect 18889 14433 18923 14467
rect 23213 14433 23247 14467
rect 2145 14365 2179 14399
rect 2237 14365 2271 14399
rect 2973 14365 3007 14399
rect 3249 14365 3283 14399
rect 13461 14365 13495 14399
rect 13737 14365 13771 14399
rect 16037 14365 16071 14399
rect 16221 14365 16255 14399
rect 16773 14365 16807 14399
rect 16957 14365 16991 14399
rect 18429 14365 18463 14399
rect 18613 14365 18647 14399
rect 20085 14365 20119 14399
rect 20269 14365 20303 14399
rect 20453 14365 20487 14399
rect 22937 14365 22971 14399
rect 26249 14365 26283 14399
rect 26342 14365 26376 14399
rect 26714 14365 26748 14399
rect 35173 14365 35207 14399
rect 35270 14365 35304 14399
rect 35909 14365 35943 14399
rect 36185 14365 36219 14399
rect 20361 14297 20395 14331
rect 26525 14297 26559 14331
rect 26617 14297 26651 14331
rect 34897 14297 34931 14331
rect 35081 14297 35115 14331
rect 36093 14297 36127 14331
rect 2789 14229 2823 14263
rect 13277 14229 13311 14263
rect 13645 14229 13679 14263
rect 16037 14229 16071 14263
rect 1685 14025 1719 14059
rect 2605 14025 2639 14059
rect 2973 14025 3007 14059
rect 4813 14025 4847 14059
rect 14289 14025 14323 14059
rect 17509 14025 17543 14059
rect 33701 14025 33735 14059
rect 3801 13957 3835 13991
rect 13176 13957 13210 13991
rect 17233 13957 17267 13991
rect 19441 13957 19475 13991
rect 22385 13957 22419 13991
rect 1869 13889 1903 13923
rect 2053 13889 2087 13923
rect 2145 13889 2179 13923
rect 3985 13889 4019 13923
rect 4169 13889 4203 13923
rect 4261 13889 4295 13923
rect 4721 13889 4755 13923
rect 9036 13889 9070 13923
rect 14933 13889 14967 13923
rect 15117 13889 15151 13923
rect 15209 13889 15243 13923
rect 17417 13889 17451 13923
rect 18705 13889 18739 13923
rect 19165 13889 19199 13923
rect 22201 13889 22235 13923
rect 22477 13889 22511 13923
rect 23397 13889 23431 13923
rect 32577 13889 32611 13923
rect 3065 13821 3099 13855
rect 3249 13821 3283 13855
rect 8769 13821 8803 13855
rect 12909 13821 12943 13855
rect 22017 13821 22051 13855
rect 32321 13821 32355 13855
rect 10149 13685 10183 13719
rect 14749 13685 14783 13719
rect 24685 13685 24719 13719
rect 2881 13481 2915 13515
rect 4169 13481 4203 13515
rect 22109 13481 22143 13515
rect 32505 13481 32539 13515
rect 18797 13413 18831 13447
rect 17877 13345 17911 13379
rect 24593 13345 24627 13379
rect 3157 13277 3191 13311
rect 12173 13277 12207 13311
rect 17141 13277 17175 13311
rect 17785 13277 17819 13311
rect 18521 13277 18555 13311
rect 18705 13277 18739 13311
rect 19441 13277 19475 13311
rect 19625 13277 19659 13311
rect 20821 13277 20855 13311
rect 26433 13277 26467 13311
rect 29929 13277 29963 13311
rect 30205 13277 30239 13311
rect 2513 13209 2547 13243
rect 2890 13209 2924 13243
rect 3985 13209 4019 13243
rect 4169 13209 4203 13243
rect 7481 13209 7515 13243
rect 7573 13209 7607 13243
rect 7941 13209 7975 13243
rect 8309 13209 8343 13243
rect 10425 13209 10459 13243
rect 14289 13209 14323 13243
rect 19809 13209 19843 13243
rect 24860 13209 24894 13243
rect 31217 13209 31251 13243
rect 4353 13141 4387 13175
rect 7205 13141 7239 13175
rect 8493 13141 8527 13175
rect 15577 13141 15611 13175
rect 25973 13141 26007 13175
rect 26617 13141 26651 13175
rect 29745 13141 29779 13175
rect 30113 13141 30147 13175
rect 3433 12937 3467 12971
rect 6009 12937 6043 12971
rect 9781 12937 9815 12971
rect 10885 12937 10919 12971
rect 14749 12937 14783 12971
rect 17509 12937 17543 12971
rect 24685 12937 24719 12971
rect 27169 12937 27203 12971
rect 29929 12937 29963 12971
rect 31401 12937 31435 12971
rect 33701 12937 33735 12971
rect 2697 12869 2731 12903
rect 3249 12869 3283 12903
rect 10517 12869 10551 12903
rect 12449 12869 12483 12903
rect 12633 12869 12667 12903
rect 19257 12869 19291 12903
rect 19349 12869 19383 12903
rect 23397 12869 23431 12903
rect 27537 12869 27571 12903
rect 28641 12869 28675 12903
rect 2605 12801 2639 12835
rect 4629 12801 4663 12835
rect 4896 12801 4930 12835
rect 10057 12801 10091 12835
rect 10149 12801 10183 12835
rect 13369 12801 13403 12835
rect 13636 12801 13670 12835
rect 15393 12801 15427 12835
rect 15577 12801 15611 12835
rect 15669 12801 15703 12835
rect 16865 12801 16899 12835
rect 16958 12801 16992 12835
rect 17141 12801 17175 12835
rect 17233 12801 17267 12835
rect 17371 12801 17405 12835
rect 18981 12801 19015 12835
rect 19129 12801 19163 12835
rect 19446 12801 19480 12835
rect 25789 12801 25823 12835
rect 25973 12801 26007 12835
rect 26065 12801 26099 12835
rect 27353 12801 27387 12835
rect 27629 12801 27663 12835
rect 31217 12801 31251 12835
rect 31493 12801 31527 12835
rect 32321 12801 32355 12835
rect 31033 12733 31067 12767
rect 32597 12733 32631 12767
rect 19625 12665 19659 12699
rect 3433 12597 3467 12631
rect 3617 12597 3651 12631
rect 11069 12597 11103 12631
rect 12633 12597 12667 12631
rect 12817 12597 12851 12631
rect 15209 12597 15243 12631
rect 25605 12597 25639 12631
rect 6837 12393 6871 12427
rect 10517 12393 10551 12427
rect 15669 12393 15703 12427
rect 20085 12393 20119 12427
rect 23305 12393 23339 12427
rect 26801 12393 26835 12427
rect 27169 12393 27203 12427
rect 28089 12393 28123 12427
rect 26893 12257 26927 12291
rect 4077 12189 4111 12223
rect 4169 12189 4203 12223
rect 5457 12189 5491 12223
rect 5713 12189 5747 12223
rect 9137 12189 9171 12223
rect 13461 12189 13495 12223
rect 13737 12189 13771 12223
rect 14289 12189 14323 12223
rect 18153 12189 18187 12223
rect 18337 12189 18371 12223
rect 18521 12189 18555 12223
rect 19441 12189 19475 12223
rect 19534 12189 19568 12223
rect 19947 12189 19981 12223
rect 21189 12189 21223 12223
rect 21465 12189 21499 12223
rect 21925 12189 21959 12223
rect 26801 12189 26835 12223
rect 28273 12189 28307 12223
rect 28365 12189 28399 12223
rect 28733 12189 28767 12223
rect 9404 12121 9438 12155
rect 14556 12121 14590 12155
rect 18429 12121 18463 12155
rect 19717 12121 19751 12155
rect 19809 12121 19843 12155
rect 22192 12121 22226 12155
rect 24593 12121 24627 12155
rect 28457 12121 28491 12155
rect 28575 12121 28609 12155
rect 30849 12121 30883 12155
rect 4353 12053 4387 12087
rect 13277 12053 13311 12087
rect 13645 12053 13679 12087
rect 18705 12053 18739 12087
rect 21005 12053 21039 12087
rect 21373 12053 21407 12087
rect 25881 12053 25915 12087
rect 32137 12053 32171 12087
rect 23489 11849 23523 11883
rect 24133 11849 24167 11883
rect 24317 11849 24351 11883
rect 26525 11849 26559 11883
rect 28457 11849 28491 11883
rect 28641 11849 28675 11883
rect 32321 11849 32355 11883
rect 32689 11849 32723 11883
rect 23949 11781 23983 11815
rect 28273 11781 28307 11815
rect 31677 11781 31711 11815
rect 13001 11713 13035 11747
rect 22376 11713 22410 11747
rect 25881 11713 25915 11747
rect 25974 11713 26008 11747
rect 26157 11713 26191 11747
rect 26249 11713 26283 11747
rect 26387 11713 26421 11747
rect 29469 11713 29503 11747
rect 31493 11713 31527 11747
rect 31769 11713 31803 11747
rect 32505 11713 32539 11747
rect 32781 11713 32815 11747
rect 14749 11645 14783 11679
rect 22109 11645 22143 11679
rect 29193 11645 29227 11679
rect 30573 11645 30607 11679
rect 24133 11509 24167 11543
rect 28457 11509 28491 11543
rect 31309 11509 31343 11543
rect 15669 11305 15703 11339
rect 23397 11305 23431 11339
rect 32597 11305 32631 11339
rect 9137 11169 9171 11203
rect 31493 11169 31527 11203
rect 6193 11101 6227 11135
rect 9404 11101 9438 11135
rect 14289 11101 14323 11135
rect 14545 11101 14579 11135
rect 22017 11101 22051 11135
rect 22273 11101 22307 11135
rect 31217 11101 31251 11135
rect 5733 11033 5767 11067
rect 5825 11033 5859 11067
rect 6561 11033 6595 11067
rect 5457 10965 5491 10999
rect 6745 10965 6779 10999
rect 10517 10965 10551 10999
rect 5273 10761 5307 10795
rect 9781 10761 9815 10795
rect 14289 10761 14323 10795
rect 29929 10761 29963 10795
rect 10885 10693 10919 10727
rect 13001 10693 13035 10727
rect 18245 10693 18279 10727
rect 28641 10693 28675 10727
rect 3893 10625 3927 10659
rect 4160 10625 4194 10659
rect 10057 10625 10091 10659
rect 10149 10625 10183 10659
rect 10517 10625 10551 10659
rect 19993 10557 20027 10591
rect 11069 10421 11103 10455
rect 5365 10217 5399 10251
rect 10517 10217 10551 10251
rect 22109 10217 22143 10251
rect 26709 10217 26743 10251
rect 27997 10217 28031 10251
rect 3985 10081 4019 10115
rect 9137 10081 9171 10115
rect 19625 10013 19659 10047
rect 19901 10013 19935 10047
rect 20821 10013 20855 10047
rect 25053 10013 25087 10047
rect 25237 10013 25271 10047
rect 25329 10013 25363 10047
rect 26157 10013 26191 10047
rect 26433 10013 26467 10047
rect 26525 10013 26559 10047
rect 29929 10013 29963 10047
rect 30205 10013 30239 10047
rect 30849 10013 30883 10047
rect 31125 10013 31159 10047
rect 4252 9945 4286 9979
rect 9382 9945 9416 9979
rect 19809 9945 19843 9979
rect 26341 9945 26375 9979
rect 27813 9945 27847 9979
rect 29745 9945 29779 9979
rect 30113 9945 30147 9979
rect 31033 9945 31067 9979
rect 19441 9877 19475 9911
rect 24869 9877 24903 9911
rect 27997 9877 28031 9911
rect 28181 9877 28215 9911
rect 30665 9877 30699 9911
rect 20085 9673 20119 9707
rect 29193 9673 29227 9707
rect 15577 9605 15611 9639
rect 18972 9605 19006 9639
rect 20729 9605 20763 9639
rect 25421 9605 25455 9639
rect 25513 9605 25547 9639
rect 29653 9605 29687 9639
rect 2697 9537 2731 9571
rect 13001 9537 13035 9571
rect 15393 9537 15427 9571
rect 15669 9537 15703 9571
rect 20545 9537 20579 9571
rect 20817 9537 20851 9571
rect 20913 9537 20947 9571
rect 25237 9537 25271 9571
rect 25605 9537 25639 9571
rect 27813 9537 27847 9571
rect 28080 9537 28114 9571
rect 18705 9469 18739 9503
rect 21097 9401 21131 9435
rect 30941 9401 30975 9435
rect 2789 9333 2823 9367
rect 14289 9333 14323 9367
rect 15209 9333 15243 9367
rect 25789 9333 25823 9367
rect 3341 9129 3375 9163
rect 15669 9129 15703 9163
rect 18705 9129 18739 9163
rect 23581 9129 23615 9163
rect 25973 9129 26007 9163
rect 29193 9129 29227 9163
rect 31125 9129 31159 9163
rect 1869 8993 1903 9027
rect 14289 8993 14323 9027
rect 1593 8925 1627 8959
rect 16313 8925 16347 8959
rect 16497 8925 16531 8959
rect 16589 8925 16623 8959
rect 18153 8925 18187 8959
rect 18521 8925 18555 8959
rect 21833 8925 21867 8959
rect 22109 8925 22143 8959
rect 24593 8925 24627 8959
rect 24860 8925 24894 8959
rect 27813 8925 27847 8959
rect 29745 8925 29779 8959
rect 14556 8857 14590 8891
rect 16129 8857 16163 8891
rect 18337 8857 18371 8891
rect 18429 8857 18463 8891
rect 19441 8857 19475 8891
rect 23397 8857 23431 8891
rect 23581 8857 23615 8891
rect 28080 8857 28114 8891
rect 29990 8857 30024 8891
rect 20729 8789 20763 8823
rect 21649 8789 21683 8823
rect 22017 8789 22051 8823
rect 23765 8789 23799 8823
rect 13921 8585 13955 8619
rect 17049 8585 17083 8619
rect 18705 8585 18739 8619
rect 20637 8585 20671 8619
rect 25973 8585 26007 8619
rect 30573 8585 30607 8619
rect 30941 8585 30975 8619
rect 2973 8517 3007 8551
rect 4896 8517 4930 8551
rect 10977 8517 11011 8551
rect 16865 8517 16899 8551
rect 18337 8517 18371 8551
rect 18521 8517 18555 8551
rect 19524 8517 19558 8551
rect 24685 8517 24719 8551
rect 2697 8449 2731 8483
rect 2789 8449 2823 8483
rect 4629 8449 4663 8483
rect 6561 8449 6595 8483
rect 6745 8449 6779 8483
rect 10149 8449 10183 8483
rect 13737 8449 13771 8483
rect 14013 8449 14047 8483
rect 14473 8449 14507 8483
rect 17325 8449 17359 8483
rect 19257 8449 19291 8483
rect 22845 8449 22879 8483
rect 23101 8449 23135 8483
rect 28733 8449 28767 8483
rect 29000 8449 29034 8483
rect 30757 8449 30791 8483
rect 31033 8449 31067 8483
rect 10057 8381 10091 8415
rect 10609 8381 10643 8415
rect 13553 8381 13587 8415
rect 6009 8313 6043 8347
rect 10517 8313 10551 8347
rect 15761 8313 15795 8347
rect 30113 8313 30147 8347
rect 6653 8245 6687 8279
rect 17049 8245 17083 8279
rect 18521 8245 18555 8279
rect 24225 8245 24259 8279
rect 6929 8041 6963 8075
rect 10885 8041 10919 8075
rect 15853 8041 15887 8075
rect 20821 8041 20855 8075
rect 22845 8041 22879 8075
rect 26249 8041 26283 8075
rect 29745 8041 29779 8075
rect 5181 7905 5215 7939
rect 9137 7905 9171 7939
rect 9413 7905 9447 7939
rect 14473 7905 14507 7939
rect 4077 7837 4111 7871
rect 11437 7837 11471 7871
rect 11621 7837 11655 7871
rect 14740 7837 14774 7871
rect 16497 7837 16531 7871
rect 16681 7837 16715 7871
rect 16773 7837 16807 7871
rect 18613 7837 18647 7871
rect 18889 7837 18923 7871
rect 19441 7837 19475 7871
rect 23029 7837 23063 7871
rect 23305 7837 23339 7871
rect 24869 7837 24903 7871
rect 29929 7837 29963 7871
rect 30205 7837 30239 7871
rect 4261 7769 4295 7803
rect 5457 7769 5491 7803
rect 11713 7769 11747 7803
rect 19708 7769 19742 7803
rect 23213 7769 23247 7803
rect 25136 7769 25170 7803
rect 30113 7769 30147 7803
rect 16313 7701 16347 7735
rect 18429 7701 18463 7735
rect 18797 7701 18831 7735
rect 7021 7497 7055 7531
rect 15761 7497 15795 7531
rect 19533 7497 19567 7531
rect 20453 7497 20487 7531
rect 20821 7497 20855 7531
rect 24685 7497 24719 7531
rect 25605 7497 25639 7531
rect 25973 7497 26007 7531
rect 29929 7497 29963 7531
rect 6929 7429 6963 7463
rect 14648 7429 14682 7463
rect 18245 7429 18279 7463
rect 23397 7429 23431 7463
rect 28641 7429 28675 7463
rect 9577 7361 9611 7395
rect 12173 7361 12207 7395
rect 12357 7361 12391 7395
rect 14381 7361 14415 7395
rect 20637 7361 20671 7395
rect 20913 7361 20947 7395
rect 25789 7361 25823 7395
rect 26065 7361 26099 7395
rect 7205 7293 7239 7327
rect 9321 7293 9355 7327
rect 6561 7157 6595 7191
rect 10701 7157 10735 7191
rect 12173 7157 12207 7191
rect 6929 6817 6963 6851
rect 7021 6817 7055 6851
rect 10977 6817 11011 6851
rect 11069 6817 11103 6851
rect 6837 6749 6871 6783
rect 10885 6749 10919 6783
rect 14473 6749 14507 6783
rect 14740 6749 14774 6783
rect 24593 6749 24627 6783
rect 24860 6681 24894 6715
rect 6469 6613 6503 6647
rect 10517 6613 10551 6647
rect 15853 6613 15887 6647
rect 25973 6613 26007 6647
rect 12173 6409 12207 6443
rect 19901 6409 19935 6443
rect 25329 6409 25363 6443
rect 25697 6409 25731 6443
rect 12081 6341 12115 6375
rect 18766 6341 18800 6375
rect 25513 6273 25547 6307
rect 25789 6273 25823 6307
rect 12265 6205 12299 6239
rect 18521 6205 18555 6239
rect 11713 6069 11747 6103
rect 6745 5865 6779 5899
rect 4629 5729 4663 5763
rect 4997 5729 5031 5763
rect 27813 5729 27847 5763
rect 10149 5661 10183 5695
rect 28080 5593 28114 5627
rect 10241 5525 10275 5559
rect 29193 5525 29227 5559
rect 10149 5321 10183 5355
rect 14473 5321 14507 5355
rect 19533 5321 19567 5355
rect 24685 5321 24719 5355
rect 29929 5321 29963 5355
rect 5733 5253 5767 5287
rect 13001 5253 13035 5287
rect 18245 5253 18279 5287
rect 23397 5253 23431 5287
rect 28641 5253 28675 5287
rect 5457 5185 5491 5219
rect 5641 5185 5675 5219
rect 9965 5185 9999 5219
rect 10149 5185 10183 5219
rect 22109 5185 22143 5219
rect 22201 4981 22235 5015
rect 11161 4777 11195 4811
rect 28917 4777 28951 4811
rect 7849 4709 7883 4743
rect 10517 4709 10551 4743
rect 14289 4709 14323 4743
rect 21557 4709 21591 4743
rect 28641 4709 28675 4743
rect 28733 4709 28767 4743
rect 8493 4641 8527 4675
rect 9597 4641 9631 4675
rect 9689 4641 9723 4675
rect 10609 4641 10643 4675
rect 22201 4641 22235 4675
rect 28825 4641 28859 4675
rect 6377 4573 6411 4607
rect 6561 4573 6595 4607
rect 8217 4573 8251 4607
rect 10333 4573 10367 4607
rect 10425 4573 10459 4607
rect 11069 4573 11103 4607
rect 11345 4573 11379 4607
rect 12725 4573 12759 4607
rect 14565 4573 14599 4607
rect 15025 4573 15059 4607
rect 17785 4573 17819 4607
rect 19625 4573 19659 4607
rect 21925 4573 21959 4607
rect 22937 4573 22971 4607
rect 23213 4573 23247 4607
rect 24593 4573 24627 4607
rect 26433 4573 26467 4607
rect 28273 4573 28307 4607
rect 6745 4505 6779 4539
rect 8309 4505 8343 4539
rect 9505 4505 9539 4539
rect 14289 4505 14323 4539
rect 26700 4505 26734 4539
rect 9137 4437 9171 4471
rect 11621 4437 11655 4471
rect 12817 4437 12851 4471
rect 14473 4437 14507 4471
rect 15117 4437 15151 4471
rect 17877 4437 17911 4471
rect 19717 4437 19751 4471
rect 22017 4437 22051 4471
rect 22753 4437 22787 4471
rect 23121 4437 23155 4471
rect 24685 4437 24719 4471
rect 27813 4437 27847 4471
rect 7941 4233 7975 4267
rect 10701 4233 10735 4267
rect 23397 4233 23431 4267
rect 28549 4233 28583 4267
rect 22284 4165 22318 4199
rect 6817 4097 6851 4131
rect 8953 4097 8987 4131
rect 12633 4097 12667 4131
rect 12900 4097 12934 4131
rect 14473 4097 14507 4131
rect 14740 4097 14774 4131
rect 16865 4097 16899 4131
rect 17693 4097 17727 4131
rect 17960 4097 17994 4131
rect 19533 4097 19567 4131
rect 19800 4097 19834 4131
rect 22017 4097 22051 4131
rect 23857 4097 23891 4131
rect 24124 4097 24158 4131
rect 27169 4097 27203 4131
rect 27425 4097 27459 4131
rect 29009 4097 29043 4131
rect 29265 4097 29299 4131
rect 6561 4029 6595 4063
rect 9229 4029 9263 4063
rect 26157 4029 26191 4063
rect 26617 4029 26651 4063
rect 15853 3961 15887 3995
rect 26525 3961 26559 3995
rect 14013 3893 14047 3927
rect 16957 3893 16991 3927
rect 19073 3893 19107 3927
rect 20913 3893 20947 3927
rect 25237 3893 25271 3927
rect 30389 3893 30423 3927
rect 7389 3689 7423 3723
rect 10885 3689 10919 3723
rect 14841 3689 14875 3723
rect 19809 3689 19843 3723
rect 23949 3689 23983 3723
rect 24593 3689 24627 3723
rect 26801 3689 26835 3723
rect 27721 3689 27755 3723
rect 29101 3689 29135 3723
rect 27629 3621 27663 3655
rect 28917 3621 28951 3655
rect 5917 3553 5951 3587
rect 15393 3553 15427 3587
rect 16589 3553 16623 3587
rect 20453 3553 20487 3587
rect 25053 3553 25087 3587
rect 25237 3553 25271 3587
rect 27813 3553 27847 3587
rect 5641 3485 5675 3519
rect 9505 3485 9539 3519
rect 20177 3485 20211 3519
rect 20269 3485 20303 3519
rect 22569 3485 22603 3519
rect 22836 3485 22870 3519
rect 26617 3485 26651 3519
rect 27261 3485 27295 3519
rect 9750 3417 9784 3451
rect 15209 3417 15243 3451
rect 16856 3417 16890 3451
rect 24961 3417 24995 3451
rect 25605 3417 25639 3451
rect 26433 3417 26467 3451
rect 28641 3417 28675 3451
rect 15301 3349 15335 3383
rect 17969 3349 18003 3383
rect 28089 3349 28123 3383
rect 14105 3145 14139 3179
rect 14565 3145 14599 3179
rect 16865 3145 16899 3179
rect 17233 3145 17267 3179
rect 17325 3145 17359 3179
rect 18429 3145 18463 3179
rect 22753 3145 22787 3179
rect 27997 3145 28031 3179
rect 1593 3009 1627 3043
rect 9873 3009 9907 3043
rect 10057 3009 10091 3043
rect 14473 3009 14507 3043
rect 18797 3009 18831 3043
rect 18889 3009 18923 3043
rect 22661 3009 22695 3043
rect 1777 2941 1811 2975
rect 10241 2941 10275 2975
rect 14749 2941 14783 2975
rect 17509 2941 17543 2975
rect 19073 2941 19107 2975
rect 27537 2941 27571 2975
rect 38117 2941 38151 2975
rect 27905 2873 27939 2907
rect 2421 2397 2455 2431
rect 3985 2397 4019 2431
rect 5365 2397 5399 2431
rect 7021 2397 7055 2431
rect 8493 2397 8527 2431
rect 9965 2397 9999 2431
rect 11897 2397 11931 2431
rect 12909 2397 12943 2431
rect 14473 2397 14507 2431
rect 15669 2397 15703 2431
rect 17141 2397 17175 2431
rect 18429 2397 18463 2431
rect 20085 2397 20119 2431
rect 22017 2397 22051 2431
rect 23029 2397 23063 2431
rect 24593 2397 24627 2431
rect 25973 2397 26007 2431
rect 27445 2397 27479 2431
rect 29745 2397 29779 2431
rect 30665 2397 30699 2431
rect 32321 2397 32355 2431
rect 33517 2397 33551 2431
rect 35081 2397 35115 2431
rect 36461 2397 36495 2431
rect 37933 2397 37967 2431
rect 2697 2329 2731 2363
rect 4261 2329 4295 2363
rect 5641 2329 5675 2363
rect 15945 2329 15979 2363
rect 17417 2329 17451 2363
rect 18705 2329 18739 2363
rect 20361 2329 20395 2363
rect 22293 2329 22327 2363
rect 23305 2329 23339 2363
rect 24869 2329 24903 2363
rect 26249 2329 26283 2363
rect 27721 2329 27755 2363
rect 30021 2329 30055 2363
rect 30941 2329 30975 2363
rect 32597 2329 32631 2363
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 17218 37408 17224 37460
rect 17276 37448 17282 37460
rect 32493 37451 32551 37457
rect 32493 37448 32505 37451
rect 17276 37420 32505 37448
rect 17276 37408 17282 37420
rect 32493 37417 32505 37420
rect 32539 37417 32551 37451
rect 32493 37411 32551 37417
rect 12069 37383 12127 37389
rect 12069 37349 12081 37383
rect 12115 37380 12127 37383
rect 14274 37380 14280 37392
rect 12115 37352 14280 37380
rect 12115 37349 12127 37352
rect 12069 37343 12127 37349
rect 14274 37340 14280 37352
rect 14332 37340 14338 37392
rect 14918 37340 14924 37392
rect 14976 37380 14982 37392
rect 28629 37383 28687 37389
rect 28629 37380 28641 37383
rect 14976 37352 28641 37380
rect 14976 37340 14982 37352
rect 28629 37349 28641 37352
rect 28675 37349 28687 37383
rect 28629 37343 28687 37349
rect 5442 37312 5448 37324
rect 5403 37284 5448 37312
rect 5442 37272 5448 37284
rect 5500 37272 5506 37324
rect 9401 37315 9459 37321
rect 9401 37281 9413 37315
rect 9447 37312 9459 37315
rect 13446 37312 13452 37324
rect 9447 37284 13452 37312
rect 9447 37281 9459 37284
rect 9401 37275 9459 37281
rect 13446 37272 13452 37284
rect 13504 37272 13510 37324
rect 37182 37272 37188 37324
rect 37240 37312 37246 37324
rect 38289 37315 38347 37321
rect 38289 37312 38301 37315
rect 37240 37284 38301 37312
rect 37240 37272 37246 37284
rect 38289 37281 38301 37284
rect 38335 37281 38347 37315
rect 38289 37275 38347 37281
rect 5074 37204 5080 37256
rect 5132 37244 5138 37256
rect 5261 37247 5319 37253
rect 5261 37244 5273 37247
rect 5132 37216 5273 37244
rect 5132 37204 5138 37216
rect 5261 37213 5273 37216
rect 5307 37213 5319 37247
rect 5261 37207 5319 37213
rect 8386 37204 8392 37256
rect 8444 37244 8450 37256
rect 9217 37247 9275 37253
rect 9217 37244 9229 37247
rect 8444 37216 9229 37244
rect 8444 37204 8450 37216
rect 9217 37213 9229 37216
rect 9263 37213 9275 37247
rect 9217 37207 9275 37213
rect 11698 37204 11704 37256
rect 11756 37244 11762 37256
rect 11885 37247 11943 37253
rect 11885 37244 11897 37247
rect 11756 37216 11897 37244
rect 11756 37204 11762 37216
rect 11885 37213 11897 37216
rect 11931 37213 11943 37247
rect 15194 37244 15200 37256
rect 15155 37216 15200 37244
rect 11885 37207 11943 37213
rect 15194 37204 15200 37216
rect 15252 37204 15258 37256
rect 18322 37204 18328 37256
rect 18380 37244 18386 37256
rect 18509 37247 18567 37253
rect 18509 37244 18521 37247
rect 18380 37216 18521 37244
rect 18380 37204 18386 37216
rect 18509 37213 18521 37216
rect 18555 37213 18567 37247
rect 18509 37207 18567 37213
rect 24946 37204 24952 37256
rect 25004 37244 25010 37256
rect 25133 37247 25191 37253
rect 25133 37244 25145 37247
rect 25004 37216 25145 37244
rect 25004 37204 25010 37216
rect 25133 37213 25145 37216
rect 25179 37213 25191 37247
rect 25133 37207 25191 37213
rect 28258 37204 28264 37256
rect 28316 37244 28322 37256
rect 28445 37247 28503 37253
rect 28445 37244 28457 37247
rect 28316 37216 28457 37244
rect 28316 37204 28322 37216
rect 28445 37213 28457 37216
rect 28491 37213 28503 37247
rect 28445 37207 28503 37213
rect 31754 37204 31760 37256
rect 31812 37244 31818 37256
rect 32401 37247 32459 37253
rect 32401 37244 32413 37247
rect 31812 37216 32413 37244
rect 31812 37204 31818 37216
rect 32401 37213 32413 37216
rect 32447 37213 32459 37247
rect 32401 37207 32459 37213
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 35069 37247 35127 37253
rect 35069 37244 35081 37247
rect 34848 37216 35081 37244
rect 34848 37204 34854 37216
rect 35069 37213 35081 37216
rect 35115 37213 35127 37247
rect 35069 37207 35127 37213
rect 38105 37247 38163 37253
rect 38105 37213 38117 37247
rect 38151 37244 38163 37247
rect 38194 37244 38200 37256
rect 38151 37216 38200 37244
rect 38151 37213 38163 37216
rect 38105 37207 38163 37213
rect 38194 37204 38200 37216
rect 38252 37204 38258 37256
rect 22094 37136 22100 37188
rect 22152 37176 22158 37188
rect 22152 37148 22197 37176
rect 22152 37136 22158 37148
rect 15286 37108 15292 37120
rect 15247 37080 15292 37108
rect 15286 37068 15292 37080
rect 15344 37068 15350 37120
rect 18598 37108 18604 37120
rect 18559 37080 18604 37108
rect 18598 37068 18604 37080
rect 18656 37068 18662 37120
rect 22186 37108 22192 37120
rect 22147 37080 22192 37108
rect 22186 37068 22192 37080
rect 22244 37068 22250 37120
rect 25222 37108 25228 37120
rect 25183 37080 25228 37108
rect 25222 37068 25228 37080
rect 25280 37068 25286 37120
rect 34514 37068 34520 37120
rect 34572 37108 34578 37120
rect 35161 37111 35219 37117
rect 35161 37108 35173 37111
rect 34572 37080 35173 37108
rect 34572 37068 34578 37080
rect 35161 37077 35173 37080
rect 35207 37077 35219 37111
rect 35161 37071 35219 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 13446 36864 13452 36916
rect 13504 36904 13510 36916
rect 14277 36907 14335 36913
rect 14277 36904 14289 36907
rect 13504 36876 14289 36904
rect 13504 36864 13510 36876
rect 14277 36873 14289 36876
rect 14323 36873 14335 36907
rect 22186 36904 22192 36916
rect 14277 36867 14335 36873
rect 15856 36876 22192 36904
rect 14185 36839 14243 36845
rect 14185 36805 14197 36839
rect 14231 36836 14243 36839
rect 15856 36836 15884 36876
rect 22186 36864 22192 36876
rect 22244 36864 22250 36916
rect 14231 36808 15884 36836
rect 14231 36805 14243 36808
rect 14185 36799 14243 36805
rect 19426 36796 19432 36848
rect 19484 36796 19490 36848
rect 18601 36771 18659 36777
rect 18601 36737 18613 36771
rect 18647 36768 18659 36771
rect 18690 36768 18696 36780
rect 18647 36740 18696 36768
rect 18647 36737 18659 36740
rect 18601 36731 18659 36737
rect 18690 36728 18696 36740
rect 18748 36728 18754 36780
rect 19061 36771 19119 36777
rect 19061 36737 19073 36771
rect 19107 36768 19119 36771
rect 20070 36768 20076 36780
rect 19107 36740 20076 36768
rect 19107 36737 19119 36740
rect 19061 36731 19119 36737
rect 20070 36728 20076 36740
rect 20128 36728 20134 36780
rect 25130 36768 25136 36780
rect 25091 36740 25136 36768
rect 25130 36728 25136 36740
rect 25188 36728 25194 36780
rect 25498 36728 25504 36780
rect 25556 36768 25562 36780
rect 25961 36771 26019 36777
rect 25961 36768 25973 36771
rect 25556 36740 25973 36768
rect 25556 36728 25562 36740
rect 25961 36737 25973 36740
rect 26007 36737 26019 36771
rect 26142 36768 26148 36780
rect 26103 36740 26148 36768
rect 25961 36731 26019 36737
rect 26142 36728 26148 36740
rect 26200 36728 26206 36780
rect 30101 36771 30159 36777
rect 30101 36737 30113 36771
rect 30147 36737 30159 36771
rect 30101 36731 30159 36737
rect 30285 36771 30343 36777
rect 30285 36737 30297 36771
rect 30331 36768 30343 36771
rect 31018 36768 31024 36780
rect 30331 36740 31024 36768
rect 30331 36737 30343 36740
rect 30285 36731 30343 36737
rect 14458 36700 14464 36712
rect 14419 36672 14464 36700
rect 14458 36660 14464 36672
rect 14516 36660 14522 36712
rect 25038 36700 25044 36712
rect 24999 36672 25044 36700
rect 25038 36660 25044 36672
rect 25096 36660 25102 36712
rect 30116 36700 30144 36731
rect 31018 36728 31024 36740
rect 31076 36728 31082 36780
rect 31202 36700 31208 36712
rect 30116 36672 31208 36700
rect 31202 36660 31208 36672
rect 31260 36660 31266 36712
rect 25501 36635 25559 36641
rect 25501 36601 25513 36635
rect 25547 36632 25559 36635
rect 26050 36632 26056 36644
rect 25547 36604 26056 36632
rect 25547 36601 25559 36604
rect 25501 36595 25559 36601
rect 26050 36592 26056 36604
rect 26108 36592 26114 36644
rect 13814 36564 13820 36576
rect 13775 36536 13820 36564
rect 13814 36524 13820 36536
rect 13872 36524 13878 36576
rect 25866 36524 25872 36576
rect 25924 36564 25930 36576
rect 25961 36567 26019 36573
rect 25961 36564 25973 36567
rect 25924 36536 25973 36564
rect 25924 36524 25930 36536
rect 25961 36533 25973 36536
rect 26007 36533 26019 36567
rect 30098 36564 30104 36576
rect 30059 36536 30104 36564
rect 25961 36527 26019 36533
rect 30098 36524 30104 36536
rect 30156 36524 30162 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 24857 36363 24915 36369
rect 24857 36329 24869 36363
rect 24903 36360 24915 36363
rect 26142 36360 26148 36372
rect 24903 36332 26148 36360
rect 24903 36329 24915 36332
rect 24857 36323 24915 36329
rect 26142 36320 26148 36332
rect 26200 36320 26206 36372
rect 30374 36320 30380 36372
rect 30432 36360 30438 36372
rect 30837 36363 30895 36369
rect 30837 36360 30849 36363
rect 30432 36332 30849 36360
rect 30432 36320 30438 36332
rect 30837 36329 30849 36332
rect 30883 36329 30895 36363
rect 31018 36360 31024 36372
rect 30979 36332 31024 36360
rect 30837 36323 30895 36329
rect 31018 36320 31024 36332
rect 31076 36320 31082 36372
rect 14182 36252 14188 36304
rect 14240 36292 14246 36304
rect 14553 36295 14611 36301
rect 14553 36292 14565 36295
rect 14240 36264 14565 36292
rect 14240 36252 14246 36264
rect 14553 36261 14565 36264
rect 14599 36261 14611 36295
rect 14553 36255 14611 36261
rect 15746 36252 15752 36304
rect 15804 36292 15810 36304
rect 37001 36295 37059 36301
rect 37001 36292 37013 36295
rect 15804 36264 37013 36292
rect 15804 36252 15810 36264
rect 37001 36261 37013 36264
rect 37047 36261 37059 36295
rect 37001 36255 37059 36261
rect 14918 36224 14924 36236
rect 14879 36196 14924 36224
rect 14918 36184 14924 36196
rect 14976 36184 14982 36236
rect 17218 36224 17224 36236
rect 17179 36196 17224 36224
rect 17218 36184 17224 36196
rect 17276 36184 17282 36236
rect 18598 36224 18604 36236
rect 17328 36196 18604 36224
rect 17328 36165 17356 36196
rect 18598 36184 18604 36196
rect 18656 36184 18662 36236
rect 25866 36224 25872 36236
rect 25827 36196 25872 36224
rect 25866 36184 25872 36196
rect 25924 36184 25930 36236
rect 26050 36224 26056 36236
rect 26011 36196 26056 36224
rect 26050 36184 26056 36196
rect 26108 36184 26114 36236
rect 29733 36227 29791 36233
rect 29733 36224 29745 36227
rect 29012 36196 29745 36224
rect 17313 36159 17371 36165
rect 17313 36125 17325 36159
rect 17359 36125 17371 36159
rect 17313 36119 17371 36125
rect 17402 36116 17408 36168
rect 17460 36156 17466 36168
rect 17497 36159 17555 36165
rect 17497 36156 17509 36159
rect 17460 36128 17509 36156
rect 17460 36116 17466 36128
rect 17497 36125 17509 36128
rect 17543 36125 17555 36159
rect 24762 36156 24768 36168
rect 24723 36128 24768 36156
rect 17497 36119 17555 36125
rect 24762 36116 24768 36128
rect 24820 36116 24826 36168
rect 29012 36165 29040 36196
rect 29733 36193 29745 36196
rect 29779 36193 29791 36227
rect 33226 36224 33232 36236
rect 33187 36196 33232 36224
rect 29733 36187 29791 36193
rect 33226 36184 33232 36196
rect 33284 36184 33290 36236
rect 28997 36159 29055 36165
rect 28997 36156 29009 36159
rect 25424 36128 29009 36156
rect 14458 36048 14464 36100
rect 14516 36088 14522 36100
rect 15105 36091 15163 36097
rect 15105 36088 15117 36091
rect 14516 36060 15117 36088
rect 14516 36048 14522 36060
rect 15105 36057 15117 36060
rect 15151 36088 15163 36091
rect 17420 36088 17448 36116
rect 15151 36060 17448 36088
rect 15151 36057 15163 36060
rect 15105 36051 15163 36057
rect 17770 36048 17776 36100
rect 17828 36088 17834 36100
rect 17957 36091 18015 36097
rect 17957 36088 17969 36091
rect 17828 36060 17969 36088
rect 17828 36048 17834 36060
rect 17957 36057 17969 36060
rect 18003 36057 18015 36091
rect 17957 36051 18015 36057
rect 15013 36023 15071 36029
rect 15013 35989 15025 36023
rect 15059 36020 15071 36023
rect 15286 36020 15292 36032
rect 15059 35992 15292 36020
rect 15059 35989 15071 35992
rect 15013 35983 15071 35989
rect 15286 35980 15292 35992
rect 15344 35980 15350 36032
rect 25424 36029 25452 36128
rect 28997 36125 29009 36128
rect 29043 36125 29055 36159
rect 28997 36119 29055 36125
rect 29086 36116 29092 36168
rect 29144 36156 29150 36168
rect 29181 36159 29239 36165
rect 29181 36156 29193 36159
rect 29144 36128 29193 36156
rect 29144 36116 29150 36128
rect 29181 36125 29193 36128
rect 29227 36156 29239 36159
rect 30009 36159 30067 36165
rect 30009 36156 30021 36159
rect 29227 36128 30021 36156
rect 29227 36125 29239 36128
rect 29181 36119 29239 36125
rect 30009 36125 30021 36128
rect 30055 36125 30067 36159
rect 30009 36119 30067 36125
rect 30193 36159 30251 36165
rect 30193 36125 30205 36159
rect 30239 36125 30251 36159
rect 30193 36119 30251 36125
rect 25777 36091 25835 36097
rect 25777 36057 25789 36091
rect 25823 36088 25835 36091
rect 26142 36088 26148 36100
rect 25823 36060 26148 36088
rect 25823 36057 25835 36060
rect 25777 36051 25835 36057
rect 26142 36048 26148 36060
rect 26200 36048 26206 36100
rect 29454 36048 29460 36100
rect 29512 36088 29518 36100
rect 30208 36088 30236 36119
rect 30374 36116 30380 36168
rect 30432 36156 30438 36168
rect 31386 36156 31392 36168
rect 30432 36128 31392 36156
rect 30432 36116 30438 36128
rect 31386 36116 31392 36128
rect 31444 36116 31450 36168
rect 33321 36159 33379 36165
rect 33321 36125 33333 36159
rect 33367 36156 33379 36159
rect 33410 36156 33416 36168
rect 33367 36128 33416 36156
rect 33367 36125 33379 36128
rect 33321 36119 33379 36125
rect 33410 36116 33416 36128
rect 33468 36116 33474 36168
rect 34149 36159 34207 36165
rect 34149 36125 34161 36159
rect 34195 36156 34207 36159
rect 34514 36156 34520 36168
rect 34195 36128 34520 36156
rect 34195 36125 34207 36128
rect 34149 36119 34207 36125
rect 34514 36116 34520 36128
rect 34572 36116 34578 36168
rect 37182 36156 37188 36168
rect 37143 36128 37188 36156
rect 37182 36116 37188 36128
rect 37240 36116 37246 36168
rect 29512 36060 30236 36088
rect 29512 36048 29518 36060
rect 30466 36048 30472 36100
rect 30524 36088 30530 36100
rect 30653 36091 30711 36097
rect 30653 36088 30665 36091
rect 30524 36060 30665 36088
rect 30524 36048 30530 36060
rect 30653 36057 30665 36060
rect 30699 36057 30711 36091
rect 30653 36051 30711 36057
rect 25409 36023 25467 36029
rect 25409 35989 25421 36023
rect 25455 35989 25467 36023
rect 29178 36020 29184 36032
rect 29139 35992 29184 36020
rect 25409 35983 25467 35989
rect 29178 35980 29184 35992
rect 29236 35980 29242 36032
rect 29917 36023 29975 36029
rect 29917 35989 29929 36023
rect 29963 36020 29975 36023
rect 30282 36020 30288 36032
rect 29963 35992 30288 36020
rect 29963 35989 29975 35992
rect 29917 35983 29975 35989
rect 30282 35980 30288 35992
rect 30340 35980 30346 36032
rect 30834 35980 30840 36032
rect 30892 36029 30898 36032
rect 30892 36023 30911 36029
rect 30899 35989 30911 36023
rect 30892 35983 30911 35989
rect 33689 36023 33747 36029
rect 33689 35989 33701 36023
rect 33735 36020 33747 36023
rect 34054 36020 34060 36032
rect 33735 35992 34060 36020
rect 33735 35989 33747 35992
rect 33689 35983 33747 35989
rect 30892 35980 30898 35983
rect 34054 35980 34060 35992
rect 34112 35980 34118 36032
rect 34238 36020 34244 36032
rect 34199 35992 34244 36020
rect 34238 35980 34244 35992
rect 34296 35980 34302 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 14274 35816 14280 35828
rect 14235 35788 14280 35816
rect 14274 35776 14280 35788
rect 14332 35776 14338 35828
rect 21453 35819 21511 35825
rect 21453 35785 21465 35819
rect 21499 35816 21511 35819
rect 22557 35819 22615 35825
rect 22557 35816 22569 35819
rect 21499 35788 22569 35816
rect 21499 35785 21511 35788
rect 21453 35779 21511 35785
rect 22557 35785 22569 35788
rect 22603 35785 22615 35819
rect 25130 35816 25136 35828
rect 22557 35779 22615 35785
rect 23032 35788 25136 35816
rect 14185 35751 14243 35757
rect 14185 35717 14197 35751
rect 14231 35748 14243 35751
rect 22830 35748 22836 35760
rect 14231 35720 22836 35748
rect 14231 35717 14243 35720
rect 14185 35711 14243 35717
rect 22830 35708 22836 35720
rect 22888 35708 22894 35760
rect 18782 35680 18788 35692
rect 18743 35652 18788 35680
rect 18782 35640 18788 35652
rect 18840 35640 18846 35692
rect 19426 35680 19432 35692
rect 19387 35652 19432 35680
rect 19426 35640 19432 35652
rect 19484 35640 19490 35692
rect 21174 35640 21180 35692
rect 21232 35680 21238 35692
rect 21269 35683 21327 35689
rect 21269 35680 21281 35683
rect 21232 35652 21281 35680
rect 21232 35640 21238 35652
rect 21269 35649 21281 35652
rect 21315 35649 21327 35683
rect 21269 35643 21327 35649
rect 21453 35683 21511 35689
rect 21453 35649 21465 35683
rect 21499 35680 21511 35683
rect 22002 35680 22008 35692
rect 21499 35652 22008 35680
rect 21499 35649 21511 35652
rect 21453 35643 21511 35649
rect 14458 35612 14464 35624
rect 14419 35584 14464 35612
rect 14458 35572 14464 35584
rect 14516 35572 14522 35624
rect 20530 35572 20536 35624
rect 20588 35612 20594 35624
rect 21468 35612 21496 35643
rect 22002 35640 22008 35652
rect 22060 35680 22066 35692
rect 22373 35683 22431 35689
rect 22373 35680 22385 35683
rect 22060 35652 22385 35680
rect 22060 35640 22066 35652
rect 22373 35649 22385 35652
rect 22419 35680 22431 35683
rect 23032 35680 23060 35788
rect 25130 35776 25136 35788
rect 25188 35816 25194 35828
rect 30466 35816 30472 35828
rect 25188 35788 30472 35816
rect 25188 35776 25194 35788
rect 30466 35776 30472 35788
rect 30524 35776 30530 35828
rect 34793 35819 34851 35825
rect 34793 35816 34805 35819
rect 31036 35788 34805 35816
rect 23106 35708 23112 35760
rect 23164 35748 23170 35760
rect 25222 35748 25228 35760
rect 23164 35720 25228 35748
rect 23164 35708 23170 35720
rect 25222 35708 25228 35720
rect 25280 35708 25286 35760
rect 28997 35751 29055 35757
rect 28997 35717 29009 35751
rect 29043 35748 29055 35751
rect 30282 35748 30288 35760
rect 29043 35720 29868 35748
rect 30243 35720 30288 35748
rect 29043 35717 29055 35720
rect 28997 35711 29055 35717
rect 23198 35680 23204 35692
rect 22419 35652 23060 35680
rect 23159 35652 23204 35680
rect 22419 35649 22431 35652
rect 22373 35643 22431 35649
rect 23198 35640 23204 35652
rect 23256 35640 23262 35692
rect 23382 35680 23388 35692
rect 23343 35652 23388 35680
rect 23382 35640 23388 35652
rect 23440 35640 23446 35692
rect 25777 35683 25835 35689
rect 25777 35680 25789 35683
rect 24780 35652 25789 35680
rect 24780 35624 24808 35652
rect 25777 35649 25789 35652
rect 25823 35649 25835 35683
rect 25777 35643 25835 35649
rect 28905 35683 28963 35689
rect 28905 35649 28917 35683
rect 28951 35680 28963 35683
rect 29089 35683 29147 35689
rect 28951 35652 29040 35680
rect 28951 35649 28963 35652
rect 28905 35643 28963 35649
rect 29012 35624 29040 35652
rect 29089 35649 29101 35683
rect 29135 35680 29147 35683
rect 29454 35680 29460 35692
rect 29135 35652 29460 35680
rect 29135 35649 29147 35652
rect 29089 35643 29147 35649
rect 29454 35640 29460 35652
rect 29512 35640 29518 35692
rect 29840 35689 29868 35720
rect 30282 35708 30288 35720
rect 30340 35708 30346 35760
rect 29825 35683 29883 35689
rect 29825 35649 29837 35683
rect 29871 35649 29883 35683
rect 29825 35643 29883 35649
rect 29917 35683 29975 35689
rect 29917 35649 29929 35683
rect 29963 35680 29975 35683
rect 30374 35680 30380 35692
rect 29963 35652 30380 35680
rect 29963 35649 29975 35652
rect 29917 35643 29975 35649
rect 30374 35640 30380 35652
rect 30432 35640 30438 35692
rect 30466 35640 30472 35692
rect 30524 35680 30530 35692
rect 31036 35680 31064 35788
rect 34793 35785 34805 35788
rect 34839 35785 34851 35819
rect 34793 35779 34851 35785
rect 31386 35748 31392 35760
rect 31347 35720 31392 35748
rect 31386 35708 31392 35720
rect 31444 35708 31450 35760
rect 31205 35683 31263 35689
rect 31205 35680 31217 35683
rect 30524 35652 31217 35680
rect 30524 35640 30530 35652
rect 31205 35649 31217 35652
rect 31251 35649 31263 35683
rect 31481 35683 31539 35689
rect 31481 35680 31493 35683
rect 31205 35643 31263 35649
rect 31312 35652 31493 35680
rect 22646 35612 22652 35624
rect 20588 35584 21496 35612
rect 22607 35584 22652 35612
rect 20588 35572 20594 35584
rect 22646 35572 22652 35584
rect 22704 35572 22710 35624
rect 23750 35612 23756 35624
rect 23308 35584 23756 35612
rect 20257 35547 20315 35553
rect 20257 35513 20269 35547
rect 20303 35544 20315 35547
rect 23308 35544 23336 35584
rect 23750 35572 23756 35584
rect 23808 35612 23814 35624
rect 24762 35612 24768 35624
rect 23808 35584 24768 35612
rect 23808 35572 23814 35584
rect 24762 35572 24768 35584
rect 24820 35572 24826 35624
rect 24946 35612 24952 35624
rect 24907 35584 24952 35612
rect 24946 35572 24952 35584
rect 25004 35572 25010 35624
rect 25498 35612 25504 35624
rect 25459 35584 25504 35612
rect 25498 35572 25504 35584
rect 25556 35572 25562 35624
rect 25961 35615 26019 35621
rect 25961 35581 25973 35615
rect 26007 35581 26019 35615
rect 25961 35575 26019 35581
rect 23474 35544 23480 35556
rect 20303 35516 23336 35544
rect 23435 35516 23480 35544
rect 20303 35513 20315 35516
rect 20257 35507 20315 35513
rect 23474 35504 23480 35516
rect 23532 35504 23538 35556
rect 24210 35504 24216 35556
rect 24268 35544 24274 35556
rect 25976 35544 26004 35575
rect 28994 35572 29000 35624
rect 29052 35572 29058 35624
rect 30009 35615 30067 35621
rect 30009 35581 30021 35615
rect 30055 35612 30067 35615
rect 30834 35612 30840 35624
rect 30055 35584 30840 35612
rect 30055 35581 30067 35584
rect 30009 35575 30067 35581
rect 30834 35572 30840 35584
rect 30892 35612 30898 35624
rect 31312 35612 31340 35652
rect 31481 35649 31493 35652
rect 31527 35649 31539 35683
rect 32950 35680 32956 35692
rect 32911 35652 32956 35680
rect 31481 35643 31539 35649
rect 32950 35640 32956 35652
rect 33008 35640 33014 35692
rect 33505 35683 33563 35689
rect 33505 35649 33517 35683
rect 33551 35649 33563 35683
rect 33781 35683 33839 35689
rect 33781 35680 33793 35683
rect 33505 35643 33563 35649
rect 33612 35652 33793 35680
rect 30892 35584 31340 35612
rect 30892 35572 30898 35584
rect 32122 35572 32128 35624
rect 32180 35612 32186 35624
rect 33520 35612 33548 35643
rect 32180 35584 33548 35612
rect 32180 35572 32186 35584
rect 33612 35556 33640 35652
rect 33781 35649 33793 35652
rect 33827 35649 33839 35683
rect 33781 35643 33839 35649
rect 34422 35640 34428 35692
rect 34480 35680 34486 35692
rect 34701 35683 34759 35689
rect 34701 35680 34713 35683
rect 34480 35652 34713 35680
rect 34480 35640 34486 35652
rect 34701 35649 34713 35652
rect 34747 35649 34759 35683
rect 34701 35643 34759 35649
rect 29638 35544 29644 35556
rect 24268 35516 29644 35544
rect 24268 35504 24274 35516
rect 29638 35504 29644 35516
rect 29696 35504 29702 35556
rect 30745 35547 30803 35553
rect 30745 35513 30757 35547
rect 30791 35544 30803 35547
rect 33594 35544 33600 35556
rect 30791 35516 33600 35544
rect 30791 35513 30803 35516
rect 30745 35507 30803 35513
rect 33594 35504 33600 35516
rect 33652 35504 33658 35556
rect 13817 35479 13875 35485
rect 13817 35445 13829 35479
rect 13863 35476 13875 35479
rect 14090 35476 14096 35488
rect 13863 35448 14096 35476
rect 13863 35445 13875 35448
rect 13817 35439 13875 35445
rect 14090 35436 14096 35448
rect 14148 35436 14154 35488
rect 22097 35479 22155 35485
rect 22097 35445 22109 35479
rect 22143 35476 22155 35479
rect 25498 35476 25504 35488
rect 22143 35448 25504 35476
rect 22143 35445 22155 35448
rect 22097 35439 22155 35445
rect 25498 35436 25504 35448
rect 25556 35436 25562 35488
rect 31202 35476 31208 35488
rect 31163 35448 31208 35476
rect 31202 35436 31208 35448
rect 31260 35436 31266 35488
rect 33134 35476 33140 35488
rect 33095 35448 33140 35476
rect 33134 35436 33140 35448
rect 33192 35436 33198 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 20070 35272 20076 35284
rect 20031 35244 20076 35272
rect 20070 35232 20076 35244
rect 20128 35232 20134 35284
rect 20622 35272 20628 35284
rect 20456 35244 20628 35272
rect 20346 35204 20352 35216
rect 19306 35176 20352 35204
rect 18877 35139 18935 35145
rect 18877 35105 18889 35139
rect 18923 35136 18935 35139
rect 19306 35136 19334 35176
rect 20346 35164 20352 35176
rect 20404 35164 20410 35216
rect 20456 35213 20484 35244
rect 20622 35232 20628 35244
rect 20680 35272 20686 35284
rect 21269 35275 21327 35281
rect 21269 35272 21281 35275
rect 20680 35244 21281 35272
rect 20680 35232 20686 35244
rect 21269 35241 21281 35244
rect 21315 35241 21327 35275
rect 21269 35235 21327 35241
rect 21729 35275 21787 35281
rect 21729 35241 21741 35275
rect 21775 35272 21787 35275
rect 22646 35272 22652 35284
rect 21775 35244 22652 35272
rect 21775 35241 21787 35244
rect 21729 35235 21787 35241
rect 22646 35232 22652 35244
rect 22704 35232 22710 35284
rect 23198 35272 23204 35284
rect 23111 35244 23204 35272
rect 23198 35232 23204 35244
rect 23256 35232 23262 35284
rect 24765 35275 24823 35281
rect 24765 35241 24777 35275
rect 24811 35272 24823 35275
rect 25038 35272 25044 35284
rect 24811 35244 25044 35272
rect 24811 35241 24823 35244
rect 24765 35235 24823 35241
rect 25038 35232 25044 35244
rect 25096 35232 25102 35284
rect 30834 35232 30840 35284
rect 30892 35272 30898 35284
rect 31941 35275 31999 35281
rect 31941 35272 31953 35275
rect 30892 35244 31953 35272
rect 30892 35232 30898 35244
rect 31941 35241 31953 35244
rect 31987 35241 31999 35275
rect 31941 35235 31999 35241
rect 20441 35207 20499 35213
rect 20441 35173 20453 35207
rect 20487 35173 20499 35207
rect 20441 35167 20499 35173
rect 20714 35164 20720 35216
rect 20772 35204 20778 35216
rect 23216 35204 23244 35232
rect 20772 35176 23244 35204
rect 20772 35164 20778 35176
rect 22756 35145 22784 35176
rect 29546 35164 29552 35216
rect 29604 35204 29610 35216
rect 29604 35176 35204 35204
rect 29604 35164 29610 35176
rect 22741 35139 22799 35145
rect 18923 35108 19334 35136
rect 20849 35108 22508 35136
rect 18923 35105 18935 35108
rect 18877 35099 18935 35105
rect 20849 35080 20877 35108
rect 22480 35080 22508 35108
rect 22741 35105 22753 35139
rect 22787 35105 22799 35139
rect 23382 35136 23388 35148
rect 22741 35099 22799 35105
rect 23216 35108 23388 35136
rect 18417 35071 18475 35077
rect 18417 35037 18429 35071
rect 18463 35037 18475 35071
rect 18690 35068 18696 35080
rect 18651 35040 18696 35068
rect 18417 35031 18475 35037
rect 18432 35000 18460 35031
rect 18690 35028 18696 35040
rect 18748 35028 18754 35080
rect 20254 35068 20260 35080
rect 20215 35040 20260 35068
rect 20254 35028 20260 35040
rect 20312 35028 20318 35080
rect 20555 35071 20613 35077
rect 20555 35068 20567 35071
rect 20548 35046 20567 35068
rect 20364 35037 20567 35046
rect 20601 35037 20613 35071
rect 20364 35031 20613 35037
rect 20717 35070 20775 35071
rect 20806 35070 20812 35080
rect 20717 35065 20812 35070
rect 20717 35031 20729 35065
rect 20763 35042 20812 35065
rect 20763 35031 20775 35042
rect 20364 35018 20576 35031
rect 20717 35025 20775 35031
rect 20806 35028 20812 35042
rect 20864 35070 20877 35080
rect 20864 35042 20955 35070
rect 21174 35068 21180 35080
rect 20864 35028 20870 35042
rect 21135 35040 21180 35068
rect 21174 35028 21180 35040
rect 21232 35028 21238 35080
rect 21545 35071 21603 35077
rect 21545 35037 21557 35071
rect 21591 35068 21603 35071
rect 21910 35068 21916 35080
rect 21591 35040 21916 35068
rect 21591 35037 21603 35040
rect 21545 35031 21603 35037
rect 19058 35000 19064 35012
rect 18432 34972 19064 35000
rect 19058 34960 19064 34972
rect 19116 35000 19122 35012
rect 20162 35000 20168 35012
rect 19116 34972 20168 35000
rect 19116 34960 19122 34972
rect 20162 34960 20168 34972
rect 20220 34960 20226 35012
rect 20364 35000 20392 35018
rect 20272 34972 20392 35000
rect 20070 34892 20076 34944
rect 20128 34932 20134 34944
rect 20272 34932 20300 34972
rect 20128 34904 20300 34932
rect 20128 34892 20134 34904
rect 20346 34892 20352 34944
rect 20404 34932 20410 34944
rect 21560 34932 21588 35031
rect 21910 35028 21916 35040
rect 21968 35028 21974 35080
rect 22462 35068 22468 35080
rect 22423 35040 22468 35068
rect 22462 35028 22468 35040
rect 22520 35028 22526 35080
rect 22646 35068 22652 35080
rect 22607 35040 22652 35068
rect 22646 35028 22652 35040
rect 22704 35068 22710 35080
rect 23216 35077 23244 35108
rect 23382 35096 23388 35108
rect 23440 35096 23446 35148
rect 27249 35139 27307 35145
rect 27249 35105 27261 35139
rect 27295 35136 27307 35139
rect 28994 35136 29000 35148
rect 27295 35108 29000 35136
rect 27295 35105 27307 35108
rect 27249 35099 27307 35105
rect 28994 35096 29000 35108
rect 29052 35136 29058 35148
rect 30006 35136 30012 35148
rect 29052 35108 30012 35136
rect 29052 35096 29058 35108
rect 30006 35096 30012 35108
rect 30064 35096 30070 35148
rect 30098 35096 30104 35148
rect 30156 35136 30162 35148
rect 30285 35139 30343 35145
rect 30285 35136 30297 35139
rect 30156 35108 30297 35136
rect 30156 35096 30162 35108
rect 30285 35105 30297 35108
rect 30331 35105 30343 35139
rect 30285 35099 30343 35105
rect 23201 35071 23259 35077
rect 23201 35068 23213 35071
rect 22704 35040 23213 35068
rect 22704 35028 22710 35040
rect 23201 35037 23213 35040
rect 23247 35037 23259 35071
rect 23201 35031 23259 35037
rect 23290 35028 23296 35080
rect 23348 35068 23354 35080
rect 23348 35040 23393 35068
rect 23348 35028 23354 35040
rect 23474 35028 23480 35080
rect 23532 35068 23538 35080
rect 24949 35071 25007 35077
rect 24949 35068 24961 35071
rect 23532 35040 24961 35068
rect 23532 35028 23538 35040
rect 24949 35037 24961 35040
rect 24995 35037 25007 35071
rect 24949 35031 25007 35037
rect 25041 35071 25099 35077
rect 25041 35037 25053 35071
rect 25087 35068 25099 35071
rect 25774 35068 25780 35080
rect 25087 35040 25780 35068
rect 25087 35037 25099 35040
rect 25041 35031 25099 35037
rect 22281 35003 22339 35009
rect 22281 34969 22293 35003
rect 22327 35000 22339 35003
rect 24486 35000 24492 35012
rect 22327 34972 24492 35000
rect 22327 34969 22339 34972
rect 22281 34963 22339 34969
rect 24486 34960 24492 34972
rect 24544 34960 24550 35012
rect 24762 35000 24768 35012
rect 24723 34972 24768 35000
rect 24762 34960 24768 34972
rect 24820 34960 24826 35012
rect 24964 35000 24992 35031
rect 25774 35028 25780 35040
rect 25832 35028 25838 35080
rect 26421 35071 26479 35077
rect 26421 35037 26433 35071
rect 26467 35037 26479 35071
rect 26786 35068 26792 35080
rect 26747 35040 26792 35068
rect 26421 35031 26479 35037
rect 26436 35000 26464 35031
rect 26786 35028 26792 35040
rect 26844 35028 26850 35080
rect 29178 35028 29184 35080
rect 29236 35068 29242 35080
rect 30193 35071 30251 35077
rect 30193 35068 30205 35071
rect 29236 35040 30205 35068
rect 29236 35028 29242 35040
rect 30193 35037 30205 35040
rect 30239 35037 30251 35071
rect 32122 35068 32128 35080
rect 32083 35040 32128 35068
rect 30193 35031 30251 35037
rect 32122 35028 32128 35040
rect 32180 35028 32186 35080
rect 32232 35068 32260 35176
rect 32306 35096 32312 35148
rect 32364 35136 32370 35148
rect 32950 35136 32956 35148
rect 32364 35108 32956 35136
rect 32364 35096 32370 35108
rect 32950 35096 32956 35108
rect 33008 35136 33014 35148
rect 33045 35139 33103 35145
rect 33045 35136 33057 35139
rect 33008 35108 33057 35136
rect 33008 35096 33014 35108
rect 33045 35105 33057 35108
rect 33091 35105 33103 35139
rect 33410 35136 33416 35148
rect 33045 35099 33103 35105
rect 33152 35108 33416 35136
rect 32401 35071 32459 35077
rect 32401 35068 32413 35071
rect 32232 35040 32413 35068
rect 32401 35037 32413 35040
rect 32447 35037 32459 35071
rect 32401 35031 32459 35037
rect 32769 35071 32827 35077
rect 32769 35037 32781 35071
rect 32815 35068 32827 35071
rect 33152 35068 33180 35108
rect 33410 35096 33416 35108
rect 33468 35096 33474 35148
rect 34241 35139 34299 35145
rect 34241 35105 34253 35139
rect 34287 35136 34299 35139
rect 35069 35139 35127 35145
rect 35069 35136 35081 35139
rect 34287 35108 35081 35136
rect 34287 35105 34299 35108
rect 34241 35099 34299 35105
rect 35069 35105 35081 35108
rect 35115 35105 35127 35139
rect 35069 35099 35127 35105
rect 32815 35040 33180 35068
rect 33229 35071 33287 35077
rect 32815 35037 32827 35040
rect 32769 35031 32827 35037
rect 33229 35037 33241 35071
rect 33275 35037 33287 35071
rect 33229 35031 33287 35037
rect 24964 34972 26464 35000
rect 29748 34972 30788 35000
rect 20404 34904 21588 34932
rect 20404 34892 20410 34904
rect 22462 34892 22468 34944
rect 22520 34932 22526 34944
rect 23290 34932 23296 34944
rect 22520 34904 23296 34932
rect 22520 34892 22526 34904
rect 23290 34892 23296 34904
rect 23348 34892 23354 34944
rect 23569 34935 23627 34941
rect 23569 34901 23581 34935
rect 23615 34932 23627 34935
rect 24670 34932 24676 34944
rect 23615 34904 24676 34932
rect 23615 34901 23627 34904
rect 23569 34895 23627 34901
rect 24670 34892 24676 34904
rect 24728 34892 24734 34944
rect 29748 34941 29776 34972
rect 29733 34935 29791 34941
rect 29733 34901 29745 34935
rect 29779 34901 29791 34935
rect 29733 34895 29791 34901
rect 30006 34892 30012 34944
rect 30064 34932 30070 34944
rect 30101 34935 30159 34941
rect 30101 34932 30113 34935
rect 30064 34904 30113 34932
rect 30064 34892 30070 34904
rect 30101 34901 30113 34904
rect 30147 34901 30159 34935
rect 30760 34932 30788 34972
rect 30834 34960 30840 35012
rect 30892 35000 30898 35012
rect 32784 35000 32812 35031
rect 30892 34972 32812 35000
rect 30892 34960 30898 34972
rect 33042 34960 33048 35012
rect 33100 35000 33106 35012
rect 33244 35000 33272 35031
rect 34054 35028 34060 35080
rect 34112 35068 34118 35080
rect 35176 35077 35204 35176
rect 34149 35071 34207 35077
rect 34149 35068 34161 35071
rect 34112 35040 34161 35068
rect 34112 35028 34118 35040
rect 34149 35037 34161 35040
rect 34195 35037 34207 35071
rect 34149 35031 34207 35037
rect 34333 35071 34391 35077
rect 34333 35037 34345 35071
rect 34379 35037 34391 35071
rect 34333 35031 34391 35037
rect 35161 35071 35219 35077
rect 35161 35037 35173 35071
rect 35207 35037 35219 35071
rect 35161 35031 35219 35037
rect 33100 34972 33272 35000
rect 33100 34960 33106 34972
rect 33594 34960 33600 35012
rect 33652 35000 33658 35012
rect 34348 35000 34376 35031
rect 33652 34972 34376 35000
rect 33652 34960 33658 34972
rect 32950 34932 32956 34944
rect 30760 34904 32956 34932
rect 30101 34895 30159 34901
rect 32950 34892 32956 34904
rect 33008 34892 33014 34944
rect 35986 34932 35992 34944
rect 35947 34904 35992 34932
rect 35986 34892 35992 34904
rect 36044 34892 36050 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 18785 34731 18843 34737
rect 18785 34697 18797 34731
rect 18831 34728 18843 34731
rect 22646 34728 22652 34740
rect 18831 34700 22652 34728
rect 18831 34697 18843 34700
rect 18785 34691 18843 34697
rect 22646 34688 22652 34700
rect 22704 34688 22710 34740
rect 30009 34731 30067 34737
rect 30009 34697 30021 34731
rect 30055 34728 30067 34731
rect 30374 34728 30380 34740
rect 30055 34700 30380 34728
rect 30055 34697 30067 34700
rect 30009 34691 30067 34697
rect 30374 34688 30380 34700
rect 30432 34688 30438 34740
rect 32585 34731 32643 34737
rect 32585 34697 32597 34731
rect 32631 34728 32643 34731
rect 33226 34728 33232 34740
rect 32631 34700 33232 34728
rect 32631 34697 32643 34700
rect 32585 34691 32643 34697
rect 33226 34688 33232 34700
rect 33284 34688 33290 34740
rect 20070 34620 20076 34672
rect 20128 34660 20134 34672
rect 20128 34632 20852 34660
rect 20128 34620 20134 34632
rect 17402 34592 17408 34604
rect 17363 34564 17408 34592
rect 17402 34552 17408 34564
rect 17460 34552 17466 34604
rect 18138 34592 18144 34604
rect 18099 34564 18144 34592
rect 18138 34552 18144 34564
rect 18196 34552 18202 34604
rect 18233 34595 18291 34601
rect 18233 34561 18245 34595
rect 18279 34561 18291 34595
rect 18233 34555 18291 34561
rect 18785 34595 18843 34601
rect 18785 34561 18797 34595
rect 18831 34592 18843 34595
rect 18874 34592 18880 34604
rect 18831 34564 18880 34592
rect 18831 34561 18843 34564
rect 18785 34555 18843 34561
rect 17218 34484 17224 34536
rect 17276 34524 17282 34536
rect 18248 34524 18276 34555
rect 18874 34552 18880 34564
rect 18932 34552 18938 34604
rect 20254 34592 20260 34604
rect 20167 34564 20260 34592
rect 20254 34552 20260 34564
rect 20312 34552 20318 34604
rect 20346 34552 20352 34604
rect 20404 34592 20410 34604
rect 20404 34564 20449 34592
rect 20404 34552 20410 34564
rect 20622 34552 20628 34604
rect 20680 34592 20686 34604
rect 20717 34595 20775 34601
rect 20717 34592 20729 34595
rect 20680 34564 20729 34592
rect 20680 34552 20686 34564
rect 20717 34561 20729 34564
rect 20763 34561 20775 34595
rect 20824 34592 20852 34632
rect 21174 34620 21180 34672
rect 21232 34660 21238 34672
rect 21232 34632 22232 34660
rect 21232 34620 21238 34632
rect 21358 34592 21364 34604
rect 20824 34564 21364 34592
rect 20717 34555 20775 34561
rect 21358 34552 21364 34564
rect 21416 34552 21422 34604
rect 22002 34592 22008 34604
rect 21963 34564 22008 34592
rect 22002 34552 22008 34564
rect 22060 34552 22066 34604
rect 22204 34601 22232 34632
rect 23750 34620 23756 34672
rect 23808 34620 23814 34672
rect 25038 34660 25044 34672
rect 24596 34632 25044 34660
rect 22189 34595 22247 34601
rect 22189 34561 22201 34595
rect 22235 34561 22247 34595
rect 23768 34592 23796 34620
rect 23950 34597 24008 34603
rect 23950 34594 23962 34597
rect 23860 34592 23962 34594
rect 23768 34566 23962 34592
rect 23768 34564 23888 34566
rect 22189 34555 22247 34561
rect 23950 34563 23962 34566
rect 23996 34563 24008 34597
rect 24210 34592 24216 34604
rect 24171 34564 24216 34592
rect 23950 34557 24008 34563
rect 24210 34552 24216 34564
rect 24268 34552 24274 34604
rect 24305 34595 24363 34601
rect 24305 34561 24317 34595
rect 24351 34592 24363 34595
rect 24486 34592 24492 34604
rect 24351 34564 24492 34592
rect 24351 34561 24363 34564
rect 24305 34555 24363 34561
rect 24486 34552 24492 34564
rect 24544 34552 24550 34604
rect 24596 34601 24624 34632
rect 25038 34620 25044 34632
rect 25096 34660 25102 34672
rect 25096 34632 25636 34660
rect 25096 34620 25102 34632
rect 24581 34595 24639 34601
rect 24581 34561 24593 34595
rect 24627 34561 24639 34595
rect 24581 34555 24639 34561
rect 24670 34552 24676 34604
rect 24728 34592 24734 34604
rect 25608 34601 25636 34632
rect 32398 34620 32404 34672
rect 32456 34660 32462 34672
rect 33042 34660 33048 34672
rect 32456 34632 33048 34660
rect 32456 34620 32462 34632
rect 33042 34620 33048 34632
rect 33100 34660 33106 34672
rect 33100 34632 33548 34660
rect 33100 34620 33106 34632
rect 24765 34595 24823 34601
rect 24765 34592 24777 34595
rect 24728 34564 24777 34592
rect 24728 34552 24734 34564
rect 24765 34561 24777 34564
rect 24811 34561 24823 34595
rect 24765 34555 24823 34561
rect 25593 34595 25651 34601
rect 25593 34561 25605 34595
rect 25639 34561 25651 34595
rect 25593 34555 25651 34561
rect 29546 34552 29552 34604
rect 29604 34592 29610 34604
rect 29825 34595 29883 34601
rect 29825 34592 29837 34595
rect 29604 34564 29837 34592
rect 29604 34552 29610 34564
rect 29825 34561 29837 34564
rect 29871 34561 29883 34595
rect 29825 34555 29883 34561
rect 30009 34595 30067 34601
rect 30009 34561 30021 34595
rect 30055 34592 30067 34595
rect 30834 34592 30840 34604
rect 30055 34564 30840 34592
rect 30055 34561 30067 34564
rect 30009 34555 30067 34561
rect 30834 34552 30840 34564
rect 30892 34552 30898 34604
rect 32306 34592 32312 34604
rect 32267 34564 32312 34592
rect 32306 34552 32312 34564
rect 32364 34552 32370 34604
rect 33134 34592 33140 34604
rect 33095 34564 33140 34592
rect 33134 34552 33140 34564
rect 33192 34552 33198 34604
rect 33520 34601 33548 34632
rect 33505 34595 33563 34601
rect 33505 34561 33517 34595
rect 33551 34561 33563 34595
rect 33505 34555 33563 34561
rect 17276 34496 18276 34524
rect 20272 34524 20300 34552
rect 20272 34496 22048 34524
rect 17276 34484 17282 34496
rect 22020 34456 22048 34496
rect 22094 34484 22100 34536
rect 22152 34524 22158 34536
rect 22152 34496 23244 34524
rect 22152 34484 22158 34496
rect 22186 34456 22192 34468
rect 22020 34428 22192 34456
rect 22186 34416 22192 34428
rect 22244 34456 22250 34468
rect 22373 34459 22431 34465
rect 22373 34456 22385 34459
rect 22244 34428 22385 34456
rect 22244 34416 22250 34428
rect 22373 34425 22385 34428
rect 22419 34425 22431 34459
rect 23216 34456 23244 34496
rect 23290 34484 23296 34536
rect 23348 34524 23354 34536
rect 25409 34527 25467 34533
rect 25409 34524 25421 34527
rect 23348 34496 25421 34524
rect 23348 34484 23354 34496
rect 25409 34493 25421 34496
rect 25455 34493 25467 34527
rect 25409 34487 25467 34493
rect 25777 34527 25835 34533
rect 25777 34493 25789 34527
rect 25823 34524 25835 34527
rect 26418 34524 26424 34536
rect 25823 34496 26424 34524
rect 25823 34493 25835 34496
rect 25777 34487 25835 34493
rect 26418 34484 26424 34496
rect 26476 34484 26482 34536
rect 32122 34484 32128 34536
rect 32180 34524 32186 34536
rect 32585 34527 32643 34533
rect 32585 34524 32597 34527
rect 32180 34496 32597 34524
rect 32180 34484 32186 34496
rect 32585 34493 32597 34496
rect 32631 34524 32643 34527
rect 32766 34524 32772 34536
rect 32631 34496 32772 34524
rect 32631 34493 32643 34496
rect 32585 34487 32643 34493
rect 32766 34484 32772 34496
rect 32824 34484 32830 34536
rect 24210 34456 24216 34468
rect 23216 34428 24216 34456
rect 22373 34419 22431 34425
rect 24210 34416 24216 34428
rect 24268 34416 24274 34468
rect 33870 34416 33876 34468
rect 33928 34456 33934 34468
rect 34333 34459 34391 34465
rect 34333 34456 34345 34459
rect 33928 34428 34345 34456
rect 33928 34416 33934 34428
rect 34333 34425 34345 34428
rect 34379 34425 34391 34459
rect 34333 34419 34391 34425
rect 21453 34391 21511 34397
rect 21453 34357 21465 34391
rect 21499 34388 21511 34391
rect 21542 34388 21548 34400
rect 21499 34360 21548 34388
rect 21499 34357 21511 34360
rect 21453 34351 21511 34357
rect 21542 34348 21548 34360
rect 21600 34348 21606 34400
rect 23569 34391 23627 34397
rect 23569 34357 23581 34391
rect 23615 34388 23627 34391
rect 25682 34388 25688 34400
rect 23615 34360 25688 34388
rect 23615 34357 23627 34360
rect 23569 34351 23627 34357
rect 25682 34348 25688 34360
rect 25740 34348 25746 34400
rect 32398 34388 32404 34400
rect 32359 34360 32404 34388
rect 32398 34348 32404 34360
rect 32456 34348 32462 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 16945 34187 17003 34193
rect 16945 34153 16957 34187
rect 16991 34184 17003 34187
rect 20714 34184 20720 34196
rect 16991 34156 20720 34184
rect 16991 34153 17003 34156
rect 16945 34147 17003 34153
rect 20714 34144 20720 34156
rect 20772 34144 20778 34196
rect 32766 34184 32772 34196
rect 32727 34156 32772 34184
rect 32766 34144 32772 34156
rect 32824 34144 32830 34196
rect 18874 34116 18880 34128
rect 17972 34088 18880 34116
rect 17313 34051 17371 34057
rect 17313 34017 17325 34051
rect 17359 34048 17371 34051
rect 17972 34048 18000 34088
rect 18874 34076 18880 34088
rect 18932 34116 18938 34128
rect 21542 34116 21548 34128
rect 18932 34088 21548 34116
rect 18932 34076 18938 34088
rect 21542 34076 21548 34088
rect 21600 34076 21606 34128
rect 26786 34116 26792 34128
rect 26747 34088 26792 34116
rect 26786 34076 26792 34088
rect 26844 34076 26850 34128
rect 17359 34020 18000 34048
rect 17359 34017 17371 34020
rect 17313 34011 17371 34017
rect 17129 33983 17187 33989
rect 17129 33949 17141 33983
rect 17175 33949 17187 33983
rect 17129 33943 17187 33949
rect 17144 33912 17172 33943
rect 17218 33940 17224 33992
rect 17276 33980 17282 33992
rect 17276 33952 17321 33980
rect 17276 33940 17282 33952
rect 17402 33940 17408 33992
rect 17460 33980 17466 33992
rect 17972 33989 18000 34020
rect 18693 34051 18751 34057
rect 18693 34017 18705 34051
rect 18739 34048 18751 34051
rect 18782 34048 18788 34060
rect 18739 34020 18788 34048
rect 18739 34017 18751 34020
rect 18693 34011 18751 34017
rect 18782 34008 18788 34020
rect 18840 34008 18846 34060
rect 20622 34008 20628 34060
rect 20680 34048 20686 34060
rect 20680 34020 21680 34048
rect 20680 34008 20686 34020
rect 17957 33983 18015 33989
rect 17460 33952 17505 33980
rect 17460 33940 17466 33952
rect 17957 33949 17969 33983
rect 18003 33949 18015 33983
rect 17957 33943 18015 33949
rect 18046 33940 18052 33992
rect 18104 33980 18110 33992
rect 18233 33983 18291 33989
rect 18104 33952 18149 33980
rect 18104 33940 18110 33952
rect 18233 33949 18245 33983
rect 18279 33949 18291 33983
rect 18233 33943 18291 33949
rect 18138 33912 18144 33924
rect 17144 33884 18144 33912
rect 18138 33872 18144 33884
rect 18196 33912 18202 33924
rect 18248 33912 18276 33943
rect 18322 33940 18328 33992
rect 18380 33980 18386 33992
rect 21177 33983 21235 33989
rect 21177 33980 21189 33983
rect 18380 33952 21189 33980
rect 18380 33940 18386 33952
rect 21177 33949 21189 33952
rect 21223 33949 21235 33983
rect 21358 33980 21364 33992
rect 21319 33952 21364 33980
rect 21177 33943 21235 33949
rect 21358 33940 21364 33952
rect 21416 33940 21422 33992
rect 21652 33989 21680 34020
rect 24762 34008 24768 34060
rect 24820 34048 24826 34060
rect 24820 34020 26174 34048
rect 24820 34008 24826 34020
rect 21637 33983 21695 33989
rect 21637 33949 21649 33983
rect 21683 33949 21695 33983
rect 21910 33980 21916 33992
rect 21871 33952 21916 33980
rect 21637 33943 21695 33949
rect 21910 33940 21916 33952
rect 21968 33940 21974 33992
rect 22186 33980 22192 33992
rect 22147 33952 22192 33980
rect 22186 33940 22192 33952
rect 22244 33940 22250 33992
rect 24946 33940 24952 33992
rect 25004 33980 25010 33992
rect 25409 33983 25467 33989
rect 25409 33980 25421 33983
rect 25004 33952 25421 33980
rect 25004 33940 25010 33952
rect 25409 33949 25421 33952
rect 25455 33949 25467 33983
rect 25409 33943 25467 33949
rect 18196 33884 18276 33912
rect 20809 33915 20867 33921
rect 18196 33872 18202 33884
rect 20809 33881 20821 33915
rect 20855 33912 20867 33915
rect 23014 33912 23020 33924
rect 20855 33884 23020 33912
rect 20855 33881 20867 33884
rect 20809 33875 20867 33881
rect 23014 33872 23020 33884
rect 23072 33872 23078 33924
rect 25424 33912 25452 33943
rect 25682 33940 25688 33992
rect 25740 33980 25746 33992
rect 25777 33983 25835 33989
rect 25777 33980 25789 33983
rect 25740 33952 25789 33980
rect 25740 33940 25746 33952
rect 25777 33949 25789 33952
rect 25823 33980 25835 33983
rect 26418 33980 26424 33992
rect 25823 33952 26280 33980
rect 26379 33952 26424 33980
rect 25823 33949 25835 33952
rect 25777 33943 25835 33949
rect 26142 33912 26148 33924
rect 25424 33884 26148 33912
rect 26142 33872 26148 33884
rect 26200 33872 26206 33924
rect 26252 33912 26280 33952
rect 26418 33940 26424 33952
rect 26476 33940 26482 33992
rect 31662 33940 31668 33992
rect 31720 33980 31726 33992
rect 32677 33983 32735 33989
rect 32677 33980 32689 33983
rect 31720 33952 32689 33980
rect 31720 33940 31726 33952
rect 32677 33949 32689 33952
rect 32723 33949 32735 33983
rect 32677 33943 32735 33949
rect 27246 33912 27252 33924
rect 26252 33884 27252 33912
rect 27246 33872 27252 33884
rect 27304 33872 27310 33924
rect 32490 33912 32496 33924
rect 32451 33884 32496 33912
rect 32490 33872 32496 33884
rect 32548 33872 32554 33924
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 25038 33640 25044 33652
rect 16132 33612 17632 33640
rect 24999 33612 25044 33640
rect 16025 33507 16083 33513
rect 16025 33473 16037 33507
rect 16071 33504 16083 33507
rect 16132 33504 16160 33612
rect 16301 33575 16359 33581
rect 16301 33541 16313 33575
rect 16347 33572 16359 33575
rect 17402 33572 17408 33584
rect 16347 33544 17408 33572
rect 16347 33541 16359 33544
rect 16301 33535 16359 33541
rect 17402 33532 17408 33544
rect 17460 33532 17466 33584
rect 17604 33516 17632 33612
rect 25038 33600 25044 33612
rect 25096 33600 25102 33652
rect 32306 33600 32312 33652
rect 32364 33640 32370 33652
rect 32769 33643 32827 33649
rect 32769 33640 32781 33643
rect 32364 33612 32781 33640
rect 32364 33600 32370 33612
rect 32769 33609 32781 33612
rect 32815 33609 32827 33643
rect 32769 33603 32827 33609
rect 18690 33532 18696 33584
rect 18748 33572 18754 33584
rect 19429 33575 19487 33581
rect 18748 33544 18920 33572
rect 18748 33532 18754 33544
rect 16071 33476 16160 33504
rect 16209 33507 16267 33513
rect 16071 33473 16083 33476
rect 16025 33467 16083 33473
rect 16209 33473 16221 33507
rect 16255 33504 16267 33507
rect 17218 33504 17224 33516
rect 16255 33476 16988 33504
rect 17179 33476 17224 33504
rect 16255 33473 16267 33476
rect 16209 33467 16267 33473
rect 16960 33368 16988 33476
rect 17218 33464 17224 33476
rect 17276 33464 17282 33516
rect 17494 33504 17500 33516
rect 17455 33476 17500 33504
rect 17494 33464 17500 33476
rect 17552 33464 17558 33516
rect 17586 33464 17592 33516
rect 17644 33504 17650 33516
rect 17681 33507 17739 33513
rect 17681 33504 17693 33507
rect 17644 33476 17693 33504
rect 17644 33464 17650 33476
rect 17681 33473 17693 33476
rect 17727 33473 17739 33507
rect 18046 33504 18052 33516
rect 17681 33467 17739 33473
rect 17788 33476 18052 33504
rect 17037 33439 17095 33445
rect 17037 33405 17049 33439
rect 17083 33436 17095 33439
rect 17788 33436 17816 33476
rect 18046 33464 18052 33476
rect 18104 33504 18110 33516
rect 18892 33513 18920 33544
rect 19429 33541 19441 33575
rect 19475 33572 19487 33575
rect 20622 33572 20628 33584
rect 19475 33544 20628 33572
rect 19475 33541 19487 33544
rect 19429 33535 19487 33541
rect 20622 33532 20628 33544
rect 20680 33532 20686 33584
rect 18325 33507 18383 33513
rect 18325 33504 18337 33507
rect 18104 33476 18337 33504
rect 18104 33464 18110 33476
rect 18325 33473 18337 33476
rect 18371 33473 18383 33507
rect 18325 33467 18383 33473
rect 18877 33507 18935 33513
rect 18877 33473 18889 33507
rect 18923 33473 18935 33507
rect 19058 33504 19064 33516
rect 19019 33476 19064 33504
rect 18877 33467 18935 33473
rect 19058 33464 19064 33476
rect 19116 33464 19122 33516
rect 25041 33507 25099 33513
rect 25041 33473 25053 33507
rect 25087 33504 25099 33507
rect 26418 33504 26424 33516
rect 25087 33476 26424 33504
rect 25087 33473 25099 33476
rect 25041 33467 25099 33473
rect 26418 33464 26424 33476
rect 26476 33464 26482 33516
rect 27341 33507 27399 33513
rect 27341 33473 27353 33507
rect 27387 33473 27399 33507
rect 27890 33504 27896 33516
rect 27851 33476 27896 33504
rect 27341 33467 27399 33473
rect 18138 33436 18144 33448
rect 17083 33408 17816 33436
rect 18099 33408 18144 33436
rect 17083 33405 17095 33408
rect 17037 33399 17095 33405
rect 18138 33396 18144 33408
rect 18196 33396 18202 33448
rect 24857 33439 24915 33445
rect 24857 33405 24869 33439
rect 24903 33405 24915 33439
rect 25406 33436 25412 33448
rect 25367 33408 25412 33436
rect 24857 33399 24915 33405
rect 17494 33368 17500 33380
rect 16960 33340 17500 33368
rect 17494 33328 17500 33340
rect 17552 33328 17558 33380
rect 24872 33368 24900 33399
rect 25406 33396 25412 33408
rect 25464 33396 25470 33448
rect 25958 33396 25964 33448
rect 26016 33436 26022 33448
rect 27356 33436 27384 33467
rect 27890 33464 27896 33476
rect 27948 33464 27954 33516
rect 28828 33504 28856 33558
rect 28902 33532 28908 33584
rect 28960 33572 28966 33584
rect 31573 33575 31631 33581
rect 28960 33544 30144 33572
rect 28960 33532 28966 33544
rect 29546 33504 29552 33516
rect 28828 33476 29552 33504
rect 29546 33464 29552 33476
rect 29604 33464 29610 33516
rect 29730 33504 29736 33516
rect 29691 33476 29736 33504
rect 29730 33464 29736 33476
rect 29788 33464 29794 33516
rect 30116 33513 30144 33544
rect 31573 33541 31585 33575
rect 31619 33572 31631 33575
rect 32398 33572 32404 33584
rect 31619 33544 32404 33572
rect 31619 33541 31631 33544
rect 31573 33535 31631 33541
rect 32398 33532 32404 33544
rect 32456 33532 32462 33584
rect 30101 33507 30159 33513
rect 30101 33473 30113 33507
rect 30147 33473 30159 33507
rect 30101 33467 30159 33473
rect 32490 33464 32496 33516
rect 32548 33504 32554 33516
rect 32585 33507 32643 33513
rect 32585 33504 32597 33507
rect 32548 33476 32597 33504
rect 32548 33464 32554 33476
rect 32585 33473 32597 33476
rect 32631 33473 32643 33507
rect 32585 33467 32643 33473
rect 26016 33408 27384 33436
rect 26016 33396 26022 33408
rect 31662 33396 31668 33448
rect 31720 33436 31726 33448
rect 32401 33439 32459 33445
rect 32401 33436 32413 33439
rect 31720 33408 32413 33436
rect 31720 33396 31726 33408
rect 32401 33405 32413 33408
rect 32447 33405 32459 33439
rect 32401 33399 32459 33405
rect 24946 33368 24952 33380
rect 24859 33340 24952 33368
rect 24946 33328 24952 33340
rect 25004 33368 25010 33380
rect 25976 33368 26004 33396
rect 25004 33340 26004 33368
rect 25004 33328 25010 33340
rect 26513 33303 26571 33309
rect 26513 33269 26525 33303
rect 26559 33300 26571 33303
rect 27430 33300 27436 33312
rect 26559 33272 27436 33300
rect 26559 33269 26571 33272
rect 26513 33263 26571 33269
rect 27430 33260 27436 33272
rect 27488 33260 27494 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 16945 33099 17003 33105
rect 16945 33065 16957 33099
rect 16991 33096 17003 33099
rect 17218 33096 17224 33108
rect 16991 33068 17224 33096
rect 16991 33065 17003 33068
rect 16945 33059 17003 33065
rect 17218 33056 17224 33068
rect 17276 33056 17282 33108
rect 24673 33099 24731 33105
rect 24673 33065 24685 33099
rect 24719 33096 24731 33099
rect 24762 33096 24768 33108
rect 24719 33068 24768 33096
rect 24719 33065 24731 33068
rect 24673 33059 24731 33065
rect 24762 33056 24768 33068
rect 24820 33056 24826 33108
rect 25774 33096 25780 33108
rect 25735 33068 25780 33096
rect 25774 33056 25780 33068
rect 25832 33056 25838 33108
rect 26973 33099 27031 33105
rect 26973 33065 26985 33099
rect 27019 33096 27031 33099
rect 27890 33096 27896 33108
rect 27019 33068 27896 33096
rect 27019 33065 27031 33068
rect 26973 33059 27031 33065
rect 27890 33056 27896 33068
rect 27948 33056 27954 33108
rect 19334 33028 19340 33040
rect 17880 33000 19340 33028
rect 16577 32963 16635 32969
rect 16577 32929 16589 32963
rect 16623 32960 16635 32963
rect 17880 32960 17908 33000
rect 19334 32988 19340 33000
rect 19392 32988 19398 33040
rect 23106 32988 23112 33040
rect 23164 33028 23170 33040
rect 23385 33031 23443 33037
rect 23385 33028 23397 33031
rect 23164 33000 23397 33028
rect 23164 32988 23170 33000
rect 23385 32997 23397 33000
rect 23431 32997 23443 33031
rect 23385 32991 23443 32997
rect 24949 33031 25007 33037
rect 24949 32997 24961 33031
rect 24995 33028 25007 33031
rect 25406 33028 25412 33040
rect 24995 33000 25412 33028
rect 24995 32997 25007 33000
rect 24949 32991 25007 32997
rect 25406 32988 25412 33000
rect 25464 33028 25470 33040
rect 26142 33028 26148 33040
rect 25464 33000 26148 33028
rect 25464 32988 25470 33000
rect 26142 32988 26148 33000
rect 26200 32988 26206 33040
rect 26234 32988 26240 33040
rect 26292 33028 26298 33040
rect 28353 33031 28411 33037
rect 26292 33000 26832 33028
rect 26292 32988 26298 33000
rect 18138 32960 18144 32972
rect 16623 32932 17908 32960
rect 18099 32932 18144 32960
rect 16623 32929 16635 32932
rect 16577 32923 16635 32929
rect 16761 32895 16819 32901
rect 16761 32861 16773 32895
rect 16807 32861 16819 32895
rect 16761 32855 16819 32861
rect 17773 32895 17831 32901
rect 17773 32861 17785 32895
rect 17819 32892 17831 32895
rect 17880 32892 17908 32932
rect 18138 32920 18144 32932
rect 18196 32920 18202 32972
rect 23569 32963 23627 32969
rect 23569 32929 23581 32963
rect 23615 32960 23627 32963
rect 25041 32963 25099 32969
rect 25041 32960 25053 32963
rect 23615 32932 25053 32960
rect 23615 32929 23627 32932
rect 23569 32923 23627 32929
rect 25041 32929 25053 32932
rect 25087 32929 25099 32963
rect 25041 32923 25099 32929
rect 25332 32932 26464 32960
rect 25332 32904 25360 32932
rect 17819 32864 17908 32892
rect 17957 32895 18015 32901
rect 17819 32861 17831 32864
rect 17773 32855 17831 32861
rect 17957 32861 17969 32895
rect 18003 32861 18015 32895
rect 17957 32855 18015 32861
rect 16776 32824 16804 32855
rect 17678 32824 17684 32836
rect 16776 32796 17684 32824
rect 17678 32784 17684 32796
rect 17736 32824 17742 32836
rect 17972 32824 18000 32855
rect 23014 32852 23020 32904
rect 23072 32892 23078 32904
rect 23109 32895 23167 32901
rect 23109 32892 23121 32895
rect 23072 32864 23121 32892
rect 23072 32852 23078 32864
rect 23109 32861 23121 32864
rect 23155 32861 23167 32895
rect 24854 32892 24860 32904
rect 24815 32864 24860 32892
rect 23109 32855 23167 32861
rect 24854 32852 24860 32864
rect 24912 32852 24918 32904
rect 25133 32895 25191 32901
rect 25133 32861 25145 32895
rect 25179 32861 25191 32895
rect 25314 32892 25320 32904
rect 25275 32864 25320 32892
rect 25133 32855 25191 32861
rect 17736 32796 18000 32824
rect 25148 32824 25176 32855
rect 25314 32852 25320 32864
rect 25372 32852 25378 32904
rect 25958 32892 25964 32904
rect 25919 32864 25964 32892
rect 25958 32852 25964 32864
rect 26016 32852 26022 32904
rect 26053 32895 26111 32901
rect 26053 32861 26065 32895
rect 26099 32861 26111 32895
rect 26053 32855 26111 32861
rect 26068 32824 26096 32855
rect 26142 32852 26148 32904
rect 26200 32892 26206 32904
rect 26436 32902 26464 32932
rect 26344 32901 26464 32902
rect 26237 32895 26295 32901
rect 26237 32892 26249 32895
rect 26200 32864 26249 32892
rect 26200 32852 26206 32864
rect 26237 32861 26249 32864
rect 26283 32861 26295 32895
rect 26237 32855 26295 32861
rect 26329 32895 26464 32901
rect 26329 32861 26341 32895
rect 26375 32874 26464 32895
rect 26804 32892 26832 33000
rect 28353 32997 28365 33031
rect 28399 33028 28411 33031
rect 29730 33028 29736 33040
rect 28399 33000 29736 33028
rect 28399 32997 28411 33000
rect 28353 32991 28411 32997
rect 29730 32988 29736 33000
rect 29788 32988 29794 33040
rect 27154 32892 27160 32904
rect 26375 32861 26387 32874
rect 26804 32864 27160 32892
rect 26329 32855 26387 32861
rect 27154 32852 27160 32864
rect 27212 32852 27218 32904
rect 27246 32852 27252 32904
rect 27304 32892 27310 32904
rect 27430 32892 27436 32904
rect 27304 32864 27349 32892
rect 27391 32864 27436 32892
rect 27304 32852 27310 32864
rect 27430 32852 27436 32864
rect 27488 32852 27494 32904
rect 27522 32852 27528 32904
rect 27580 32892 27586 32904
rect 28074 32892 28080 32904
rect 27580 32864 27625 32892
rect 28035 32864 28080 32892
rect 27580 32852 27586 32864
rect 28074 32852 28080 32864
rect 28132 32852 28138 32904
rect 28626 32892 28632 32904
rect 28587 32864 28632 32892
rect 28626 32852 28632 32864
rect 28684 32852 28690 32904
rect 28905 32895 28963 32901
rect 28905 32861 28917 32895
rect 28951 32861 28963 32895
rect 28905 32855 28963 32861
rect 26418 32824 26424 32836
rect 25148 32796 26424 32824
rect 17736 32784 17742 32796
rect 26418 32784 26424 32796
rect 26476 32784 26482 32836
rect 27172 32824 27200 32852
rect 28920 32824 28948 32855
rect 27172 32796 28948 32824
rect 21266 32716 21272 32768
rect 21324 32756 21330 32768
rect 22002 32756 22008 32768
rect 21324 32728 22008 32756
rect 21324 32716 21330 32728
rect 22002 32716 22008 32728
rect 22060 32716 22066 32768
rect 27246 32716 27252 32768
rect 27304 32756 27310 32768
rect 27798 32756 27804 32768
rect 27304 32728 27804 32756
rect 27304 32716 27310 32728
rect 27798 32716 27804 32728
rect 27856 32756 27862 32768
rect 28626 32756 28632 32768
rect 27856 32728 28632 32756
rect 27856 32716 27862 32728
rect 28626 32716 28632 32728
rect 28684 32716 28690 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 17494 32552 17500 32564
rect 17455 32524 17500 32552
rect 17494 32512 17500 32524
rect 17552 32512 17558 32564
rect 17586 32512 17592 32564
rect 17644 32552 17650 32564
rect 18693 32555 18751 32561
rect 18693 32552 18705 32555
rect 17644 32524 18705 32552
rect 17644 32512 17650 32524
rect 18693 32521 18705 32524
rect 18739 32521 18751 32555
rect 18693 32515 18751 32521
rect 26142 32512 26148 32564
rect 26200 32552 26206 32564
rect 27522 32552 27528 32564
rect 26200 32524 27528 32552
rect 26200 32512 26206 32524
rect 27522 32512 27528 32524
rect 27580 32552 27586 32564
rect 28077 32555 28135 32561
rect 28077 32552 28089 32555
rect 27580 32524 28089 32552
rect 27580 32512 27586 32524
rect 28077 32521 28089 32524
rect 28123 32521 28135 32555
rect 34422 32552 34428 32564
rect 28077 32515 28135 32521
rect 33888 32524 34428 32552
rect 18322 32484 18328 32496
rect 17512 32456 18328 32484
rect 17512 32425 17540 32456
rect 18322 32444 18328 32456
rect 18380 32444 18386 32496
rect 18541 32487 18599 32493
rect 18541 32484 18553 32487
rect 18432 32456 18553 32484
rect 17497 32419 17555 32425
rect 17497 32385 17509 32419
rect 17543 32385 17555 32419
rect 18432 32416 18460 32456
rect 18541 32453 18553 32456
rect 18587 32484 18599 32487
rect 18874 32484 18880 32496
rect 18587 32456 18880 32484
rect 18587 32453 18599 32456
rect 18541 32447 18599 32453
rect 18874 32444 18880 32456
rect 18932 32444 18938 32496
rect 21085 32487 21143 32493
rect 21085 32453 21097 32487
rect 21131 32484 21143 32487
rect 21358 32484 21364 32496
rect 21131 32456 21364 32484
rect 21131 32453 21143 32456
rect 21085 32447 21143 32453
rect 21358 32444 21364 32456
rect 21416 32444 21422 32496
rect 23014 32444 23020 32496
rect 23072 32484 23078 32496
rect 23382 32484 23388 32496
rect 23072 32456 23388 32484
rect 23072 32444 23078 32456
rect 23382 32444 23388 32456
rect 23440 32484 23446 32496
rect 24946 32484 24952 32496
rect 23440 32456 23520 32484
rect 24426 32456 24952 32484
rect 23440 32444 23446 32456
rect 20806 32416 20812 32428
rect 17497 32379 17555 32385
rect 17604 32388 18460 32416
rect 20767 32388 20812 32416
rect 17313 32351 17371 32357
rect 17313 32317 17325 32351
rect 17359 32348 17371 32351
rect 17604 32348 17632 32388
rect 20806 32376 20812 32388
rect 20864 32376 20870 32428
rect 20993 32419 21051 32425
rect 20993 32385 21005 32419
rect 21039 32416 21051 32419
rect 21266 32416 21272 32428
rect 21039 32388 21272 32416
rect 21039 32385 21051 32388
rect 20993 32379 21051 32385
rect 21266 32376 21272 32388
rect 21324 32376 21330 32428
rect 23106 32416 23112 32428
rect 23067 32388 23112 32416
rect 23106 32376 23112 32388
rect 23164 32376 23170 32428
rect 23492 32425 23520 32456
rect 24946 32444 24952 32456
rect 25004 32444 25010 32496
rect 28905 32487 28963 32493
rect 28905 32484 28917 32487
rect 27264 32456 28917 32484
rect 27264 32425 27292 32456
rect 23477 32419 23535 32425
rect 23477 32385 23489 32419
rect 23523 32385 23535 32419
rect 23477 32379 23535 32385
rect 27249 32419 27307 32425
rect 27249 32385 27261 32419
rect 27295 32385 27307 32419
rect 27249 32379 27307 32385
rect 27338 32376 27344 32428
rect 27396 32416 27402 32428
rect 28276 32425 28304 32456
rect 28905 32453 28917 32456
rect 28951 32453 28963 32487
rect 28905 32447 28963 32453
rect 27985 32419 28043 32425
rect 27985 32416 27997 32419
rect 27396 32388 27997 32416
rect 27396 32376 27402 32388
rect 27985 32385 27997 32388
rect 28031 32385 28043 32419
rect 27985 32379 28043 32385
rect 28261 32419 28319 32425
rect 28261 32385 28273 32419
rect 28307 32385 28319 32419
rect 28810 32416 28816 32428
rect 28771 32388 28816 32416
rect 28261 32379 28319 32385
rect 17862 32348 17868 32360
rect 17359 32320 17632 32348
rect 17823 32320 17868 32348
rect 17359 32317 17371 32320
rect 17313 32311 17371 32317
rect 17862 32308 17868 32320
rect 17920 32308 17926 32360
rect 18322 32308 18328 32360
rect 18380 32348 18386 32360
rect 19150 32348 19156 32360
rect 18380 32320 19156 32348
rect 18380 32308 18386 32320
rect 19150 32308 19156 32320
rect 19208 32308 19214 32360
rect 26418 32240 26424 32292
rect 26476 32280 26482 32292
rect 27249 32283 27307 32289
rect 27249 32280 27261 32283
rect 26476 32252 27261 32280
rect 26476 32240 26482 32252
rect 27249 32249 27261 32252
rect 27295 32249 27307 32283
rect 28000 32280 28028 32379
rect 28810 32376 28816 32388
rect 28868 32376 28874 32428
rect 28997 32419 29055 32425
rect 28997 32416 29009 32419
rect 28920 32388 29009 32416
rect 28350 32308 28356 32360
rect 28408 32348 28414 32360
rect 28920 32348 28948 32388
rect 28997 32385 29009 32388
rect 29043 32385 29055 32419
rect 28997 32379 29055 32385
rect 29638 32376 29644 32428
rect 29696 32416 29702 32428
rect 33888 32425 33916 32524
rect 34422 32512 34428 32524
rect 34480 32512 34486 32564
rect 34149 32487 34207 32493
rect 34149 32453 34161 32487
rect 34195 32484 34207 32487
rect 34514 32484 34520 32496
rect 34195 32456 34520 32484
rect 34195 32453 34207 32456
rect 34149 32447 34207 32453
rect 34514 32444 34520 32456
rect 34572 32444 34578 32496
rect 34716 32456 35296 32484
rect 33873 32419 33931 32425
rect 33873 32416 33885 32419
rect 29696 32388 33885 32416
rect 29696 32376 29702 32388
rect 33873 32385 33885 32388
rect 33919 32385 33931 32419
rect 34609 32419 34667 32425
rect 34609 32416 34621 32419
rect 33873 32379 33931 32385
rect 34164 32388 34621 32416
rect 28408 32320 28948 32348
rect 28408 32308 28414 32320
rect 32950 32308 32956 32360
rect 33008 32348 33014 32360
rect 34164 32357 34192 32388
rect 34609 32385 34621 32388
rect 34655 32385 34667 32419
rect 34609 32379 34667 32385
rect 34149 32351 34207 32357
rect 34149 32348 34161 32351
rect 33008 32320 34161 32348
rect 33008 32308 33014 32320
rect 34149 32317 34161 32320
rect 34195 32317 34207 32351
rect 34716 32348 34744 32456
rect 35268 32425 35296 32456
rect 34793 32419 34851 32425
rect 34793 32385 34805 32419
rect 34839 32385 34851 32419
rect 34793 32379 34851 32385
rect 35253 32419 35311 32425
rect 35253 32385 35265 32419
rect 35299 32416 35311 32419
rect 35986 32416 35992 32428
rect 35299 32388 35992 32416
rect 35299 32385 35311 32388
rect 35253 32379 35311 32385
rect 34149 32311 34207 32317
rect 34440 32320 34744 32348
rect 34808 32348 34836 32379
rect 35986 32376 35992 32388
rect 36044 32376 36050 32428
rect 35342 32348 35348 32360
rect 34808 32320 35348 32348
rect 31662 32280 31668 32292
rect 28000 32252 31668 32280
rect 27249 32243 27307 32249
rect 31662 32240 31668 32252
rect 31720 32240 31726 32292
rect 17862 32172 17868 32224
rect 17920 32212 17926 32224
rect 18509 32215 18567 32221
rect 18509 32212 18521 32215
rect 17920 32184 18521 32212
rect 17920 32172 17926 32184
rect 18509 32181 18521 32184
rect 18555 32181 18567 32215
rect 18509 32175 18567 32181
rect 33502 32172 33508 32224
rect 33560 32212 33566 32224
rect 33965 32215 34023 32221
rect 33965 32212 33977 32215
rect 33560 32184 33977 32212
rect 33560 32172 33566 32184
rect 33965 32181 33977 32184
rect 34011 32212 34023 32215
rect 34440 32212 34468 32320
rect 35342 32308 35348 32320
rect 35400 32308 35406 32360
rect 34606 32212 34612 32224
rect 34011 32184 34468 32212
rect 34567 32184 34612 32212
rect 34011 32181 34023 32184
rect 33965 32175 34023 32181
rect 34606 32172 34612 32184
rect 34664 32172 34670 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 17586 31968 17592 32020
rect 17644 32008 17650 32020
rect 23198 32008 23204 32020
rect 17644 31980 23204 32008
rect 17644 31968 17650 31980
rect 23198 31968 23204 31980
rect 23256 32008 23262 32020
rect 23569 32011 23627 32017
rect 23256 31980 23520 32008
rect 23256 31968 23262 31980
rect 17678 31940 17684 31952
rect 17639 31912 17684 31940
rect 17678 31900 17684 31912
rect 17736 31900 17742 31952
rect 23382 31940 23388 31952
rect 23343 31912 23388 31940
rect 23382 31900 23388 31912
rect 23440 31900 23446 31952
rect 23492 31940 23520 31980
rect 23569 31977 23581 32011
rect 23615 32008 23627 32011
rect 24854 32008 24860 32020
rect 23615 31980 24860 32008
rect 23615 31977 23627 31980
rect 23569 31971 23627 31977
rect 24854 31968 24860 31980
rect 24912 31968 24918 32020
rect 28074 31940 28080 31952
rect 23492 31912 28080 31940
rect 28074 31900 28080 31912
rect 28132 31900 28138 31952
rect 17218 31832 17224 31884
rect 17276 31872 17282 31884
rect 23106 31872 23112 31884
rect 17276 31844 17724 31872
rect 17276 31832 17282 31844
rect 5442 31764 5448 31816
rect 5500 31804 5506 31816
rect 14369 31807 14427 31813
rect 14369 31804 14381 31807
rect 5500 31776 14381 31804
rect 5500 31764 5506 31776
rect 14369 31773 14381 31776
rect 14415 31773 14427 31807
rect 14369 31767 14427 31773
rect 17402 31764 17408 31816
rect 17460 31804 17466 31816
rect 17497 31807 17555 31813
rect 17497 31804 17509 31807
rect 17460 31776 17509 31804
rect 17460 31764 17466 31776
rect 17497 31773 17509 31776
rect 17543 31804 17555 31807
rect 17586 31804 17592 31816
rect 17543 31776 17592 31804
rect 17543 31773 17555 31776
rect 17497 31767 17555 31773
rect 17586 31764 17592 31776
rect 17644 31764 17650 31816
rect 17696 31813 17724 31844
rect 22066 31844 23112 31872
rect 17681 31807 17739 31813
rect 17681 31773 17693 31807
rect 17727 31804 17739 31807
rect 22066 31804 22094 31844
rect 23106 31832 23112 31844
rect 23164 31832 23170 31884
rect 27706 31872 27712 31884
rect 27667 31844 27712 31872
rect 27706 31832 27712 31844
rect 27764 31832 27770 31884
rect 33226 31832 33232 31884
rect 33284 31872 33290 31884
rect 34241 31875 34299 31881
rect 33284 31844 33732 31872
rect 33284 31832 33290 31844
rect 17727 31776 22094 31804
rect 17727 31773 17739 31776
rect 17681 31767 17739 31773
rect 27154 31764 27160 31816
rect 27212 31804 27218 31816
rect 27617 31807 27675 31813
rect 27617 31804 27629 31807
rect 27212 31776 27629 31804
rect 27212 31764 27218 31776
rect 27617 31773 27629 31776
rect 27663 31773 27675 31807
rect 27798 31804 27804 31816
rect 27759 31776 27804 31804
rect 27617 31767 27675 31773
rect 27798 31764 27804 31776
rect 27856 31764 27862 31816
rect 33502 31804 33508 31816
rect 33463 31776 33508 31804
rect 33502 31764 33508 31776
rect 33560 31764 33566 31816
rect 33704 31813 33732 31844
rect 34241 31841 34253 31875
rect 34287 31872 34299 31875
rect 34790 31872 34796 31884
rect 34287 31844 34796 31872
rect 34287 31841 34299 31844
rect 34241 31835 34299 31841
rect 34790 31832 34796 31844
rect 34848 31832 34854 31884
rect 35434 31872 35440 31884
rect 35395 31844 35440 31872
rect 35434 31832 35440 31844
rect 35492 31832 35498 31884
rect 33689 31807 33747 31813
rect 33689 31773 33701 31807
rect 33735 31773 33747 31807
rect 33689 31767 33747 31773
rect 33778 31764 33784 31816
rect 33836 31804 33842 31816
rect 34149 31807 34207 31813
rect 34149 31804 34161 31807
rect 33836 31776 34161 31804
rect 33836 31764 33842 31776
rect 34149 31773 34161 31776
rect 34195 31773 34207 31807
rect 34149 31767 34207 31773
rect 34333 31807 34391 31813
rect 34333 31773 34345 31807
rect 34379 31773 34391 31807
rect 34333 31767 34391 31773
rect 14921 31739 14979 31745
rect 14921 31705 14933 31739
rect 14967 31736 14979 31739
rect 15102 31736 15108 31748
rect 14967 31708 15108 31736
rect 14967 31705 14979 31708
rect 14921 31699 14979 31705
rect 15102 31696 15108 31708
rect 15160 31696 15166 31748
rect 34348 31736 34376 31767
rect 34606 31764 34612 31816
rect 34664 31804 34670 31816
rect 35345 31807 35403 31813
rect 35345 31804 35357 31807
rect 34664 31776 35357 31804
rect 34664 31764 34670 31776
rect 35345 31773 35357 31776
rect 35391 31773 35403 31807
rect 35345 31767 35403 31773
rect 34164 31708 34376 31736
rect 34164 31680 34192 31708
rect 33689 31671 33747 31677
rect 33689 31637 33701 31671
rect 33735 31668 33747 31671
rect 34054 31668 34060 31680
rect 33735 31640 34060 31668
rect 33735 31637 33747 31640
rect 33689 31631 33747 31637
rect 34054 31628 34060 31640
rect 34112 31628 34118 31680
rect 34146 31628 34152 31680
rect 34204 31628 34210 31680
rect 34606 31628 34612 31680
rect 34664 31668 34670 31680
rect 34885 31671 34943 31677
rect 34885 31668 34897 31671
rect 34664 31640 34897 31668
rect 34664 31628 34670 31640
rect 34885 31637 34897 31640
rect 34931 31637 34943 31671
rect 34885 31631 34943 31637
rect 35253 31671 35311 31677
rect 35253 31637 35265 31671
rect 35299 31668 35311 31671
rect 35342 31668 35348 31680
rect 35299 31640 35348 31668
rect 35299 31637 35311 31640
rect 35253 31631 35311 31637
rect 35342 31628 35348 31640
rect 35400 31628 35406 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 13814 31464 13820 31476
rect 12912 31436 13820 31464
rect 12912 31405 12940 31436
rect 13814 31424 13820 31436
rect 13872 31424 13878 31476
rect 17221 31467 17279 31473
rect 17221 31433 17233 31467
rect 17267 31464 17279 31467
rect 17862 31464 17868 31476
rect 17267 31436 17868 31464
rect 17267 31433 17279 31436
rect 17221 31427 17279 31433
rect 17862 31424 17868 31436
rect 17920 31424 17926 31476
rect 12897 31399 12955 31405
rect 12897 31365 12909 31399
rect 12943 31365 12955 31399
rect 15289 31399 15347 31405
rect 15289 31396 15301 31399
rect 14122 31368 15301 31396
rect 12897 31359 12955 31365
rect 15289 31365 15301 31368
rect 15335 31365 15347 31399
rect 20714 31396 20720 31408
rect 15289 31359 15347 31365
rect 19720 31368 20720 31396
rect 5261 31331 5319 31337
rect 5261 31297 5273 31331
rect 5307 31328 5319 31331
rect 6730 31328 6736 31340
rect 5307 31300 6736 31328
rect 5307 31297 5319 31300
rect 5261 31291 5319 31297
rect 6730 31288 6736 31300
rect 6788 31288 6794 31340
rect 12618 31328 12624 31340
rect 12579 31300 12624 31328
rect 12618 31288 12624 31300
rect 12676 31288 12682 31340
rect 15013 31331 15071 31337
rect 15013 31297 15025 31331
rect 15059 31297 15071 31331
rect 15013 31291 15071 31297
rect 5534 31260 5540 31272
rect 5495 31232 5540 31260
rect 5534 31220 5540 31232
rect 5592 31220 5598 31272
rect 15028 31260 15056 31291
rect 15102 31288 15108 31340
rect 15160 31328 15166 31340
rect 17126 31328 17132 31340
rect 15160 31300 15205 31328
rect 17087 31300 17132 31328
rect 15160 31288 15166 31300
rect 17126 31288 17132 31300
rect 17184 31288 17190 31340
rect 19720 31337 19748 31368
rect 20714 31356 20720 31368
rect 20772 31356 20778 31408
rect 30561 31399 30619 31405
rect 30561 31365 30573 31399
rect 30607 31396 30619 31399
rect 31018 31396 31024 31408
rect 30607 31368 31024 31396
rect 30607 31365 30619 31368
rect 30561 31359 30619 31365
rect 31018 31356 31024 31368
rect 31076 31356 31082 31408
rect 34514 31396 34520 31408
rect 34475 31368 34520 31396
rect 34514 31356 34520 31368
rect 34572 31356 34578 31408
rect 19705 31331 19763 31337
rect 19705 31297 19717 31331
rect 19751 31297 19763 31331
rect 19705 31291 19763 31297
rect 19797 31331 19855 31337
rect 19797 31297 19809 31331
rect 19843 31297 19855 31331
rect 19978 31328 19984 31340
rect 19939 31300 19984 31328
rect 19797 31291 19855 31297
rect 15838 31260 15844 31272
rect 15028 31232 15844 31260
rect 15838 31220 15844 31232
rect 15896 31220 15902 31272
rect 18874 31220 18880 31272
rect 18932 31260 18938 31272
rect 19153 31263 19211 31269
rect 19153 31260 19165 31263
rect 18932 31232 19165 31260
rect 18932 31220 18938 31232
rect 19153 31229 19165 31232
rect 19199 31229 19211 31263
rect 19153 31223 19211 31229
rect 19242 31220 19248 31272
rect 19300 31260 19306 31272
rect 19812 31260 19840 31291
rect 19978 31288 19984 31300
rect 20036 31288 20042 31340
rect 20530 31328 20536 31340
rect 20491 31300 20536 31328
rect 20530 31288 20536 31300
rect 20588 31288 20594 31340
rect 22278 31288 22284 31340
rect 22336 31328 22342 31340
rect 22373 31331 22431 31337
rect 22373 31328 22385 31331
rect 22336 31300 22385 31328
rect 22336 31288 22342 31300
rect 22373 31297 22385 31300
rect 22419 31297 22431 31331
rect 22373 31291 22431 31297
rect 23385 31331 23443 31337
rect 23385 31297 23397 31331
rect 23431 31328 23443 31331
rect 23566 31328 23572 31340
rect 23431 31300 23572 31328
rect 23431 31297 23443 31300
rect 23385 31291 23443 31297
rect 23566 31288 23572 31300
rect 23624 31288 23630 31340
rect 30377 31331 30435 31337
rect 30377 31297 30389 31331
rect 30423 31328 30435 31331
rect 30466 31328 30472 31340
rect 30423 31300 30472 31328
rect 30423 31297 30435 31300
rect 30377 31291 30435 31297
rect 30466 31288 30472 31300
rect 30524 31288 30530 31340
rect 30650 31288 30656 31340
rect 30708 31328 30714 31340
rect 34054 31328 34060 31340
rect 30708 31300 30753 31328
rect 34015 31300 34060 31328
rect 30708 31288 30714 31300
rect 34054 31288 34060 31300
rect 34112 31288 34118 31340
rect 34146 31288 34152 31340
rect 34204 31328 34210 31340
rect 34204 31300 34249 31328
rect 34204 31288 34210 31300
rect 20254 31260 20260 31272
rect 19300 31232 19840 31260
rect 20215 31232 20260 31260
rect 19300 31220 19306 31232
rect 20254 31220 20260 31232
rect 20312 31220 20318 31272
rect 33778 31260 33784 31272
rect 33739 31232 33784 31260
rect 33778 31220 33784 31232
rect 33836 31220 33842 31272
rect 5353 31195 5411 31201
rect 5353 31161 5365 31195
rect 5399 31192 5411 31195
rect 6822 31192 6828 31204
rect 5399 31164 6828 31192
rect 5399 31161 5411 31164
rect 5353 31155 5411 31161
rect 6822 31152 6828 31164
rect 6880 31152 6886 31204
rect 23198 31192 23204 31204
rect 23159 31164 23204 31192
rect 23198 31152 23204 31164
rect 23256 31152 23262 31204
rect 34422 31152 34428 31204
rect 34480 31192 34486 31204
rect 34701 31195 34759 31201
rect 34701 31192 34713 31195
rect 34480 31164 34713 31192
rect 34480 31152 34486 31164
rect 34701 31161 34713 31164
rect 34747 31161 34759 31195
rect 34701 31155 34759 31161
rect 5442 31084 5448 31136
rect 5500 31124 5506 31136
rect 5500 31096 5545 31124
rect 5500 31084 5506 31096
rect 12066 31084 12072 31136
rect 12124 31124 12130 31136
rect 14369 31127 14427 31133
rect 14369 31124 14381 31127
rect 12124 31096 14381 31124
rect 12124 31084 12130 31096
rect 14369 31093 14381 31096
rect 14415 31093 14427 31127
rect 22370 31124 22376 31136
rect 22331 31096 22376 31124
rect 14369 31087 14427 31093
rect 22370 31084 22376 31096
rect 22428 31084 22434 31136
rect 29822 31084 29828 31136
rect 29880 31124 29886 31136
rect 30193 31127 30251 31133
rect 30193 31124 30205 31127
rect 29880 31096 30205 31124
rect 29880 31084 29886 31096
rect 30193 31093 30205 31096
rect 30239 31093 30251 31127
rect 30193 31087 30251 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 29638 30880 29644 30932
rect 29696 30920 29702 30932
rect 33873 30923 33931 30929
rect 29696 30892 30144 30920
rect 29696 30880 29702 30892
rect 14366 30852 14372 30864
rect 14327 30824 14372 30852
rect 14366 30812 14372 30824
rect 14424 30812 14430 30864
rect 18230 30812 18236 30864
rect 18288 30852 18294 30864
rect 19978 30852 19984 30864
rect 18288 30824 19984 30852
rect 18288 30812 18294 30824
rect 19978 30812 19984 30824
rect 20036 30852 20042 30864
rect 21085 30855 21143 30861
rect 20036 30824 20116 30852
rect 20036 30812 20042 30824
rect 4341 30787 4399 30793
rect 4341 30753 4353 30787
rect 4387 30784 4399 30787
rect 5258 30784 5264 30796
rect 4387 30756 5264 30784
rect 4387 30753 4399 30756
rect 4341 30747 4399 30753
rect 5258 30744 5264 30756
rect 5316 30744 5322 30796
rect 10318 30744 10324 30796
rect 10376 30784 10382 30796
rect 11057 30787 11115 30793
rect 11057 30784 11069 30787
rect 10376 30756 11069 30784
rect 10376 30744 10382 30756
rect 11057 30753 11069 30756
rect 11103 30753 11115 30787
rect 19242 30784 19248 30796
rect 11057 30747 11115 30753
rect 18432 30756 19248 30784
rect 18432 30728 18460 30756
rect 19242 30744 19248 30756
rect 19300 30784 19306 30796
rect 19300 30756 20024 30784
rect 19300 30744 19306 30756
rect 4614 30716 4620 30728
rect 4575 30688 4620 30716
rect 4614 30676 4620 30688
rect 4672 30676 4678 30728
rect 8478 30676 8484 30728
rect 8536 30716 8542 30728
rect 9861 30719 9919 30725
rect 9861 30716 9873 30719
rect 8536 30688 9873 30716
rect 8536 30676 8542 30688
rect 9861 30685 9873 30688
rect 9907 30685 9919 30719
rect 9861 30679 9919 30685
rect 10873 30719 10931 30725
rect 10873 30685 10885 30719
rect 10919 30716 10931 30719
rect 12066 30716 12072 30728
rect 10919 30688 12072 30716
rect 10919 30685 10931 30688
rect 10873 30679 10931 30685
rect 12066 30676 12072 30688
rect 12124 30676 12130 30728
rect 14369 30719 14427 30725
rect 14369 30685 14381 30719
rect 14415 30685 14427 30719
rect 14550 30716 14556 30728
rect 14511 30688 14556 30716
rect 14369 30679 14427 30685
rect 5994 30648 6000 30660
rect 5955 30620 6000 30648
rect 5994 30608 6000 30620
rect 6052 30608 6058 30660
rect 9677 30651 9735 30657
rect 9677 30617 9689 30651
rect 9723 30648 9735 30651
rect 9766 30648 9772 30660
rect 9723 30620 9772 30648
rect 9723 30617 9735 30620
rect 9677 30611 9735 30617
rect 9766 30608 9772 30620
rect 9824 30608 9830 30660
rect 14384 30648 14412 30679
rect 14550 30676 14556 30688
rect 14608 30716 14614 30728
rect 15102 30716 15108 30728
rect 14608 30688 15108 30716
rect 14608 30676 14614 30688
rect 15102 30676 15108 30688
rect 15160 30676 15166 30728
rect 18138 30716 18144 30728
rect 18099 30688 18144 30716
rect 18138 30676 18144 30688
rect 18196 30676 18202 30728
rect 18414 30716 18420 30728
rect 18375 30688 18420 30716
rect 18414 30676 18420 30688
rect 18472 30676 18478 30728
rect 19996 30725 20024 30756
rect 19889 30719 19947 30725
rect 19889 30685 19901 30719
rect 19935 30685 19947 30719
rect 19889 30679 19947 30685
rect 19981 30719 20039 30725
rect 19981 30685 19993 30719
rect 20027 30685 20039 30719
rect 20088 30716 20116 30824
rect 21085 30821 21097 30855
rect 21131 30852 21143 30855
rect 21174 30852 21180 30864
rect 21131 30824 21180 30852
rect 21131 30821 21143 30824
rect 21085 30815 21143 30821
rect 21174 30812 21180 30824
rect 21232 30812 21238 30864
rect 29089 30855 29147 30861
rect 29089 30821 29101 30855
rect 29135 30852 29147 30855
rect 29914 30852 29920 30864
rect 29135 30824 29920 30852
rect 29135 30821 29147 30824
rect 29089 30815 29147 30821
rect 29914 30812 29920 30824
rect 29972 30812 29978 30864
rect 20806 30744 20812 30796
rect 20864 30784 20870 30796
rect 20864 30756 21220 30784
rect 20864 30744 20870 30756
rect 20349 30719 20407 30725
rect 20349 30716 20361 30719
rect 20088 30688 20361 30716
rect 19981 30679 20039 30685
rect 20349 30685 20361 30688
rect 20395 30685 20407 30719
rect 20898 30716 20904 30728
rect 20859 30688 20904 30716
rect 20349 30679 20407 30685
rect 15838 30648 15844 30660
rect 14384 30620 15844 30648
rect 15838 30608 15844 30620
rect 15896 30608 15902 30660
rect 19904 30648 19932 30679
rect 20898 30676 20904 30688
rect 20956 30676 20962 30728
rect 21192 30725 21220 30756
rect 29730 30744 29736 30796
rect 29788 30784 29794 30796
rect 30116 30793 30144 30892
rect 33873 30889 33885 30923
rect 33919 30920 33931 30923
rect 34146 30920 34152 30932
rect 33919 30892 34152 30920
rect 33919 30889 33931 30892
rect 33873 30883 33931 30889
rect 34146 30880 34152 30892
rect 34204 30880 34210 30932
rect 35434 30852 35440 30864
rect 31128 30824 35112 30852
rect 35395 30824 35440 30852
rect 30009 30787 30067 30793
rect 30009 30784 30021 30787
rect 29788 30756 30021 30784
rect 29788 30744 29794 30756
rect 30009 30753 30021 30756
rect 30055 30753 30067 30787
rect 30009 30747 30067 30753
rect 30101 30787 30159 30793
rect 30101 30753 30113 30787
rect 30147 30753 30159 30787
rect 30101 30747 30159 30753
rect 30466 30744 30472 30796
rect 30524 30784 30530 30796
rect 31128 30793 31156 30824
rect 31113 30787 31171 30793
rect 31113 30784 31125 30787
rect 30524 30756 31125 30784
rect 30524 30744 30530 30756
rect 31113 30753 31125 30756
rect 31159 30753 31171 30787
rect 31113 30747 31171 30753
rect 31205 30787 31263 30793
rect 31205 30753 31217 30787
rect 31251 30784 31263 30787
rect 34606 30784 34612 30796
rect 31251 30756 34612 30784
rect 31251 30753 31263 30756
rect 31205 30747 31263 30753
rect 21177 30719 21235 30725
rect 21177 30685 21189 30719
rect 21223 30685 21235 30719
rect 21177 30679 21235 30685
rect 29917 30719 29975 30725
rect 29917 30685 29929 30719
rect 29963 30685 29975 30719
rect 29917 30679 29975 30685
rect 20714 30648 20720 30660
rect 19904 30620 20720 30648
rect 20714 30608 20720 30620
rect 20772 30608 20778 30660
rect 28074 30608 28080 30660
rect 28132 30648 28138 30660
rect 28721 30651 28779 30657
rect 28721 30648 28733 30651
rect 28132 30620 28733 30648
rect 28132 30608 28138 30620
rect 28721 30617 28733 30620
rect 28767 30617 28779 30651
rect 29932 30648 29960 30679
rect 30190 30676 30196 30728
rect 30248 30716 30254 30728
rect 30248 30688 30293 30716
rect 30248 30676 30254 30688
rect 30558 30676 30564 30728
rect 30616 30716 30622 30728
rect 30929 30719 30987 30725
rect 30929 30716 30941 30719
rect 30616 30688 30941 30716
rect 30616 30676 30622 30688
rect 30929 30685 30941 30688
rect 30975 30685 30987 30719
rect 30929 30679 30987 30685
rect 31018 30676 31024 30728
rect 31076 30716 31082 30728
rect 31076 30688 31121 30716
rect 31076 30676 31082 30688
rect 31220 30648 31248 30747
rect 34606 30744 34612 30756
rect 34664 30744 34670 30796
rect 34790 30744 34796 30796
rect 34848 30784 34854 30796
rect 34977 30787 35035 30793
rect 34977 30784 34989 30787
rect 34848 30756 34989 30784
rect 34848 30744 34854 30756
rect 34977 30753 34989 30756
rect 35023 30753 35035 30787
rect 34977 30747 35035 30753
rect 33781 30719 33839 30725
rect 33781 30685 33793 30719
rect 33827 30716 33839 30719
rect 33870 30716 33876 30728
rect 33827 30688 33876 30716
rect 33827 30685 33839 30688
rect 33781 30679 33839 30685
rect 33870 30676 33876 30688
rect 33928 30676 33934 30728
rect 35084 30725 35112 30824
rect 35434 30812 35440 30824
rect 35492 30812 35498 30864
rect 33965 30719 34023 30725
rect 33965 30685 33977 30719
rect 34011 30685 34023 30719
rect 33965 30679 34023 30685
rect 35069 30719 35127 30725
rect 35069 30685 35081 30719
rect 35115 30685 35127 30719
rect 35069 30679 35127 30685
rect 29932 30620 31248 30648
rect 28721 30611 28779 30617
rect 33410 30608 33416 30660
rect 33468 30648 33474 30660
rect 33686 30648 33692 30660
rect 33468 30620 33692 30648
rect 33468 30608 33474 30620
rect 33686 30608 33692 30620
rect 33744 30648 33750 30660
rect 33980 30648 34008 30679
rect 33744 30620 34008 30648
rect 33744 30608 33750 30620
rect 9398 30540 9404 30592
rect 9456 30580 9462 30592
rect 10045 30583 10103 30589
rect 10045 30580 10057 30583
rect 9456 30552 10057 30580
rect 9456 30540 9462 30552
rect 10045 30549 10057 30552
rect 10091 30549 10103 30583
rect 17954 30580 17960 30592
rect 17915 30552 17960 30580
rect 10045 30543 10103 30549
rect 17954 30540 17960 30552
rect 18012 30540 18018 30592
rect 18322 30580 18328 30592
rect 18283 30552 18328 30580
rect 18322 30540 18328 30552
rect 18380 30540 18386 30592
rect 29178 30580 29184 30592
rect 29139 30552 29184 30580
rect 29178 30540 29184 30552
rect 29236 30540 29242 30592
rect 29270 30540 29276 30592
rect 29328 30580 29334 30592
rect 29733 30583 29791 30589
rect 29733 30580 29745 30583
rect 29328 30552 29745 30580
rect 29328 30540 29334 30552
rect 29733 30549 29745 30552
rect 29779 30549 29791 30583
rect 29733 30543 29791 30549
rect 29914 30540 29920 30592
rect 29972 30580 29978 30592
rect 30745 30583 30803 30589
rect 30745 30580 30757 30583
rect 29972 30552 30757 30580
rect 29972 30540 29978 30552
rect 30745 30549 30757 30552
rect 30791 30549 30803 30583
rect 30745 30543 30803 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 4614 30336 4620 30388
rect 4672 30376 4678 30388
rect 4801 30379 4859 30385
rect 4801 30376 4813 30379
rect 4672 30348 4813 30376
rect 4672 30336 4678 30348
rect 4801 30345 4813 30348
rect 4847 30345 4859 30379
rect 4801 30339 4859 30345
rect 18782 30336 18788 30388
rect 18840 30376 18846 30388
rect 18877 30379 18935 30385
rect 18877 30376 18889 30379
rect 18840 30348 18889 30376
rect 18840 30336 18846 30348
rect 18877 30345 18889 30348
rect 18923 30345 18935 30379
rect 18877 30339 18935 30345
rect 19058 30336 19064 30388
rect 19116 30376 19122 30388
rect 19116 30348 20576 30376
rect 19116 30336 19122 30348
rect 5442 30308 5448 30320
rect 5403 30280 5448 30308
rect 5442 30268 5448 30280
rect 5500 30268 5506 30320
rect 6730 30308 6736 30320
rect 6691 30280 6736 30308
rect 6730 30268 6736 30280
rect 6788 30308 6794 30320
rect 7098 30308 7104 30320
rect 6788 30280 7104 30308
rect 6788 30268 6794 30280
rect 7098 30268 7104 30280
rect 7156 30268 7162 30320
rect 8772 30280 9628 30308
rect 5077 30243 5135 30249
rect 5077 30209 5089 30243
rect 5123 30240 5135 30243
rect 6362 30240 6368 30252
rect 5123 30212 6368 30240
rect 5123 30209 5135 30212
rect 5077 30203 5135 30209
rect 6362 30200 6368 30212
rect 6420 30200 6426 30252
rect 6454 30200 6460 30252
rect 6512 30240 6518 30252
rect 6549 30243 6607 30249
rect 6549 30240 6561 30243
rect 6512 30212 6561 30240
rect 6512 30200 6518 30212
rect 6549 30209 6561 30212
rect 6595 30209 6607 30243
rect 6549 30203 6607 30209
rect 6822 30200 6828 30252
rect 6880 30240 6886 30252
rect 6880 30212 6925 30240
rect 6880 30200 6886 30212
rect 8386 30200 8392 30252
rect 8444 30240 8450 30252
rect 8772 30249 8800 30280
rect 8757 30243 8815 30249
rect 8757 30240 8769 30243
rect 8444 30212 8769 30240
rect 8444 30200 8450 30212
rect 8757 30209 8769 30212
rect 8803 30209 8815 30243
rect 8757 30203 8815 30209
rect 8941 30243 8999 30249
rect 8941 30209 8953 30243
rect 8987 30209 8999 30243
rect 9600 30226 9628 30280
rect 9766 30268 9772 30320
rect 9824 30308 9830 30320
rect 10229 30311 10287 30317
rect 10229 30308 10241 30311
rect 9824 30280 10241 30308
rect 9824 30268 9830 30280
rect 10229 30277 10241 30280
rect 10275 30277 10287 30311
rect 14366 30308 14372 30320
rect 14306 30280 14372 30308
rect 10229 30271 10287 30277
rect 14366 30268 14372 30280
rect 14424 30268 14430 30320
rect 17221 30311 17279 30317
rect 17221 30277 17233 30311
rect 17267 30308 17279 30311
rect 18138 30308 18144 30320
rect 17267 30280 18144 30308
rect 17267 30277 17279 30280
rect 17221 30271 17279 30277
rect 18138 30268 18144 30280
rect 18196 30268 18202 30320
rect 20548 30308 20576 30348
rect 20714 30336 20720 30388
rect 20772 30376 20778 30388
rect 20834 30379 20892 30385
rect 20834 30376 20846 30379
rect 20772 30348 20846 30376
rect 20772 30336 20778 30348
rect 20834 30345 20846 30348
rect 20880 30345 20892 30379
rect 33870 30376 33876 30388
rect 20834 30339 20892 30345
rect 33612 30348 33876 30376
rect 22278 30308 22284 30320
rect 20548 30280 22284 30308
rect 10962 30240 10968 30252
rect 10923 30212 10968 30240
rect 8941 30203 8999 30209
rect 4985 30175 5043 30181
rect 4985 30141 4997 30175
rect 5031 30141 5043 30175
rect 4985 30135 5043 30141
rect 5353 30175 5411 30181
rect 5353 30141 5365 30175
rect 5399 30141 5411 30175
rect 5353 30135 5411 30141
rect 5000 30036 5028 30135
rect 5368 30104 5396 30135
rect 5994 30132 6000 30184
rect 6052 30172 6058 30184
rect 6638 30172 6644 30184
rect 6052 30144 6644 30172
rect 6052 30132 6058 30144
rect 6638 30132 6644 30144
rect 6696 30172 6702 30184
rect 8846 30172 8852 30184
rect 6696 30144 8852 30172
rect 6696 30132 6702 30144
rect 8846 30132 8852 30144
rect 8904 30132 8910 30184
rect 6549 30107 6607 30113
rect 6549 30104 6561 30107
rect 5368 30076 6561 30104
rect 6549 30073 6561 30076
rect 6595 30073 6607 30107
rect 8956 30104 8984 30203
rect 10962 30200 10968 30212
rect 11020 30200 11026 30252
rect 15105 30243 15163 30249
rect 15105 30209 15117 30243
rect 15151 30209 15163 30243
rect 15105 30203 15163 30209
rect 9677 30175 9735 30181
rect 9677 30141 9689 30175
rect 9723 30141 9735 30175
rect 9677 30135 9735 30141
rect 9692 30104 9720 30135
rect 10778 30132 10784 30184
rect 10836 30172 10842 30184
rect 10836 30144 12434 30172
rect 10836 30132 10842 30144
rect 11146 30104 11152 30116
rect 8956 30076 11152 30104
rect 6549 30067 6607 30073
rect 11146 30064 11152 30076
rect 11204 30064 11210 30116
rect 5718 30036 5724 30048
rect 5000 30008 5724 30036
rect 5718 29996 5724 30008
rect 5776 29996 5782 30048
rect 6914 29996 6920 30048
rect 6972 30036 6978 30048
rect 8849 30039 8907 30045
rect 8849 30036 8861 30039
rect 6972 30008 8861 30036
rect 6972 29996 6978 30008
rect 8849 30005 8861 30008
rect 8895 30005 8907 30039
rect 11054 30036 11060 30048
rect 11015 30008 11060 30036
rect 8849 29999 8907 30005
rect 11054 29996 11060 30008
rect 11112 29996 11118 30048
rect 12406 30036 12434 30144
rect 12710 30132 12716 30184
rect 12768 30172 12774 30184
rect 12805 30175 12863 30181
rect 12805 30172 12817 30175
rect 12768 30144 12817 30172
rect 12768 30132 12774 30144
rect 12805 30141 12817 30144
rect 12851 30141 12863 30175
rect 12805 30135 12863 30141
rect 13081 30175 13139 30181
rect 13081 30141 13093 30175
rect 13127 30172 13139 30175
rect 14090 30172 14096 30184
rect 13127 30144 14096 30172
rect 13127 30141 13139 30144
rect 13081 30135 13139 30141
rect 14090 30132 14096 30144
rect 14148 30172 14154 30184
rect 15120 30172 15148 30203
rect 15194 30200 15200 30252
rect 15252 30240 15258 30252
rect 15289 30243 15347 30249
rect 15289 30240 15301 30243
rect 15252 30212 15301 30240
rect 15252 30200 15258 30212
rect 15289 30209 15301 30212
rect 15335 30209 15347 30243
rect 15289 30203 15347 30209
rect 16666 30200 16672 30252
rect 16724 30240 16730 30252
rect 17126 30240 17132 30252
rect 16724 30212 17132 30240
rect 16724 30200 16730 30212
rect 17126 30200 17132 30212
rect 17184 30200 17190 30252
rect 17313 30243 17371 30249
rect 17313 30209 17325 30243
rect 17359 30240 17371 30243
rect 17402 30240 17408 30252
rect 17359 30212 17408 30240
rect 17359 30209 17371 30212
rect 17313 30203 17371 30209
rect 17402 30200 17408 30212
rect 17460 30200 17466 30252
rect 17954 30200 17960 30252
rect 18012 30240 18018 30252
rect 20548 30249 20576 30280
rect 22278 30268 22284 30280
rect 22336 30268 22342 30320
rect 28353 30311 28411 30317
rect 28353 30277 28365 30311
rect 28399 30308 28411 30311
rect 29178 30308 29184 30320
rect 28399 30280 29184 30308
rect 28399 30277 28411 30280
rect 28353 30271 28411 30277
rect 29178 30268 29184 30280
rect 29236 30268 29242 30320
rect 29914 30308 29920 30320
rect 29472 30280 29920 30308
rect 20533 30243 20591 30249
rect 18012 30212 18630 30240
rect 18012 30200 18018 30212
rect 20533 30209 20545 30243
rect 20579 30209 20591 30243
rect 20714 30240 20720 30252
rect 20675 30212 20720 30240
rect 20533 30203 20591 30209
rect 20714 30200 20720 30212
rect 20772 30200 20778 30252
rect 21266 30240 21272 30252
rect 21227 30212 21272 30240
rect 21266 30200 21272 30212
rect 21324 30200 21330 30252
rect 24302 30240 24308 30252
rect 24263 30212 24308 30240
rect 24302 30200 24308 30212
rect 24360 30200 24366 30252
rect 24489 30243 24547 30249
rect 24489 30209 24501 30243
rect 24535 30240 24547 30243
rect 24946 30240 24952 30252
rect 24535 30212 24952 30240
rect 24535 30209 24547 30212
rect 24489 30203 24547 30209
rect 24946 30200 24952 30212
rect 25004 30200 25010 30252
rect 28166 30240 28172 30252
rect 28127 30212 28172 30240
rect 28166 30200 28172 30212
rect 28224 30200 28230 30252
rect 28445 30243 28503 30249
rect 28445 30209 28457 30243
rect 28491 30240 28503 30243
rect 29270 30240 29276 30252
rect 28491 30212 29276 30240
rect 28491 30209 28503 30212
rect 28445 30203 28503 30209
rect 29270 30200 29276 30212
rect 29328 30200 29334 30252
rect 29472 30249 29500 30280
rect 29914 30268 29920 30280
rect 29972 30268 29978 30320
rect 31018 30308 31024 30320
rect 30760 30280 31024 30308
rect 29457 30243 29515 30249
rect 29457 30209 29469 30243
rect 29503 30209 29515 30243
rect 29641 30243 29699 30249
rect 29641 30240 29653 30243
rect 29457 30203 29515 30209
rect 29564 30212 29653 30240
rect 14148 30144 15148 30172
rect 17865 30175 17923 30181
rect 14148 30132 14154 30144
rect 17865 30141 17877 30175
rect 17911 30172 17923 30175
rect 18690 30172 18696 30184
rect 17911 30144 18696 30172
rect 17911 30141 17923 30144
rect 17865 30135 17923 30141
rect 18690 30132 18696 30144
rect 18748 30132 18754 30184
rect 18874 30132 18880 30184
rect 18932 30132 18938 30184
rect 20254 30132 20260 30184
rect 20312 30172 20318 30184
rect 20312 30144 20838 30172
rect 20312 30132 20318 30144
rect 22370 30132 22376 30184
rect 22428 30172 22434 30184
rect 25314 30172 25320 30184
rect 22428 30144 25320 30172
rect 22428 30132 22434 30144
rect 25314 30132 25320 30144
rect 25372 30172 25378 30184
rect 25958 30172 25964 30184
rect 25372 30144 25964 30172
rect 25372 30132 25378 30144
rect 25958 30132 25964 30144
rect 26016 30132 26022 30184
rect 28074 30132 28080 30184
rect 28132 30172 28138 30184
rect 29564 30172 29592 30212
rect 29641 30209 29653 30212
rect 29687 30209 29699 30243
rect 29822 30240 29828 30252
rect 29783 30212 29828 30240
rect 29641 30203 29699 30209
rect 29822 30200 29828 30212
rect 29880 30200 29886 30252
rect 30558 30240 30564 30252
rect 30519 30212 30564 30240
rect 30558 30200 30564 30212
rect 30616 30200 30622 30252
rect 30760 30249 30788 30280
rect 31018 30268 31024 30280
rect 31076 30308 31082 30320
rect 32401 30311 32459 30317
rect 32401 30308 32413 30311
rect 31076 30280 32413 30308
rect 31076 30268 31082 30280
rect 32401 30277 32413 30280
rect 32447 30277 32459 30311
rect 32401 30271 32459 30277
rect 30745 30243 30803 30249
rect 30745 30209 30757 30243
rect 30791 30209 30803 30243
rect 30745 30203 30803 30209
rect 32214 30200 32220 30252
rect 32272 30240 32278 30252
rect 32309 30243 32367 30249
rect 32309 30240 32321 30243
rect 32272 30212 32321 30240
rect 32272 30200 32278 30212
rect 32309 30209 32321 30212
rect 32355 30209 32367 30243
rect 32309 30203 32367 30209
rect 32677 30243 32735 30249
rect 32677 30209 32689 30243
rect 32723 30209 32735 30243
rect 32950 30240 32956 30252
rect 32911 30212 32956 30240
rect 32677 30203 32735 30209
rect 28132 30144 29592 30172
rect 28132 30132 28138 30144
rect 32398 30132 32404 30184
rect 32456 30172 32462 30184
rect 32692 30172 32720 30203
rect 32950 30200 32956 30212
rect 33008 30200 33014 30252
rect 33134 30200 33140 30252
rect 33192 30240 33198 30252
rect 33612 30249 33640 30348
rect 33870 30336 33876 30348
rect 33928 30336 33934 30388
rect 33686 30268 33692 30320
rect 33744 30308 33750 30320
rect 33781 30311 33839 30317
rect 33781 30308 33793 30311
rect 33744 30280 33793 30308
rect 33744 30268 33750 30280
rect 33781 30277 33793 30280
rect 33827 30277 33839 30311
rect 33781 30271 33839 30277
rect 33597 30243 33655 30249
rect 33597 30240 33609 30243
rect 33192 30212 33609 30240
rect 33192 30200 33198 30212
rect 33597 30209 33609 30212
rect 33643 30209 33655 30243
rect 33597 30203 33655 30209
rect 33873 30243 33931 30249
rect 33873 30209 33885 30243
rect 33919 30240 33931 30243
rect 34422 30240 34428 30252
rect 33919 30212 34428 30240
rect 33919 30209 33931 30212
rect 33873 30203 33931 30209
rect 33413 30175 33471 30181
rect 33413 30172 33425 30175
rect 32456 30144 33425 30172
rect 32456 30132 32462 30144
rect 33413 30141 33425 30144
rect 33459 30141 33471 30175
rect 33413 30135 33471 30141
rect 18598 30064 18604 30116
rect 18656 30104 18662 30116
rect 18656 30076 28304 30104
rect 18656 30064 18662 30076
rect 14553 30039 14611 30045
rect 14553 30036 14565 30039
rect 12406 30008 14565 30036
rect 14553 30005 14565 30008
rect 14599 30005 14611 30039
rect 14553 29999 14611 30005
rect 14826 29996 14832 30048
rect 14884 30036 14890 30048
rect 15197 30039 15255 30045
rect 15197 30036 15209 30039
rect 14884 30008 15209 30036
rect 14884 29996 14890 30008
rect 15197 30005 15209 30008
rect 15243 30005 15255 30039
rect 15197 29999 15255 30005
rect 23934 29996 23940 30048
rect 23992 30036 23998 30048
rect 24305 30039 24363 30045
rect 24305 30036 24317 30039
rect 23992 30008 24317 30036
rect 23992 29996 23998 30008
rect 24305 30005 24317 30008
rect 24351 30005 24363 30039
rect 24305 29999 24363 30005
rect 27982 29996 27988 30048
rect 28040 30036 28046 30048
rect 28169 30039 28227 30045
rect 28169 30036 28181 30039
rect 28040 30008 28181 30036
rect 28040 29996 28046 30008
rect 28169 30005 28181 30008
rect 28215 30005 28227 30039
rect 28276 30036 28304 30076
rect 28350 30064 28356 30116
rect 28408 30104 28414 30116
rect 29273 30107 29331 30113
rect 29273 30104 29285 30107
rect 28408 30076 29285 30104
rect 28408 30064 28414 30076
rect 29273 30073 29285 30076
rect 29319 30073 29331 30107
rect 29273 30067 29331 30073
rect 29380 30076 30880 30104
rect 29380 30036 29408 30076
rect 28276 30008 29408 30036
rect 28169 29999 28227 30005
rect 29730 29996 29736 30048
rect 29788 30036 29794 30048
rect 30653 30039 30711 30045
rect 30653 30036 30665 30039
rect 29788 30008 30665 30036
rect 29788 29996 29794 30008
rect 30653 30005 30665 30008
rect 30699 30005 30711 30039
rect 30852 30036 30880 30076
rect 33318 30064 33324 30116
rect 33376 30104 33382 30116
rect 33888 30104 33916 30203
rect 34422 30200 34428 30212
rect 34480 30200 34486 30252
rect 33376 30076 33916 30104
rect 33376 30064 33382 30076
rect 34238 30036 34244 30048
rect 30852 30008 34244 30036
rect 30653 29999 30711 30005
rect 34238 29996 34244 30008
rect 34296 29996 34302 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 6454 29832 6460 29844
rect 6415 29804 6460 29832
rect 6454 29792 6460 29804
rect 6512 29792 6518 29844
rect 6638 29792 6644 29844
rect 6696 29792 6702 29844
rect 6730 29792 6736 29844
rect 6788 29792 6794 29844
rect 6822 29792 6828 29844
rect 6880 29832 6886 29844
rect 7561 29835 7619 29841
rect 7561 29832 7573 29835
rect 6880 29804 7573 29832
rect 6880 29792 6886 29804
rect 7561 29801 7573 29804
rect 7607 29801 7619 29835
rect 10778 29832 10784 29844
rect 7561 29795 7619 29801
rect 8128 29804 10784 29832
rect 5169 29699 5227 29705
rect 5169 29665 5181 29699
rect 5215 29696 5227 29699
rect 5350 29696 5356 29708
rect 5215 29668 5356 29696
rect 5215 29665 5227 29668
rect 5169 29659 5227 29665
rect 5350 29656 5356 29668
rect 5408 29656 5414 29708
rect 6656 29696 6684 29792
rect 6748 29764 6776 29792
rect 6748 29736 6960 29764
rect 6932 29705 6960 29736
rect 7098 29724 7104 29776
rect 7156 29764 7162 29776
rect 8018 29764 8024 29776
rect 7156 29736 8024 29764
rect 7156 29724 7162 29736
rect 8018 29724 8024 29736
rect 8076 29724 8082 29776
rect 6733 29699 6791 29705
rect 6733 29696 6745 29699
rect 6656 29668 6745 29696
rect 6733 29665 6745 29668
rect 6779 29665 6791 29699
rect 6733 29659 6791 29665
rect 6917 29699 6975 29705
rect 6917 29665 6929 29699
rect 6963 29665 6975 29699
rect 8128 29696 8156 29804
rect 10778 29792 10784 29804
rect 10836 29792 10842 29844
rect 18414 29792 18420 29844
rect 18472 29832 18478 29844
rect 18509 29835 18567 29841
rect 18509 29832 18521 29835
rect 18472 29804 18521 29832
rect 18472 29792 18478 29804
rect 18509 29801 18521 29804
rect 18555 29801 18567 29835
rect 24765 29835 24823 29841
rect 18509 29795 18567 29801
rect 19352 29804 20852 29832
rect 8294 29764 8300 29776
rect 8255 29736 8300 29764
rect 8294 29724 8300 29736
rect 8352 29724 8358 29776
rect 9125 29767 9183 29773
rect 9125 29733 9137 29767
rect 9171 29764 9183 29767
rect 9674 29764 9680 29776
rect 9171 29736 9680 29764
rect 9171 29733 9183 29736
rect 9125 29727 9183 29733
rect 9674 29724 9680 29736
rect 9732 29724 9738 29776
rect 10962 29764 10968 29776
rect 9968 29736 10968 29764
rect 9766 29696 9772 29708
rect 6917 29659 6975 29665
rect 7392 29668 8156 29696
rect 8312 29668 9772 29696
rect 4157 29631 4215 29637
rect 4157 29597 4169 29631
rect 4203 29597 4215 29631
rect 4157 29591 4215 29597
rect 4341 29631 4399 29637
rect 4341 29597 4353 29631
rect 4387 29628 4399 29631
rect 4982 29628 4988 29640
rect 4387 29600 4988 29628
rect 4387 29597 4399 29600
rect 4341 29591 4399 29597
rect 4172 29492 4200 29591
rect 4982 29588 4988 29600
rect 5040 29588 5046 29640
rect 5534 29588 5540 29640
rect 5592 29588 5598 29640
rect 6641 29631 6699 29637
rect 6641 29597 6653 29631
rect 6687 29597 6699 29631
rect 6641 29591 6699 29597
rect 6825 29631 6883 29637
rect 6825 29597 6837 29631
rect 6871 29628 6883 29631
rect 7392 29628 7420 29668
rect 8312 29637 8340 29668
rect 9766 29656 9772 29668
rect 9824 29656 9830 29708
rect 6871 29600 7420 29628
rect 7469 29631 7527 29637
rect 6871 29597 6883 29600
rect 6825 29591 6883 29597
rect 7469 29597 7481 29631
rect 7515 29597 7527 29631
rect 7469 29591 7527 29597
rect 8297 29631 8355 29637
rect 8297 29597 8309 29631
rect 8343 29597 8355 29631
rect 8478 29628 8484 29640
rect 8439 29600 8484 29628
rect 8297 29591 8355 29597
rect 4433 29563 4491 29569
rect 4433 29529 4445 29563
rect 4479 29560 4491 29563
rect 5552 29560 5580 29588
rect 4479 29532 5580 29560
rect 5997 29563 6055 29569
rect 4479 29529 4491 29532
rect 4433 29523 4491 29529
rect 5997 29529 6009 29563
rect 6043 29560 6055 29563
rect 6086 29560 6092 29572
rect 6043 29532 6092 29560
rect 6043 29529 6055 29532
rect 5997 29523 6055 29529
rect 6086 29520 6092 29532
rect 6144 29520 6150 29572
rect 6656 29560 6684 29591
rect 7484 29560 7512 29591
rect 8478 29588 8484 29600
rect 8536 29588 8542 29640
rect 9306 29628 9312 29640
rect 8680 29600 9312 29628
rect 6656 29532 7512 29560
rect 5166 29492 5172 29504
rect 4172 29464 5172 29492
rect 5166 29452 5172 29464
rect 5224 29452 5230 29504
rect 5442 29452 5448 29504
rect 5500 29492 5506 29504
rect 6656 29492 6684 29532
rect 5500 29464 6684 29492
rect 7484 29492 7512 29532
rect 8018 29520 8024 29572
rect 8076 29560 8082 29572
rect 8680 29560 8708 29600
rect 9306 29588 9312 29600
rect 9364 29588 9370 29640
rect 9401 29631 9459 29637
rect 9401 29597 9413 29631
rect 9447 29628 9459 29631
rect 9968 29628 9996 29736
rect 10962 29724 10968 29736
rect 11020 29724 11026 29776
rect 11146 29764 11152 29776
rect 11107 29736 11152 29764
rect 11146 29724 11152 29736
rect 11204 29724 11210 29776
rect 19352 29764 19380 29804
rect 19978 29764 19984 29776
rect 16546 29736 19380 29764
rect 19536 29736 19984 29764
rect 13814 29696 13820 29708
rect 13556 29668 13820 29696
rect 10318 29628 10324 29640
rect 9447 29600 9996 29628
rect 10279 29600 10324 29628
rect 9447 29597 9459 29600
rect 9401 29591 9459 29597
rect 10318 29588 10324 29600
rect 10376 29588 10382 29640
rect 10962 29588 10968 29640
rect 11020 29628 11026 29640
rect 13556 29637 13584 29668
rect 13814 29656 13820 29668
rect 13872 29656 13878 29708
rect 16546 29696 16574 29736
rect 18138 29696 18144 29708
rect 15120 29668 16574 29696
rect 17696 29668 18144 29696
rect 11241 29631 11299 29637
rect 11241 29628 11253 29631
rect 11020 29600 11253 29628
rect 11020 29588 11026 29600
rect 11241 29597 11253 29600
rect 11287 29628 11299 29631
rect 13541 29631 13599 29637
rect 11287 29600 12434 29628
rect 11287 29597 11299 29600
rect 11241 29591 11299 29597
rect 8076 29532 8708 29560
rect 9125 29563 9183 29569
rect 8076 29520 8082 29532
rect 9125 29529 9137 29563
rect 9171 29560 9183 29563
rect 10226 29560 10232 29572
rect 9171 29532 10232 29560
rect 9171 29529 9183 29532
rect 9125 29523 9183 29529
rect 10226 29520 10232 29532
rect 10284 29520 10290 29572
rect 12406 29560 12434 29600
rect 13541 29597 13553 29631
rect 13587 29597 13599 29631
rect 13541 29591 13599 29597
rect 13725 29631 13783 29637
rect 13725 29597 13737 29631
rect 13771 29628 13783 29631
rect 14458 29628 14464 29640
rect 13771 29600 14464 29628
rect 13771 29597 13783 29600
rect 13725 29591 13783 29597
rect 14458 29588 14464 29600
rect 14516 29588 14522 29640
rect 14826 29628 14832 29640
rect 14787 29600 14832 29628
rect 14826 29588 14832 29600
rect 14884 29588 14890 29640
rect 15120 29637 15148 29668
rect 15105 29631 15163 29637
rect 15105 29597 15117 29631
rect 15151 29597 15163 29631
rect 15105 29591 15163 29597
rect 15197 29631 15255 29637
rect 15197 29597 15209 29631
rect 15243 29597 15255 29631
rect 15473 29631 15531 29637
rect 15473 29628 15485 29631
rect 15197 29591 15255 29597
rect 15304 29600 15485 29628
rect 14369 29563 14427 29569
rect 14369 29560 14381 29563
rect 12406 29532 14381 29560
rect 14369 29529 14381 29532
rect 14415 29529 14427 29563
rect 14369 29523 14427 29529
rect 14918 29520 14924 29572
rect 14976 29560 14982 29572
rect 15212 29560 15240 29591
rect 14976 29532 15240 29560
rect 14976 29520 14982 29532
rect 13354 29492 13360 29504
rect 7484 29464 13360 29492
rect 5500 29452 5506 29464
rect 13354 29452 13360 29464
rect 13412 29452 13418 29504
rect 13725 29495 13783 29501
rect 13725 29461 13737 29495
rect 13771 29492 13783 29495
rect 14274 29492 14280 29504
rect 13771 29464 14280 29492
rect 13771 29461 13783 29464
rect 13725 29455 13783 29461
rect 14274 29452 14280 29464
rect 14332 29452 14338 29504
rect 14458 29452 14464 29504
rect 14516 29492 14522 29504
rect 15102 29492 15108 29504
rect 14516 29464 15108 29492
rect 14516 29452 14522 29464
rect 15102 29452 15108 29464
rect 15160 29492 15166 29504
rect 15304 29492 15332 29600
rect 15473 29597 15485 29600
rect 15519 29597 15531 29631
rect 15746 29628 15752 29640
rect 15707 29600 15752 29628
rect 15473 29591 15531 29597
rect 15746 29588 15752 29600
rect 15804 29588 15810 29640
rect 17696 29637 17724 29668
rect 18138 29656 18144 29668
rect 18196 29656 18202 29708
rect 18782 29696 18788 29708
rect 18524 29668 18788 29696
rect 17681 29631 17739 29637
rect 17681 29597 17693 29631
rect 17727 29597 17739 29631
rect 17681 29591 17739 29597
rect 17865 29631 17923 29637
rect 17865 29597 17877 29631
rect 17911 29597 17923 29631
rect 17865 29591 17923 29597
rect 17957 29631 18015 29637
rect 17957 29597 17969 29631
rect 18003 29628 18015 29631
rect 18230 29628 18236 29640
rect 18003 29600 18236 29628
rect 18003 29597 18015 29600
rect 17957 29591 18015 29597
rect 15160 29464 15332 29492
rect 17880 29492 17908 29591
rect 18230 29588 18236 29600
rect 18288 29588 18294 29640
rect 18524 29637 18552 29668
rect 18782 29656 18788 29668
rect 18840 29656 18846 29708
rect 19536 29696 19564 29736
rect 19978 29724 19984 29736
rect 20036 29724 20042 29776
rect 20162 29724 20168 29776
rect 20220 29764 20226 29776
rect 20717 29767 20775 29773
rect 20717 29764 20729 29767
rect 20220 29736 20729 29764
rect 20220 29724 20226 29736
rect 20717 29733 20729 29736
rect 20763 29733 20775 29767
rect 20824 29764 20852 29804
rect 24765 29801 24777 29835
rect 24811 29801 24823 29835
rect 24946 29832 24952 29844
rect 24907 29804 24952 29832
rect 24765 29795 24823 29801
rect 22094 29764 22100 29776
rect 20824 29736 22100 29764
rect 20717 29727 20775 29733
rect 22094 29724 22100 29736
rect 22152 29724 22158 29776
rect 23566 29724 23572 29776
rect 23624 29764 23630 29776
rect 24780 29764 24808 29795
rect 24946 29792 24952 29804
rect 25004 29792 25010 29844
rect 28445 29835 28503 29841
rect 28445 29801 28457 29835
rect 28491 29832 28503 29835
rect 29270 29832 29276 29844
rect 28491 29804 29276 29832
rect 28491 29801 28503 29804
rect 28445 29795 28503 29801
rect 29270 29792 29276 29804
rect 29328 29792 29334 29844
rect 29733 29835 29791 29841
rect 29733 29801 29745 29835
rect 29779 29832 29791 29835
rect 30190 29832 30196 29844
rect 29779 29804 30196 29832
rect 29779 29801 29791 29804
rect 29733 29795 29791 29801
rect 30190 29792 30196 29804
rect 30248 29792 30254 29844
rect 30558 29792 30564 29844
rect 30616 29832 30622 29844
rect 32033 29835 32091 29841
rect 32033 29832 32045 29835
rect 30616 29804 32045 29832
rect 30616 29792 30622 29804
rect 32033 29801 32045 29804
rect 32079 29801 32091 29835
rect 33226 29832 33232 29844
rect 32033 29795 32091 29801
rect 32876 29804 33232 29832
rect 25590 29764 25596 29776
rect 23624 29736 24532 29764
rect 24780 29736 25596 29764
rect 23624 29724 23630 29736
rect 20180 29696 20208 29724
rect 20898 29696 20904 29708
rect 19352 29668 19564 29696
rect 19628 29668 20208 29696
rect 20859 29668 20904 29696
rect 19352 29640 19380 29668
rect 18509 29631 18567 29637
rect 18509 29597 18521 29631
rect 18555 29597 18567 29631
rect 18509 29591 18567 29597
rect 18693 29631 18751 29637
rect 18693 29597 18705 29631
rect 18739 29628 18751 29631
rect 19334 29628 19340 29640
rect 18739 29600 19340 29628
rect 18739 29597 18751 29600
rect 18693 29591 18751 29597
rect 19334 29588 19340 29600
rect 19392 29588 19398 29640
rect 19628 29637 19656 29668
rect 20898 29656 20904 29668
rect 20956 29656 20962 29708
rect 23750 29696 23756 29708
rect 23711 29668 23756 29696
rect 23750 29656 23756 29668
rect 23808 29656 23814 29708
rect 23934 29696 23940 29708
rect 23895 29668 23940 29696
rect 23934 29656 23940 29668
rect 23992 29656 23998 29708
rect 19613 29631 19671 29637
rect 19613 29597 19625 29631
rect 19659 29597 19671 29631
rect 19613 29591 19671 29597
rect 19705 29631 19763 29637
rect 19705 29597 19717 29631
rect 19751 29597 19763 29631
rect 19705 29591 19763 29597
rect 19889 29631 19947 29637
rect 19889 29597 19901 29631
rect 19935 29597 19947 29631
rect 19889 29591 19947 29597
rect 18322 29492 18328 29504
rect 17880 29464 18328 29492
rect 15160 29452 15166 29464
rect 18322 29452 18328 29464
rect 18380 29492 18386 29504
rect 19429 29495 19487 29501
rect 19429 29492 19441 29495
rect 18380 29464 19441 29492
rect 18380 29452 18386 29464
rect 19429 29461 19441 29464
rect 19475 29461 19487 29495
rect 19720 29492 19748 29591
rect 19904 29560 19932 29591
rect 19978 29588 19984 29640
rect 20036 29628 20042 29640
rect 21361 29631 21419 29637
rect 21361 29628 21373 29631
rect 20036 29600 21373 29628
rect 20036 29588 20042 29600
rect 21361 29597 21373 29600
rect 21407 29597 21419 29631
rect 21361 29591 21419 29597
rect 21545 29631 21603 29637
rect 21545 29597 21557 29631
rect 21591 29628 21603 29631
rect 23474 29628 23480 29640
rect 21591 29600 23480 29628
rect 21591 29597 21603 29600
rect 21545 29591 21603 29597
rect 20070 29560 20076 29572
rect 19904 29532 20076 29560
rect 20070 29520 20076 29532
rect 20128 29520 20134 29572
rect 20346 29520 20352 29572
rect 20404 29560 20410 29572
rect 20441 29563 20499 29569
rect 20441 29560 20453 29563
rect 20404 29532 20453 29560
rect 20404 29520 20410 29532
rect 20441 29529 20453 29532
rect 20487 29560 20499 29563
rect 21453 29563 21511 29569
rect 21453 29560 21465 29563
rect 20487 29532 21465 29560
rect 20487 29529 20499 29532
rect 20441 29523 20499 29529
rect 21453 29529 21465 29532
rect 21499 29529 21511 29563
rect 21453 29523 21511 29529
rect 21560 29492 21588 29591
rect 23474 29588 23480 29600
rect 23532 29588 23538 29640
rect 23658 29628 23664 29640
rect 23619 29600 23664 29628
rect 23658 29588 23664 29600
rect 23716 29588 23722 29640
rect 23842 29588 23848 29640
rect 23900 29628 23906 29640
rect 24504 29628 24532 29736
rect 25590 29724 25596 29736
rect 25648 29764 25654 29776
rect 25648 29736 26234 29764
rect 25648 29724 25654 29736
rect 24578 29656 24584 29708
rect 24636 29696 24642 29708
rect 26050 29696 26056 29708
rect 24636 29668 24808 29696
rect 26011 29668 26056 29696
rect 24636 29656 24642 29668
rect 23900 29600 23945 29628
rect 24504 29600 24716 29628
rect 23900 29588 23906 29600
rect 24688 29572 24716 29600
rect 23382 29520 23388 29572
rect 23440 29560 23446 29572
rect 24581 29563 24639 29569
rect 23440 29532 24532 29560
rect 23440 29520 23446 29532
rect 19720 29464 21588 29492
rect 19429 29455 19487 29461
rect 22830 29452 22836 29504
rect 22888 29492 22894 29504
rect 23477 29495 23535 29501
rect 23477 29492 23489 29495
rect 22888 29464 23489 29492
rect 22888 29452 22894 29464
rect 23477 29461 23489 29464
rect 23523 29461 23535 29495
rect 24504 29492 24532 29532
rect 24581 29529 24593 29563
rect 24627 29560 24639 29563
rect 24670 29560 24676 29572
rect 24627 29532 24676 29560
rect 24627 29529 24639 29532
rect 24581 29523 24639 29529
rect 24670 29520 24676 29532
rect 24728 29520 24734 29572
rect 24780 29560 24808 29668
rect 26050 29656 26056 29668
rect 26108 29656 26114 29708
rect 26206 29696 26234 29736
rect 28350 29724 28356 29776
rect 28408 29764 28414 29776
rect 32876 29764 32904 29804
rect 33226 29792 33232 29804
rect 33284 29792 33290 29844
rect 28408 29736 30052 29764
rect 28408 29724 28414 29736
rect 28537 29699 28595 29705
rect 26206 29668 28488 29696
rect 25958 29628 25964 29640
rect 25919 29600 25964 29628
rect 25958 29588 25964 29600
rect 26016 29588 26022 29640
rect 27982 29588 27988 29640
rect 28040 29628 28046 29640
rect 28261 29631 28319 29637
rect 28261 29628 28273 29631
rect 28040 29600 28273 29628
rect 28040 29588 28046 29600
rect 28261 29597 28273 29600
rect 28307 29597 28319 29631
rect 28460 29628 28488 29668
rect 28537 29665 28549 29699
rect 28583 29696 28595 29699
rect 29178 29696 29184 29708
rect 28583 29668 29184 29696
rect 28583 29665 28595 29668
rect 28537 29659 28595 29665
rect 29178 29656 29184 29668
rect 29236 29656 29242 29708
rect 29730 29628 29736 29640
rect 28460 29600 29592 29628
rect 29691 29600 29736 29628
rect 28261 29591 28319 29597
rect 28718 29560 28724 29572
rect 24780 29532 28724 29560
rect 28718 29520 28724 29532
rect 28776 29520 28782 29572
rect 29564 29560 29592 29600
rect 29730 29588 29736 29600
rect 29788 29588 29794 29640
rect 30024 29637 30052 29736
rect 32048 29736 32904 29764
rect 30009 29631 30067 29637
rect 30009 29597 30021 29631
rect 30055 29597 30067 29631
rect 30009 29591 30067 29597
rect 31662 29560 31668 29572
rect 29564 29532 31668 29560
rect 31662 29520 31668 29532
rect 31720 29520 31726 29572
rect 24781 29495 24839 29501
rect 24781 29492 24793 29495
rect 24504 29464 24793 29492
rect 23477 29455 23535 29461
rect 24781 29461 24793 29464
rect 24827 29492 24839 29495
rect 25866 29492 25872 29504
rect 24827 29464 25872 29492
rect 24827 29461 24839 29464
rect 24781 29455 24839 29461
rect 25866 29452 25872 29464
rect 25924 29452 25930 29504
rect 26329 29495 26387 29501
rect 26329 29461 26341 29495
rect 26375 29492 26387 29495
rect 27706 29492 27712 29504
rect 26375 29464 27712 29492
rect 26375 29461 26387 29464
rect 26329 29455 26387 29461
rect 27706 29452 27712 29464
rect 27764 29452 27770 29504
rect 27798 29452 27804 29504
rect 27856 29492 27862 29504
rect 28077 29495 28135 29501
rect 28077 29492 28089 29495
rect 27856 29464 28089 29492
rect 27856 29452 27862 29464
rect 28077 29461 28089 29464
rect 28123 29461 28135 29495
rect 28077 29455 28135 29461
rect 29546 29452 29552 29504
rect 29604 29492 29610 29504
rect 29822 29492 29828 29504
rect 29604 29464 29828 29492
rect 29604 29452 29610 29464
rect 29822 29452 29828 29464
rect 29880 29492 29886 29504
rect 29917 29495 29975 29501
rect 29917 29492 29929 29495
rect 29880 29464 29929 29492
rect 29880 29452 29886 29464
rect 29917 29461 29929 29464
rect 29963 29492 29975 29495
rect 32048 29492 32076 29736
rect 32950 29724 32956 29776
rect 33008 29764 33014 29776
rect 33045 29767 33103 29773
rect 33045 29764 33057 29767
rect 33008 29736 33057 29764
rect 33008 29724 33014 29736
rect 33045 29733 33057 29736
rect 33091 29733 33103 29767
rect 33045 29727 33103 29733
rect 33060 29696 33088 29727
rect 32508 29668 33088 29696
rect 32214 29628 32220 29640
rect 32127 29600 32220 29628
rect 32214 29588 32220 29600
rect 32272 29588 32278 29640
rect 32398 29628 32404 29640
rect 32359 29600 32404 29628
rect 32398 29588 32404 29600
rect 32456 29588 32462 29640
rect 32508 29637 32536 29668
rect 32493 29631 32551 29637
rect 32493 29597 32505 29631
rect 32539 29597 32551 29631
rect 33134 29628 33140 29640
rect 33095 29600 33140 29628
rect 32493 29591 32551 29597
rect 33134 29588 33140 29600
rect 33192 29588 33198 29640
rect 33226 29588 33232 29640
rect 33284 29628 33290 29640
rect 33686 29628 33692 29640
rect 33284 29600 33692 29628
rect 33284 29588 33290 29600
rect 33686 29588 33692 29600
rect 33744 29588 33750 29640
rect 29963 29464 32076 29492
rect 32232 29492 32260 29588
rect 32953 29563 33011 29569
rect 32953 29529 32965 29563
rect 32999 29560 33011 29563
rect 33318 29560 33324 29572
rect 32999 29532 33324 29560
rect 32999 29529 33011 29532
rect 32953 29523 33011 29529
rect 33318 29520 33324 29532
rect 33376 29520 33382 29572
rect 33502 29492 33508 29504
rect 32232 29464 33508 29492
rect 29963 29461 29975 29464
rect 29917 29455 29975 29461
rect 33502 29452 33508 29464
rect 33560 29452 33566 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 5074 29248 5080 29300
rect 5132 29288 5138 29300
rect 5994 29288 6000 29300
rect 5132 29260 6000 29288
rect 5132 29248 5138 29260
rect 5994 29248 6000 29260
rect 6052 29248 6058 29300
rect 6362 29248 6368 29300
rect 6420 29288 6426 29300
rect 6549 29291 6607 29297
rect 6549 29288 6561 29291
rect 6420 29260 6561 29288
rect 6420 29248 6426 29260
rect 6549 29257 6561 29260
rect 6595 29257 6607 29291
rect 8386 29288 8392 29300
rect 6549 29251 6607 29257
rect 6748 29260 8248 29288
rect 8347 29260 8392 29288
rect 5166 29180 5172 29232
rect 5224 29220 5230 29232
rect 6748 29220 6776 29260
rect 8110 29220 8116 29232
rect 5224 29192 6776 29220
rect 6840 29192 8116 29220
rect 5224 29180 5230 29192
rect 4982 29152 4988 29164
rect 4943 29124 4988 29152
rect 4982 29112 4988 29124
rect 5040 29112 5046 29164
rect 5442 29152 5448 29164
rect 5403 29124 5448 29152
rect 5442 29112 5448 29124
rect 5500 29112 5506 29164
rect 5534 29112 5540 29164
rect 5592 29152 5598 29164
rect 6840 29161 6868 29192
rect 8110 29180 8116 29192
rect 8168 29180 8174 29232
rect 6825 29155 6883 29161
rect 6825 29152 6837 29155
rect 5592 29124 6837 29152
rect 5592 29112 5598 29124
rect 6825 29121 6837 29124
rect 6871 29121 6883 29155
rect 6825 29115 6883 29121
rect 6914 29112 6920 29164
rect 6972 29152 6978 29164
rect 8220 29161 8248 29260
rect 8386 29248 8392 29260
rect 8444 29248 8450 29300
rect 9306 29248 9312 29300
rect 9364 29288 9370 29300
rect 10318 29288 10324 29300
rect 9364 29260 10324 29288
rect 9364 29248 9370 29260
rect 10318 29248 10324 29260
rect 10376 29248 10382 29300
rect 18782 29288 18788 29300
rect 18743 29260 18788 29288
rect 18782 29248 18788 29260
rect 18840 29248 18846 29300
rect 19426 29288 19432 29300
rect 18984 29260 19432 29288
rect 14458 29220 14464 29232
rect 14200 29192 14464 29220
rect 14200 29161 14228 29192
rect 14458 29180 14464 29192
rect 14516 29180 14522 29232
rect 8205 29155 8263 29161
rect 6972 29124 7017 29152
rect 6972 29112 6978 29124
rect 8205 29121 8217 29155
rect 8251 29121 8263 29155
rect 14093 29155 14151 29161
rect 8205 29115 8263 29121
rect 8864 29124 10548 29152
rect 6086 29044 6092 29096
rect 6144 29084 6150 29096
rect 6733 29087 6791 29093
rect 6733 29084 6745 29087
rect 6144 29056 6745 29084
rect 6144 29044 6150 29056
rect 6733 29053 6745 29056
rect 6779 29053 6791 29087
rect 6733 29047 6791 29053
rect 7009 29087 7067 29093
rect 7009 29053 7021 29087
rect 7055 29084 7067 29087
rect 7742 29084 7748 29096
rect 7055 29056 7748 29084
rect 7055 29053 7067 29056
rect 7009 29047 7067 29053
rect 7742 29044 7748 29056
rect 7800 29044 7806 29096
rect 8021 29087 8079 29093
rect 8021 29053 8033 29087
rect 8067 29084 8079 29087
rect 8864 29084 8892 29124
rect 8067 29056 8892 29084
rect 8941 29087 8999 29093
rect 8067 29053 8079 29056
rect 8021 29047 8079 29053
rect 8941 29053 8953 29087
rect 8987 29053 8999 29087
rect 9214 29084 9220 29096
rect 9175 29056 9220 29084
rect 8941 29047 8999 29053
rect 5350 29016 5356 29028
rect 5311 28988 5356 29016
rect 5350 28976 5356 28988
rect 5408 28976 5414 29028
rect 7926 29016 7932 29028
rect 5460 28988 7932 29016
rect 5258 28908 5264 28960
rect 5316 28948 5322 28960
rect 5460 28948 5488 28988
rect 7926 28976 7932 28988
rect 7984 29016 7990 29028
rect 8956 29016 8984 29047
rect 9214 29044 9220 29056
rect 9272 29044 9278 29096
rect 7984 28988 8984 29016
rect 7984 28976 7990 28988
rect 10520 28957 10548 29124
rect 14093 29121 14105 29155
rect 14139 29121 14151 29155
rect 14093 29115 14151 29121
rect 14185 29155 14243 29161
rect 14185 29121 14197 29155
rect 14231 29121 14243 29155
rect 14185 29115 14243 29121
rect 14108 29084 14136 29115
rect 14274 29112 14280 29164
rect 14332 29152 14338 29164
rect 18984 29161 19012 29260
rect 19426 29248 19432 29260
rect 19484 29248 19490 29300
rect 20073 29291 20131 29297
rect 20073 29257 20085 29291
rect 20119 29288 20131 29291
rect 20254 29288 20260 29300
rect 20119 29260 20260 29288
rect 20119 29257 20131 29260
rect 20073 29251 20131 29257
rect 20254 29248 20260 29260
rect 20312 29248 20318 29300
rect 23750 29288 23756 29300
rect 23663 29260 23756 29288
rect 23750 29248 23756 29260
rect 23808 29248 23814 29300
rect 23934 29288 23940 29300
rect 23895 29260 23940 29288
rect 23934 29248 23940 29260
rect 23992 29248 23998 29300
rect 24762 29248 24768 29300
rect 24820 29248 24826 29300
rect 24854 29248 24860 29300
rect 24912 29288 24918 29300
rect 25777 29291 25835 29297
rect 25777 29288 25789 29291
rect 24912 29260 25789 29288
rect 24912 29248 24918 29260
rect 25777 29257 25789 29260
rect 25823 29257 25835 29291
rect 25777 29251 25835 29257
rect 25866 29248 25872 29300
rect 25924 29288 25930 29300
rect 28074 29288 28080 29300
rect 25924 29260 26234 29288
rect 28035 29260 28080 29288
rect 25924 29248 25930 29260
rect 22370 29220 22376 29232
rect 20548 29192 22376 29220
rect 14369 29155 14427 29161
rect 14369 29152 14381 29155
rect 14332 29124 14381 29152
rect 14332 29112 14338 29124
rect 14369 29121 14381 29124
rect 14415 29121 14427 29155
rect 14369 29115 14427 29121
rect 18969 29155 19027 29161
rect 18969 29121 18981 29155
rect 19015 29121 19027 29155
rect 18969 29115 19027 29121
rect 19150 29112 19156 29164
rect 19208 29152 19214 29164
rect 20257 29155 20315 29161
rect 19208 29124 19253 29152
rect 19208 29112 19214 29124
rect 20257 29121 20269 29155
rect 20303 29121 20315 29155
rect 20257 29115 20315 29121
rect 18598 29084 18604 29096
rect 14108 29056 18604 29084
rect 18598 29044 18604 29056
rect 18656 29044 18662 29096
rect 19061 29087 19119 29093
rect 19061 29053 19073 29087
rect 19107 29053 19119 29087
rect 19061 29047 19119 29053
rect 13814 28976 13820 29028
rect 13872 29016 13878 29028
rect 13909 29019 13967 29025
rect 13909 29016 13921 29019
rect 13872 28988 13921 29016
rect 13872 28976 13878 28988
rect 13909 28985 13921 28988
rect 13955 28985 13967 29019
rect 13909 28979 13967 28985
rect 14277 29019 14335 29025
rect 14277 28985 14289 29019
rect 14323 29016 14335 29019
rect 14918 29016 14924 29028
rect 14323 28988 14924 29016
rect 14323 28985 14335 28988
rect 14277 28979 14335 28985
rect 14918 28976 14924 28988
rect 14976 28976 14982 29028
rect 17402 28976 17408 29028
rect 17460 29016 17466 29028
rect 19076 29016 19104 29047
rect 19242 29044 19248 29096
rect 19300 29084 19306 29096
rect 20070 29084 20076 29096
rect 19300 29056 20076 29084
rect 19300 29044 19306 29056
rect 20070 29044 20076 29056
rect 20128 29044 20134 29096
rect 20272 29084 20300 29115
rect 20346 29112 20352 29164
rect 20404 29152 20410 29164
rect 20548 29161 20576 29192
rect 22370 29180 22376 29192
rect 22428 29180 22434 29232
rect 23658 29180 23664 29232
rect 23716 29180 23722 29232
rect 23768 29220 23796 29248
rect 24780 29220 24808 29248
rect 25590 29220 25596 29232
rect 23768 29192 25084 29220
rect 25551 29192 25596 29220
rect 20533 29155 20591 29161
rect 20404 29124 20449 29152
rect 20404 29112 20410 29124
rect 20533 29121 20545 29155
rect 20579 29121 20591 29155
rect 20533 29115 20591 29121
rect 20622 29112 20628 29164
rect 20680 29152 20686 29164
rect 20717 29155 20775 29161
rect 20717 29152 20729 29155
rect 20680 29124 20729 29152
rect 20680 29112 20686 29124
rect 20717 29121 20729 29124
rect 20763 29121 20775 29155
rect 23676 29152 23704 29180
rect 23676 29124 24072 29152
rect 20717 29115 20775 29121
rect 24044 29096 24072 29124
rect 24670 29112 24676 29164
rect 24728 29152 24734 29164
rect 24765 29155 24823 29161
rect 24765 29152 24777 29155
rect 24728 29124 24777 29152
rect 24728 29112 24734 29124
rect 24765 29121 24777 29124
rect 24811 29121 24823 29155
rect 24765 29115 24823 29121
rect 24857 29155 24915 29161
rect 24857 29121 24869 29155
rect 24903 29152 24915 29155
rect 24946 29152 24952 29164
rect 24903 29124 24952 29152
rect 24903 29121 24915 29124
rect 24857 29115 24915 29121
rect 24946 29112 24952 29124
rect 25004 29112 25010 29164
rect 25056 29161 25084 29192
rect 25590 29180 25596 29192
rect 25648 29180 25654 29232
rect 26206 29220 26234 29260
rect 28074 29248 28080 29260
rect 28132 29248 28138 29300
rect 26206 29192 28028 29220
rect 25041 29155 25099 29161
rect 25041 29121 25053 29155
rect 25087 29121 25099 29155
rect 25866 29152 25872 29164
rect 25827 29124 25872 29152
rect 25041 29115 25099 29121
rect 25866 29112 25872 29124
rect 25924 29112 25930 29164
rect 27801 29155 27859 29161
rect 27801 29152 27813 29155
rect 26206 29124 27813 29152
rect 21266 29084 21272 29096
rect 20272 29056 21272 29084
rect 21266 29044 21272 29056
rect 21324 29044 21330 29096
rect 22465 29087 22523 29093
rect 22465 29053 22477 29087
rect 22511 29084 22523 29087
rect 23385 29087 23443 29093
rect 23385 29084 23397 29087
rect 22511 29056 23397 29084
rect 22511 29053 22523 29056
rect 22465 29047 22523 29053
rect 23385 29053 23397 29056
rect 23431 29053 23443 29087
rect 23385 29047 23443 29053
rect 23569 29087 23627 29093
rect 23569 29053 23581 29087
rect 23615 29053 23627 29087
rect 23569 29047 23627 29053
rect 23661 29087 23719 29093
rect 23661 29053 23673 29087
rect 23707 29084 23719 29087
rect 23934 29084 23940 29096
rect 23707 29056 23940 29084
rect 23707 29053 23719 29056
rect 23661 29047 23719 29053
rect 20162 29016 20168 29028
rect 17460 28988 19012 29016
rect 19076 28988 20168 29016
rect 17460 28976 17466 28988
rect 5316 28920 5488 28948
rect 10505 28951 10563 28957
rect 5316 28908 5322 28920
rect 10505 28917 10517 28951
rect 10551 28948 10563 28951
rect 10594 28948 10600 28960
rect 10551 28920 10600 28948
rect 10551 28917 10563 28920
rect 10505 28911 10563 28917
rect 10594 28908 10600 28920
rect 10652 28908 10658 28960
rect 18984 28948 19012 28988
rect 20162 28976 20168 28988
rect 20220 28976 20226 29028
rect 20438 28976 20444 29028
rect 20496 29016 20502 29028
rect 22830 29016 22836 29028
rect 20496 28988 20541 29016
rect 22791 28988 22836 29016
rect 20496 28976 20502 28988
rect 22830 28976 22836 28988
rect 22888 28976 22894 29028
rect 23584 29016 23612 29047
rect 23934 29044 23940 29056
rect 23992 29044 23998 29096
rect 24026 29044 24032 29096
rect 24084 29084 24090 29096
rect 24486 29084 24492 29096
rect 24084 29056 24492 29084
rect 24084 29044 24090 29056
rect 24486 29044 24492 29056
rect 24544 29044 24550 29096
rect 24581 29087 24639 29093
rect 24581 29053 24593 29087
rect 24627 29084 24639 29087
rect 26050 29084 26056 29096
rect 24627 29056 26056 29084
rect 24627 29053 24639 29056
rect 24581 29047 24639 29053
rect 26050 29044 26056 29056
rect 26108 29084 26114 29096
rect 26206 29084 26234 29124
rect 27801 29121 27813 29124
rect 27847 29121 27859 29155
rect 27801 29115 27859 29121
rect 26108 29056 26234 29084
rect 27617 29087 27675 29093
rect 26108 29044 26114 29056
rect 27617 29053 27629 29087
rect 27663 29053 27675 29087
rect 27617 29047 27675 29053
rect 23584 28988 24256 29016
rect 19334 28948 19340 28960
rect 18984 28920 19340 28948
rect 19334 28908 19340 28920
rect 19392 28908 19398 28960
rect 22370 28908 22376 28960
rect 22428 28948 22434 28960
rect 22925 28951 22983 28957
rect 22925 28948 22937 28951
rect 22428 28920 22937 28948
rect 22428 28908 22434 28920
rect 22925 28917 22937 28920
rect 22971 28917 22983 28951
rect 24228 28948 24256 28988
rect 24302 28976 24308 29028
rect 24360 29016 24366 29028
rect 24949 29019 25007 29025
rect 24949 29016 24961 29019
rect 24360 28988 24961 29016
rect 24360 28976 24366 28988
rect 24949 28985 24961 28988
rect 24995 29016 25007 29019
rect 25593 29019 25651 29025
rect 25593 29016 25605 29019
rect 24995 28988 25605 29016
rect 24995 28985 25007 28988
rect 24949 28979 25007 28985
rect 25593 28985 25605 28988
rect 25639 28985 25651 29019
rect 27632 29016 27660 29047
rect 28000 29016 28028 29192
rect 28718 29152 28724 29164
rect 28679 29124 28724 29152
rect 28718 29112 28724 29124
rect 28776 29112 28782 29164
rect 28169 29087 28227 29093
rect 28169 29053 28181 29087
rect 28215 29084 28227 29087
rect 29178 29084 29184 29096
rect 28215 29056 29184 29084
rect 28215 29053 28227 29056
rect 28169 29047 28227 29053
rect 29178 29044 29184 29056
rect 29236 29044 29242 29096
rect 29270 29044 29276 29096
rect 29328 29084 29334 29096
rect 29328 29056 29373 29084
rect 29328 29044 29334 29056
rect 31110 29016 31116 29028
rect 27632 28988 27936 29016
rect 28000 28988 31116 29016
rect 25593 28979 25651 28985
rect 24854 28948 24860 28960
rect 24228 28920 24860 28948
rect 22925 28911 22983 28917
rect 24854 28908 24860 28920
rect 24912 28908 24918 28960
rect 27908 28948 27936 28988
rect 31110 28976 31116 28988
rect 31168 29016 31174 29028
rect 33318 29016 33324 29028
rect 31168 28988 33324 29016
rect 31168 28976 31174 28988
rect 33318 28976 33324 28988
rect 33376 28976 33382 29028
rect 29086 28948 29092 28960
rect 27908 28920 29092 28948
rect 29086 28908 29092 28920
rect 29144 28908 29150 28960
rect 29270 28908 29276 28960
rect 29328 28948 29334 28960
rect 29730 28948 29736 28960
rect 29328 28920 29736 28948
rect 29328 28908 29334 28920
rect 29730 28908 29736 28920
rect 29788 28948 29794 28960
rect 33226 28948 33232 28960
rect 29788 28920 33232 28948
rect 29788 28908 29794 28920
rect 33226 28908 33232 28920
rect 33284 28908 33290 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 9214 28744 9220 28756
rect 9175 28716 9220 28744
rect 9214 28704 9220 28716
rect 9272 28704 9278 28756
rect 10226 28704 10232 28756
rect 10284 28744 10290 28756
rect 10321 28747 10379 28753
rect 10321 28744 10333 28747
rect 10284 28716 10333 28744
rect 10284 28704 10290 28716
rect 10321 28713 10333 28716
rect 10367 28713 10379 28747
rect 11054 28744 11060 28756
rect 10321 28707 10379 28713
rect 10520 28716 11060 28744
rect 5534 28608 5540 28620
rect 5495 28580 5540 28608
rect 5534 28568 5540 28580
rect 5592 28568 5598 28620
rect 6086 28608 6092 28620
rect 6047 28580 6092 28608
rect 6086 28568 6092 28580
rect 6144 28568 6150 28620
rect 8294 28568 8300 28620
rect 8352 28608 8358 28620
rect 8352 28580 9628 28608
rect 8352 28568 8358 28580
rect 5721 28543 5779 28549
rect 5721 28509 5733 28543
rect 5767 28540 5779 28543
rect 6914 28540 6920 28552
rect 5767 28512 6920 28540
rect 5767 28509 5779 28512
rect 5721 28503 5779 28509
rect 6914 28500 6920 28512
rect 6972 28500 6978 28552
rect 9398 28540 9404 28552
rect 9359 28512 9404 28540
rect 9398 28500 9404 28512
rect 9456 28500 9462 28552
rect 9600 28549 9628 28580
rect 9585 28543 9643 28549
rect 9585 28509 9597 28543
rect 9631 28509 9643 28543
rect 9585 28503 9643 28509
rect 9674 28500 9680 28552
rect 9732 28549 9738 28552
rect 9732 28543 9761 28549
rect 9749 28509 9761 28543
rect 9858 28540 9864 28552
rect 9819 28512 9864 28540
rect 9732 28503 9761 28509
rect 9732 28500 9738 28503
rect 9858 28500 9864 28512
rect 9916 28500 9922 28552
rect 10318 28500 10324 28552
rect 10376 28540 10382 28552
rect 10520 28549 10548 28716
rect 11054 28704 11060 28716
rect 11112 28704 11118 28756
rect 14918 28744 14924 28756
rect 14879 28716 14924 28744
rect 14918 28704 14924 28716
rect 14976 28704 14982 28756
rect 18785 28747 18843 28753
rect 18785 28713 18797 28747
rect 18831 28744 18843 28747
rect 19242 28744 19248 28756
rect 18831 28716 19248 28744
rect 18831 28713 18843 28716
rect 18785 28707 18843 28713
rect 19242 28704 19248 28716
rect 19300 28704 19306 28756
rect 19889 28747 19947 28753
rect 19889 28713 19901 28747
rect 19935 28744 19947 28747
rect 19978 28744 19984 28756
rect 19935 28716 19984 28744
rect 19935 28713 19947 28716
rect 19889 28707 19947 28713
rect 19978 28704 19984 28716
rect 20036 28704 20042 28756
rect 20073 28747 20131 28753
rect 20073 28713 20085 28747
rect 20119 28744 20131 28747
rect 20438 28744 20444 28756
rect 20119 28716 20444 28744
rect 20119 28713 20131 28716
rect 20073 28707 20131 28713
rect 20438 28704 20444 28716
rect 20496 28704 20502 28756
rect 23934 28744 23940 28756
rect 23895 28716 23940 28744
rect 23934 28704 23940 28716
rect 23992 28704 23998 28756
rect 29914 28744 29920 28756
rect 28276 28716 29920 28744
rect 28276 28688 28304 28716
rect 29914 28704 29920 28716
rect 29972 28704 29978 28756
rect 10778 28676 10784 28688
rect 10704 28648 10784 28676
rect 10704 28617 10732 28648
rect 10778 28636 10784 28648
rect 10836 28636 10842 28688
rect 27338 28676 27344 28688
rect 24596 28648 27344 28676
rect 24596 28617 24624 28648
rect 27338 28636 27344 28648
rect 27396 28636 27402 28688
rect 28258 28676 28264 28688
rect 28171 28648 28264 28676
rect 28258 28636 28264 28648
rect 28316 28636 28322 28688
rect 29178 28636 29184 28688
rect 29236 28676 29242 28688
rect 30101 28679 30159 28685
rect 30101 28676 30113 28679
rect 29236 28648 30113 28676
rect 29236 28636 29242 28648
rect 30101 28645 30113 28648
rect 30147 28645 30159 28679
rect 33502 28676 33508 28688
rect 33463 28648 33508 28676
rect 30101 28639 30159 28645
rect 33502 28636 33508 28648
rect 33560 28636 33566 28688
rect 10689 28611 10747 28617
rect 10689 28577 10701 28611
rect 10735 28577 10747 28611
rect 10689 28571 10747 28577
rect 24581 28611 24639 28617
rect 24581 28577 24593 28611
rect 24627 28577 24639 28611
rect 24581 28571 24639 28577
rect 32953 28611 33011 28617
rect 32953 28577 32965 28611
rect 32999 28608 33011 28611
rect 34330 28608 34336 28620
rect 32999 28580 34336 28608
rect 32999 28577 33011 28580
rect 32953 28571 33011 28577
rect 34330 28568 34336 28580
rect 34388 28568 34394 28620
rect 10505 28543 10563 28549
rect 10505 28540 10517 28543
rect 10376 28512 10517 28540
rect 10376 28500 10382 28512
rect 10505 28509 10517 28512
rect 10551 28509 10563 28543
rect 10505 28503 10563 28509
rect 10594 28500 10600 28552
rect 10652 28540 10658 28552
rect 10781 28543 10839 28549
rect 10652 28512 10697 28540
rect 10652 28500 10658 28512
rect 10781 28509 10793 28543
rect 10827 28509 10839 28543
rect 10781 28503 10839 28509
rect 6822 28432 6828 28484
rect 6880 28472 6886 28484
rect 9493 28475 9551 28481
rect 9493 28472 9505 28475
rect 6880 28444 9505 28472
rect 6880 28432 6886 28444
rect 9493 28441 9505 28444
rect 9539 28472 9551 28475
rect 10796 28472 10824 28503
rect 14734 28500 14740 28552
rect 14792 28540 14798 28552
rect 14829 28543 14887 28549
rect 14829 28540 14841 28543
rect 14792 28512 14841 28540
rect 14792 28500 14798 28512
rect 14829 28509 14841 28512
rect 14875 28509 14887 28543
rect 14829 28503 14887 28509
rect 18414 28500 18420 28552
rect 18472 28540 18478 28552
rect 18693 28543 18751 28549
rect 18693 28540 18705 28543
rect 18472 28512 18705 28540
rect 18472 28500 18478 28512
rect 18693 28509 18705 28512
rect 18739 28540 18751 28543
rect 19521 28543 19579 28549
rect 19521 28540 19533 28543
rect 18739 28512 19533 28540
rect 18739 28509 18751 28512
rect 18693 28503 18751 28509
rect 19521 28509 19533 28512
rect 19567 28509 19579 28543
rect 22738 28540 22744 28552
rect 22699 28512 22744 28540
rect 19521 28503 19579 28509
rect 22738 28500 22744 28512
rect 22796 28500 22802 28552
rect 23566 28540 23572 28552
rect 23124 28512 23572 28540
rect 9539 28444 10824 28472
rect 9539 28441 9551 28444
rect 9493 28435 9551 28441
rect 19150 28432 19156 28484
rect 19208 28472 19214 28484
rect 19889 28475 19947 28481
rect 19889 28472 19901 28475
rect 19208 28444 19901 28472
rect 19208 28432 19214 28444
rect 19889 28441 19901 28444
rect 19935 28472 19947 28475
rect 23124 28472 23152 28512
rect 23566 28500 23572 28512
rect 23624 28500 23630 28552
rect 23845 28543 23903 28549
rect 23845 28509 23857 28543
rect 23891 28509 23903 28543
rect 23845 28503 23903 28509
rect 19935 28444 23152 28472
rect 23293 28475 23351 28481
rect 19935 28441 19947 28444
rect 19889 28435 19947 28441
rect 23293 28441 23305 28475
rect 23339 28441 23351 28475
rect 23860 28472 23888 28503
rect 24394 28500 24400 28552
rect 24452 28540 24458 28552
rect 24765 28543 24823 28549
rect 24765 28540 24777 28543
rect 24452 28512 24777 28540
rect 24452 28500 24458 28512
rect 24765 28509 24777 28512
rect 24811 28509 24823 28543
rect 24765 28503 24823 28509
rect 27706 28500 27712 28552
rect 27764 28540 27770 28552
rect 28629 28543 28687 28549
rect 28629 28540 28641 28543
rect 27764 28512 28641 28540
rect 27764 28500 27770 28512
rect 28629 28509 28641 28512
rect 28675 28509 28687 28543
rect 28629 28503 28687 28509
rect 33042 28500 33048 28552
rect 33100 28540 33106 28552
rect 33137 28543 33195 28549
rect 33137 28540 33149 28543
rect 33100 28512 33149 28540
rect 33100 28500 33106 28512
rect 33137 28509 33149 28512
rect 33183 28509 33195 28543
rect 33137 28503 33195 28509
rect 33410 28500 33416 28552
rect 33468 28540 33474 28552
rect 33505 28543 33563 28549
rect 33505 28540 33517 28543
rect 33468 28512 33517 28540
rect 33468 28500 33474 28512
rect 33505 28509 33517 28512
rect 33551 28509 33563 28543
rect 33505 28503 33563 28509
rect 33873 28543 33931 28549
rect 33873 28509 33885 28543
rect 33919 28509 33931 28543
rect 33873 28503 33931 28509
rect 24670 28472 24676 28484
rect 23860 28444 24676 28472
rect 23293 28435 23351 28441
rect 5718 28404 5724 28416
rect 5679 28376 5724 28404
rect 5718 28364 5724 28376
rect 5776 28364 5782 28416
rect 22554 28364 22560 28416
rect 22612 28404 22618 28416
rect 23308 28404 23336 28435
rect 24670 28432 24676 28444
rect 24728 28472 24734 28484
rect 24949 28475 25007 28481
rect 24949 28472 24961 28475
rect 24728 28444 24961 28472
rect 24728 28432 24734 28444
rect 24949 28441 24961 28444
rect 24995 28441 25007 28475
rect 24949 28435 25007 28441
rect 28445 28475 28503 28481
rect 28445 28441 28457 28475
rect 28491 28472 28503 28475
rect 28718 28472 28724 28484
rect 28491 28444 28724 28472
rect 28491 28441 28503 28444
rect 28445 28435 28503 28441
rect 28718 28432 28724 28444
rect 28776 28472 28782 28484
rect 29730 28472 29736 28484
rect 28776 28444 29592 28472
rect 29691 28444 29736 28472
rect 28776 28432 28782 28444
rect 29564 28416 29592 28444
rect 29730 28432 29736 28444
rect 29788 28432 29794 28484
rect 33318 28432 33324 28484
rect 33376 28472 33382 28484
rect 33888 28472 33916 28503
rect 33376 28444 33916 28472
rect 33376 28432 33382 28444
rect 25038 28404 25044 28416
rect 22612 28376 25044 28404
rect 22612 28364 22618 28376
rect 25038 28364 25044 28376
rect 25096 28364 25102 28416
rect 27614 28364 27620 28416
rect 27672 28404 27678 28416
rect 28350 28404 28356 28416
rect 27672 28376 28356 28404
rect 27672 28364 27678 28376
rect 28350 28364 28356 28376
rect 28408 28404 28414 28416
rect 28537 28407 28595 28413
rect 28537 28404 28549 28407
rect 28408 28376 28549 28404
rect 28408 28364 28414 28376
rect 28537 28373 28549 28376
rect 28583 28373 28595 28407
rect 28810 28404 28816 28416
rect 28771 28376 28816 28404
rect 28537 28367 28595 28373
rect 28810 28364 28816 28376
rect 28868 28364 28874 28416
rect 29546 28364 29552 28416
rect 29604 28404 29610 28416
rect 29933 28407 29991 28413
rect 29933 28404 29945 28407
rect 29604 28376 29945 28404
rect 29604 28364 29610 28376
rect 29933 28373 29945 28376
rect 29979 28373 29991 28407
rect 29933 28367 29991 28373
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 5258 28160 5264 28212
rect 5316 28209 5322 28212
rect 5316 28203 5335 28209
rect 5323 28169 5335 28203
rect 5316 28163 5335 28169
rect 9309 28203 9367 28209
rect 9309 28169 9321 28203
rect 9355 28200 9367 28203
rect 9858 28200 9864 28212
rect 9355 28172 9864 28200
rect 9355 28169 9367 28172
rect 9309 28163 9367 28169
rect 5316 28160 5322 28163
rect 9858 28160 9864 28172
rect 9916 28160 9922 28212
rect 19978 28160 19984 28212
rect 20036 28200 20042 28212
rect 24762 28200 24768 28212
rect 20036 28172 24624 28200
rect 24723 28172 24768 28200
rect 20036 28160 20042 28172
rect 5074 28132 5080 28144
rect 5035 28104 5080 28132
rect 5074 28092 5080 28104
rect 5132 28092 5138 28144
rect 6914 28092 6920 28144
rect 6972 28132 6978 28144
rect 9677 28135 9735 28141
rect 9677 28132 9689 28135
rect 6972 28104 9689 28132
rect 6972 28092 6978 28104
rect 9677 28101 9689 28104
rect 9723 28101 9735 28135
rect 9677 28095 9735 28101
rect 16025 28135 16083 28141
rect 16025 28101 16037 28135
rect 16071 28132 16083 28135
rect 16666 28132 16672 28144
rect 16071 28104 16672 28132
rect 16071 28101 16083 28104
rect 16025 28095 16083 28101
rect 16666 28092 16672 28104
rect 16724 28092 16730 28144
rect 22554 28132 22560 28144
rect 22515 28104 22560 28132
rect 22554 28092 22560 28104
rect 22612 28092 22618 28144
rect 24596 28141 24624 28172
rect 24762 28160 24768 28172
rect 24820 28160 24826 28212
rect 29086 28200 29092 28212
rect 29047 28172 29092 28200
rect 29086 28160 29092 28172
rect 29144 28160 29150 28212
rect 29457 28203 29515 28209
rect 29457 28169 29469 28203
rect 29503 28200 29515 28203
rect 29914 28200 29920 28212
rect 29503 28172 29920 28200
rect 29503 28169 29515 28172
rect 29457 28163 29515 28169
rect 29914 28160 29920 28172
rect 29972 28200 29978 28212
rect 31205 28203 31263 28209
rect 31205 28200 31217 28203
rect 29972 28172 31217 28200
rect 29972 28160 29978 28172
rect 31205 28169 31217 28172
rect 31251 28169 31263 28203
rect 31205 28163 31263 28169
rect 24581 28135 24639 28141
rect 24581 28101 24593 28135
rect 24627 28101 24639 28135
rect 33042 28132 33048 28144
rect 24581 28095 24639 28101
rect 31680 28104 33048 28132
rect 5626 28024 5632 28076
rect 5684 28064 5690 28076
rect 6822 28064 6828 28076
rect 5684 28036 6828 28064
rect 5684 28024 5690 28036
rect 6822 28024 6828 28036
rect 6880 28064 6886 28076
rect 7561 28067 7619 28073
rect 7561 28064 7573 28067
rect 6880 28036 7573 28064
rect 6880 28024 6886 28036
rect 7561 28033 7573 28036
rect 7607 28033 7619 28067
rect 7561 28027 7619 28033
rect 8386 28024 8392 28076
rect 8444 28064 8450 28076
rect 9493 28067 9551 28073
rect 9493 28064 9505 28067
rect 8444 28036 9505 28064
rect 8444 28024 8450 28036
rect 9493 28033 9505 28036
rect 9539 28033 9551 28067
rect 9493 28027 9551 28033
rect 9769 28067 9827 28073
rect 9769 28033 9781 28067
rect 9815 28064 9827 28067
rect 10318 28064 10324 28076
rect 9815 28036 10324 28064
rect 9815 28033 9827 28036
rect 9769 28027 9827 28033
rect 10318 28024 10324 28036
rect 10376 28024 10382 28076
rect 15841 28067 15899 28073
rect 15841 28033 15853 28067
rect 15887 28064 15899 28067
rect 16117 28067 16175 28073
rect 15887 28036 16068 28064
rect 15887 28033 15899 28036
rect 15841 28027 15899 28033
rect 16040 28008 16068 28036
rect 16117 28033 16129 28067
rect 16163 28064 16175 28067
rect 16482 28064 16488 28076
rect 16163 28036 16488 28064
rect 16163 28033 16175 28036
rect 16117 28027 16175 28033
rect 16482 28024 16488 28036
rect 16540 28024 16546 28076
rect 16758 28024 16764 28076
rect 16816 28064 16822 28076
rect 16945 28067 17003 28073
rect 16945 28064 16957 28067
rect 16816 28036 16957 28064
rect 16816 28024 16822 28036
rect 16945 28033 16957 28036
rect 16991 28033 17003 28067
rect 22186 28064 22192 28076
rect 22147 28036 22192 28064
rect 16945 28027 17003 28033
rect 22186 28024 22192 28036
rect 22244 28024 22250 28076
rect 22370 28064 22376 28076
rect 22331 28036 22376 28064
rect 22370 28024 22376 28036
rect 22428 28024 22434 28076
rect 24394 28064 24400 28076
rect 24355 28036 24400 28064
rect 24394 28024 24400 28036
rect 24452 28024 24458 28076
rect 27614 28024 27620 28076
rect 27672 28064 27678 28076
rect 28166 28064 28172 28076
rect 27672 28036 28172 28064
rect 27672 28024 27678 28036
rect 28166 28024 28172 28036
rect 28224 28024 28230 28076
rect 28442 28064 28448 28076
rect 28403 28036 28448 28064
rect 28442 28024 28448 28036
rect 28500 28024 28506 28076
rect 28629 28067 28687 28073
rect 28629 28033 28641 28067
rect 28675 28064 28687 28067
rect 28810 28064 28816 28076
rect 28675 28036 28816 28064
rect 28675 28033 28687 28036
rect 28629 28027 28687 28033
rect 28810 28024 28816 28036
rect 28868 28024 28874 28076
rect 29270 28064 29276 28076
rect 29231 28036 29276 28064
rect 29270 28024 29276 28036
rect 29328 28024 29334 28076
rect 29546 28064 29552 28076
rect 29507 28036 29552 28064
rect 29546 28024 29552 28036
rect 29604 28024 29610 28076
rect 31110 28024 31116 28076
rect 31168 28064 31174 28076
rect 31680 28073 31708 28104
rect 33042 28092 33048 28104
rect 33100 28132 33106 28144
rect 33100 28104 34468 28132
rect 33100 28092 33106 28104
rect 31389 28067 31447 28073
rect 31389 28064 31401 28067
rect 31168 28036 31401 28064
rect 31168 28024 31174 28036
rect 31389 28033 31401 28036
rect 31435 28033 31447 28067
rect 31389 28027 31447 28033
rect 31481 28067 31539 28073
rect 31481 28033 31493 28067
rect 31527 28033 31539 28067
rect 31481 28027 31539 28033
rect 31665 28067 31723 28073
rect 31665 28033 31677 28067
rect 31711 28033 31723 28067
rect 31665 28027 31723 28033
rect 16022 27956 16028 28008
rect 16080 27956 16086 28008
rect 22094 27888 22100 27940
rect 22152 27928 22158 27940
rect 22189 27931 22247 27937
rect 22189 27928 22201 27931
rect 22152 27900 22201 27928
rect 22152 27888 22158 27900
rect 22189 27897 22201 27900
rect 22235 27897 22247 27931
rect 22189 27891 22247 27897
rect 5166 27820 5172 27872
rect 5224 27860 5230 27872
rect 5261 27863 5319 27869
rect 5261 27860 5273 27863
rect 5224 27832 5273 27860
rect 5224 27820 5230 27832
rect 5261 27829 5273 27832
rect 5307 27829 5319 27863
rect 5442 27860 5448 27872
rect 5403 27832 5448 27860
rect 5261 27823 5319 27829
rect 5442 27820 5448 27832
rect 5500 27820 5506 27872
rect 7742 27860 7748 27872
rect 7703 27832 7748 27860
rect 7742 27820 7748 27832
rect 7800 27820 7806 27872
rect 15657 27863 15715 27869
rect 15657 27829 15669 27863
rect 15703 27860 15715 27863
rect 15746 27860 15752 27872
rect 15703 27832 15752 27860
rect 15703 27829 15715 27832
rect 15657 27823 15715 27829
rect 15746 27820 15752 27832
rect 15804 27820 15810 27872
rect 17034 27860 17040 27872
rect 16995 27832 17040 27860
rect 17034 27820 17040 27832
rect 17092 27820 17098 27872
rect 27985 27863 28043 27869
rect 27985 27829 27997 27863
rect 28031 27860 28043 27863
rect 28166 27860 28172 27872
rect 28031 27832 28172 27860
rect 28031 27829 28043 27832
rect 27985 27823 28043 27829
rect 28166 27820 28172 27832
rect 28224 27820 28230 27872
rect 31404 27860 31432 28027
rect 31496 27940 31524 28027
rect 31846 28024 31852 28076
rect 31904 28064 31910 28076
rect 32309 28067 32367 28073
rect 32309 28064 32321 28067
rect 31904 28036 32321 28064
rect 31904 28024 31910 28036
rect 32309 28033 32321 28036
rect 32355 28033 32367 28067
rect 32309 28027 32367 28033
rect 32493 28067 32551 28073
rect 32493 28033 32505 28067
rect 32539 28033 32551 28067
rect 33410 28064 33416 28076
rect 33371 28036 33416 28064
rect 32493 28027 32551 28033
rect 31573 27999 31631 28005
rect 31573 27965 31585 27999
rect 31619 27965 31631 27999
rect 31573 27959 31631 27965
rect 31478 27888 31484 27940
rect 31536 27888 31542 27940
rect 31588 27928 31616 27959
rect 31754 27956 31760 28008
rect 31812 27996 31818 28008
rect 32508 27996 32536 28027
rect 33410 28024 33416 28036
rect 33468 28024 33474 28076
rect 33597 28067 33655 28073
rect 33597 28033 33609 28067
rect 33643 28033 33655 28067
rect 33597 28027 33655 28033
rect 31812 27968 32536 27996
rect 31812 27956 31818 27968
rect 33134 27956 33140 28008
rect 33192 27996 33198 28008
rect 33612 27996 33640 28027
rect 33686 28024 33692 28076
rect 33744 28064 33750 28076
rect 34057 28067 34115 28073
rect 34057 28064 34069 28067
rect 33744 28036 34069 28064
rect 33744 28024 33750 28036
rect 34057 28033 34069 28036
rect 34103 28033 34115 28067
rect 34330 28064 34336 28076
rect 34291 28036 34336 28064
rect 34057 28027 34115 28033
rect 34330 28024 34336 28036
rect 34388 28024 34394 28076
rect 34440 28073 34468 28104
rect 34425 28067 34483 28073
rect 34425 28033 34437 28067
rect 34471 28033 34483 28067
rect 34425 28027 34483 28033
rect 33778 27996 33784 28008
rect 33192 27968 33640 27996
rect 33739 27968 33784 27996
rect 33192 27956 33198 27968
rect 33778 27956 33784 27968
rect 33836 27956 33842 28008
rect 33042 27928 33048 27940
rect 31588 27900 33048 27928
rect 33042 27888 33048 27900
rect 33100 27888 33106 27940
rect 32030 27860 32036 27872
rect 31404 27832 32036 27860
rect 32030 27820 32036 27832
rect 32088 27820 32094 27872
rect 32306 27860 32312 27872
rect 32267 27832 32312 27860
rect 32306 27820 32312 27832
rect 32364 27820 32370 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 19352 27628 19932 27656
rect 4341 27591 4399 27597
rect 4341 27557 4353 27591
rect 4387 27588 4399 27591
rect 5718 27588 5724 27600
rect 4387 27560 5724 27588
rect 4387 27557 4399 27560
rect 4341 27551 4399 27557
rect 5718 27548 5724 27560
rect 5776 27548 5782 27600
rect 6914 27548 6920 27600
rect 6972 27588 6978 27600
rect 7193 27591 7251 27597
rect 7193 27588 7205 27591
rect 6972 27560 7205 27588
rect 6972 27548 6978 27560
rect 7193 27557 7205 27560
rect 7239 27557 7251 27591
rect 7193 27551 7251 27557
rect 18138 27548 18144 27600
rect 18196 27588 18202 27600
rect 19352 27588 19380 27628
rect 18196 27560 19380 27588
rect 18196 27548 18202 27560
rect 19426 27548 19432 27600
rect 19484 27588 19490 27600
rect 19797 27591 19855 27597
rect 19797 27588 19809 27591
rect 19484 27560 19809 27588
rect 19484 27548 19490 27560
rect 19797 27557 19809 27560
rect 19843 27557 19855 27591
rect 19904 27588 19932 27628
rect 29546 27616 29552 27668
rect 29604 27656 29610 27668
rect 32125 27659 32183 27665
rect 32125 27656 32137 27659
rect 29604 27628 32137 27656
rect 29604 27616 29610 27628
rect 32125 27625 32137 27628
rect 32171 27625 32183 27659
rect 33410 27656 33416 27668
rect 32125 27619 32183 27625
rect 32784 27628 33416 27656
rect 26234 27588 26240 27600
rect 19904 27560 26240 27588
rect 19797 27551 19855 27557
rect 26234 27548 26240 27560
rect 26292 27548 26298 27600
rect 27338 27548 27344 27600
rect 27396 27588 27402 27600
rect 32674 27588 32680 27600
rect 27396 27560 32680 27588
rect 27396 27548 27402 27560
rect 4522 27520 4528 27532
rect 4483 27492 4528 27520
rect 4522 27480 4528 27492
rect 4580 27480 4586 27532
rect 14366 27480 14372 27532
rect 14424 27520 14430 27532
rect 14829 27523 14887 27529
rect 14829 27520 14841 27523
rect 14424 27492 14841 27520
rect 14424 27480 14430 27492
rect 14829 27489 14841 27492
rect 14875 27520 14887 27523
rect 22738 27520 22744 27532
rect 14875 27492 22744 27520
rect 14875 27489 14887 27492
rect 14829 27483 14887 27489
rect 22738 27480 22744 27492
rect 22796 27480 22802 27532
rect 24394 27480 24400 27532
rect 24452 27520 24458 27532
rect 25409 27523 25467 27529
rect 25409 27520 25421 27523
rect 24452 27492 25421 27520
rect 24452 27480 24458 27492
rect 4249 27455 4307 27461
rect 4249 27421 4261 27455
rect 4295 27421 4307 27455
rect 7098 27452 7104 27464
rect 7059 27424 7104 27452
rect 4249 27415 4307 27421
rect 4264 27384 4292 27415
rect 7098 27412 7104 27424
rect 7156 27412 7162 27464
rect 14274 27412 14280 27464
rect 14332 27452 14338 27464
rect 14458 27452 14464 27464
rect 14332 27424 14464 27452
rect 14332 27412 14338 27424
rect 14458 27412 14464 27424
rect 14516 27412 14522 27464
rect 14734 27452 14740 27464
rect 14695 27424 14740 27452
rect 14734 27412 14740 27424
rect 14792 27412 14798 27464
rect 15470 27412 15476 27464
rect 15528 27452 15534 27464
rect 15933 27455 15991 27461
rect 15933 27452 15945 27455
rect 15528 27424 15945 27452
rect 15528 27412 15534 27424
rect 15933 27421 15945 27424
rect 15979 27421 15991 27455
rect 15933 27415 15991 27421
rect 16209 27455 16267 27461
rect 16209 27421 16221 27455
rect 16255 27452 16267 27455
rect 16850 27452 16856 27464
rect 16255 27424 16856 27452
rect 16255 27421 16267 27424
rect 16209 27415 16267 27421
rect 16850 27412 16856 27424
rect 16908 27412 16914 27464
rect 18233 27455 18291 27461
rect 18233 27421 18245 27455
rect 18279 27421 18291 27455
rect 18506 27452 18512 27464
rect 18467 27424 18512 27452
rect 18233 27415 18291 27421
rect 4614 27384 4620 27396
rect 4264 27356 4620 27384
rect 4614 27344 4620 27356
rect 4672 27384 4678 27396
rect 5442 27384 5448 27396
rect 4672 27356 5448 27384
rect 4672 27344 4678 27356
rect 5442 27344 5448 27356
rect 5500 27344 5506 27396
rect 18248 27384 18276 27415
rect 18506 27412 18512 27424
rect 18564 27412 18570 27464
rect 19429 27455 19487 27461
rect 19429 27421 19441 27455
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 19583 27455 19641 27461
rect 19583 27421 19595 27455
rect 19629 27452 19641 27455
rect 19978 27452 19984 27464
rect 19629 27424 19984 27452
rect 19629 27421 19641 27424
rect 19583 27415 19641 27421
rect 18690 27384 18696 27396
rect 18248 27356 18696 27384
rect 18690 27344 18696 27356
rect 18748 27344 18754 27396
rect 19444 27384 19472 27415
rect 19978 27412 19984 27424
rect 20036 27412 20042 27464
rect 22462 27412 22468 27464
rect 22520 27452 22526 27464
rect 24026 27452 24032 27464
rect 22520 27424 24032 27452
rect 22520 27412 22526 27424
rect 24026 27412 24032 27424
rect 24084 27452 24090 27464
rect 24780 27461 24808 27492
rect 25409 27489 25421 27492
rect 25455 27489 25467 27523
rect 28442 27520 28448 27532
rect 28403 27492 28448 27520
rect 25409 27483 25467 27489
rect 28442 27480 28448 27492
rect 28500 27480 28506 27532
rect 24581 27455 24639 27461
rect 24581 27452 24593 27455
rect 24084 27424 24593 27452
rect 24084 27412 24090 27424
rect 24581 27421 24593 27424
rect 24627 27421 24639 27455
rect 24581 27415 24639 27421
rect 24765 27455 24823 27461
rect 24765 27421 24777 27455
rect 24811 27421 24823 27455
rect 25314 27452 25320 27464
rect 25275 27424 25320 27452
rect 24765 27415 24823 27421
rect 25314 27412 25320 27424
rect 25372 27412 25378 27464
rect 25501 27455 25559 27461
rect 25501 27421 25513 27455
rect 25547 27421 25559 27455
rect 25501 27415 25559 27421
rect 20622 27384 20628 27396
rect 19444 27356 20628 27384
rect 20622 27344 20628 27356
rect 20680 27344 20686 27396
rect 25516 27384 25544 27415
rect 27706 27412 27712 27464
rect 27764 27452 27770 27464
rect 28169 27455 28227 27461
rect 28169 27452 28181 27455
rect 27764 27424 28181 27452
rect 27764 27412 27770 27424
rect 28169 27421 28181 27424
rect 28215 27421 28227 27455
rect 28169 27415 28227 27421
rect 28258 27412 28264 27464
rect 28316 27452 28322 27464
rect 28573 27455 28631 27461
rect 28316 27424 28488 27452
rect 28316 27412 28322 27424
rect 24596 27356 26234 27384
rect 4525 27319 4583 27325
rect 4525 27285 4537 27319
rect 4571 27316 4583 27319
rect 4706 27316 4712 27328
rect 4571 27288 4712 27316
rect 4571 27285 4583 27288
rect 4525 27279 4583 27285
rect 4706 27276 4712 27288
rect 4764 27276 4770 27328
rect 17218 27276 17224 27328
rect 17276 27316 17282 27328
rect 17313 27319 17371 27325
rect 17313 27316 17325 27319
rect 17276 27288 17325 27316
rect 17276 27276 17282 27288
rect 17313 27285 17325 27288
rect 17359 27285 17371 27319
rect 18046 27316 18052 27328
rect 18007 27288 18052 27316
rect 17313 27279 17371 27285
rect 18046 27276 18052 27288
rect 18104 27276 18110 27328
rect 18414 27316 18420 27328
rect 18375 27288 18420 27316
rect 18414 27276 18420 27288
rect 18472 27276 18478 27328
rect 19334 27276 19340 27328
rect 19392 27316 19398 27328
rect 24596 27316 24624 27356
rect 24762 27316 24768 27328
rect 19392 27288 24624 27316
rect 24723 27288 24768 27316
rect 19392 27276 19398 27288
rect 24762 27276 24768 27288
rect 24820 27276 24826 27328
rect 26206 27316 26234 27356
rect 27614 27344 27620 27396
rect 27672 27384 27678 27396
rect 28350 27384 28356 27396
rect 27672 27356 28356 27384
rect 27672 27344 27678 27356
rect 28350 27344 28356 27356
rect 28408 27344 28414 27396
rect 28460 27393 28488 27424
rect 28573 27421 28585 27455
rect 28619 27452 28631 27455
rect 28718 27452 28724 27464
rect 28619 27424 28724 27452
rect 28619 27421 28631 27424
rect 28573 27415 28631 27421
rect 28718 27412 28724 27424
rect 28776 27412 28782 27464
rect 31220 27461 31248 27560
rect 32674 27548 32680 27560
rect 32732 27548 32738 27600
rect 31478 27480 31484 27532
rect 31536 27520 31542 27532
rect 31573 27523 31631 27529
rect 31573 27520 31585 27523
rect 31536 27492 31585 27520
rect 31536 27480 31542 27492
rect 31573 27489 31585 27492
rect 31619 27520 31631 27523
rect 32784 27520 32812 27628
rect 33410 27616 33416 27628
rect 33468 27616 33474 27668
rect 34057 27591 34115 27597
rect 34057 27588 34069 27591
rect 31619 27492 32812 27520
rect 31619 27489 31631 27492
rect 31573 27483 31631 27489
rect 31205 27455 31263 27461
rect 31205 27421 31217 27455
rect 31251 27421 31263 27455
rect 32030 27452 32036 27464
rect 31991 27424 32036 27452
rect 31205 27415 31263 27421
rect 32030 27412 32036 27424
rect 32088 27412 32094 27464
rect 32677 27455 32735 27461
rect 32677 27421 32689 27455
rect 32723 27452 32735 27455
rect 32784 27452 32812 27492
rect 33336 27560 34069 27588
rect 32950 27452 32956 27464
rect 32723 27424 32812 27452
rect 32911 27424 32956 27452
rect 32723 27421 32735 27424
rect 32677 27415 32735 27421
rect 32950 27412 32956 27424
rect 33008 27412 33014 27464
rect 33042 27412 33048 27464
rect 33100 27452 33106 27464
rect 33336 27461 33364 27560
rect 34057 27557 34069 27560
rect 34103 27557 34115 27591
rect 34057 27551 34115 27557
rect 34072 27492 34284 27520
rect 34072 27461 34100 27492
rect 33321 27455 33379 27461
rect 33321 27452 33333 27455
rect 33100 27424 33333 27452
rect 33100 27412 33106 27424
rect 33321 27421 33333 27424
rect 33367 27421 33379 27455
rect 33321 27415 33379 27421
rect 34057 27455 34115 27461
rect 34057 27421 34069 27455
rect 34103 27421 34115 27455
rect 34057 27415 34115 27421
rect 34149 27455 34207 27461
rect 34149 27421 34161 27455
rect 34195 27421 34207 27455
rect 34149 27415 34207 27421
rect 28445 27387 28503 27393
rect 28445 27353 28457 27387
rect 28491 27353 28503 27387
rect 28445 27347 28503 27353
rect 31021 27387 31079 27393
rect 31021 27353 31033 27387
rect 31067 27384 31079 27387
rect 32306 27384 32312 27396
rect 31067 27356 32312 27384
rect 31067 27353 31079 27356
rect 31021 27347 31079 27353
rect 32306 27344 32312 27356
rect 32364 27344 32370 27396
rect 32766 27344 32772 27396
rect 32824 27384 32830 27396
rect 34164 27384 34192 27415
rect 32824 27356 34192 27384
rect 32824 27344 32830 27356
rect 31386 27316 31392 27328
rect 26206 27288 31392 27316
rect 31386 27276 31392 27288
rect 31444 27316 31450 27328
rect 31662 27316 31668 27328
rect 31444 27288 31668 27316
rect 31444 27276 31450 27288
rect 31662 27276 31668 27288
rect 31720 27276 31726 27328
rect 32324 27316 32352 27344
rect 33042 27316 33048 27328
rect 32324 27288 33048 27316
rect 33042 27276 33048 27288
rect 33100 27316 33106 27328
rect 34256 27316 34284 27492
rect 33100 27288 34284 27316
rect 33100 27276 33106 27288
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 16114 27072 16120 27124
rect 16172 27112 16178 27124
rect 18138 27112 18144 27124
rect 16172 27084 18144 27112
rect 16172 27072 16178 27084
rect 18138 27072 18144 27084
rect 18196 27072 18202 27124
rect 18233 27115 18291 27121
rect 18233 27081 18245 27115
rect 18279 27112 18291 27115
rect 18414 27112 18420 27124
rect 18279 27084 18420 27112
rect 18279 27081 18291 27084
rect 18233 27075 18291 27081
rect 18414 27072 18420 27084
rect 18472 27072 18478 27124
rect 22005 27115 22063 27121
rect 22005 27081 22017 27115
rect 22051 27112 22063 27115
rect 22186 27112 22192 27124
rect 22051 27084 22192 27112
rect 22051 27081 22063 27084
rect 22005 27075 22063 27081
rect 22186 27072 22192 27084
rect 22244 27072 22250 27124
rect 22373 27115 22431 27121
rect 22373 27081 22385 27115
rect 22419 27112 22431 27115
rect 23382 27112 23388 27124
rect 22419 27084 23388 27112
rect 22419 27081 22431 27084
rect 22373 27075 22431 27081
rect 23382 27072 23388 27084
rect 23440 27072 23446 27124
rect 25314 27072 25320 27124
rect 25372 27112 25378 27124
rect 25593 27115 25651 27121
rect 25593 27112 25605 27115
rect 25372 27084 25605 27112
rect 25372 27072 25378 27084
rect 25593 27081 25605 27084
rect 25639 27112 25651 27115
rect 28718 27112 28724 27124
rect 25639 27084 28724 27112
rect 25639 27081 25651 27084
rect 25593 27075 25651 27081
rect 28718 27072 28724 27084
rect 28776 27072 28782 27124
rect 32677 27115 32735 27121
rect 32677 27081 32689 27115
rect 32723 27112 32735 27115
rect 32950 27112 32956 27124
rect 32723 27084 32956 27112
rect 32723 27081 32735 27084
rect 32677 27075 32735 27081
rect 32950 27072 32956 27084
rect 33008 27072 33014 27124
rect 5074 27044 5080 27056
rect 3160 27016 5080 27044
rect 3160 26985 3188 27016
rect 5074 27004 5080 27016
rect 5132 27004 5138 27056
rect 15838 27044 15844 27056
rect 15799 27016 15844 27044
rect 15838 27004 15844 27016
rect 15896 27004 15902 27056
rect 15930 27004 15936 27056
rect 15988 27044 15994 27056
rect 16025 27047 16083 27053
rect 16025 27044 16037 27047
rect 15988 27016 16037 27044
rect 15988 27004 15994 27016
rect 16025 27013 16037 27016
rect 16071 27044 16083 27047
rect 17120 27047 17178 27053
rect 16071 27016 17080 27044
rect 16071 27013 16083 27016
rect 16025 27007 16083 27013
rect 3145 26979 3203 26985
rect 3145 26945 3157 26979
rect 3191 26945 3203 26979
rect 4614 26976 4620 26988
rect 4575 26948 4620 26976
rect 3145 26939 3203 26945
rect 4614 26936 4620 26948
rect 4672 26936 4678 26988
rect 4893 26979 4951 26985
rect 4893 26945 4905 26979
rect 4939 26976 4951 26979
rect 5626 26976 5632 26988
rect 4939 26948 5632 26976
rect 4939 26945 4951 26948
rect 4893 26939 4951 26945
rect 5626 26936 5632 26948
rect 5684 26936 5690 26988
rect 12437 26979 12495 26985
rect 12437 26945 12449 26979
rect 12483 26976 12495 26979
rect 13814 26976 13820 26988
rect 12483 26948 13820 26976
rect 12483 26945 12495 26948
rect 12437 26939 12495 26945
rect 13814 26936 13820 26948
rect 13872 26936 13878 26988
rect 13909 26979 13967 26985
rect 13909 26945 13921 26979
rect 13955 26945 13967 26979
rect 14274 26976 14280 26988
rect 14235 26948 14280 26976
rect 13909 26939 13967 26945
rect 3053 26911 3111 26917
rect 3053 26877 3065 26911
rect 3099 26908 3111 26911
rect 3513 26911 3571 26917
rect 3099 26880 3188 26908
rect 3099 26877 3111 26880
rect 3053 26871 3111 26877
rect 3160 26852 3188 26880
rect 3513 26877 3525 26911
rect 3559 26908 3571 26911
rect 4522 26908 4528 26920
rect 3559 26880 4528 26908
rect 3559 26877 3571 26880
rect 3513 26871 3571 26877
rect 4522 26868 4528 26880
rect 4580 26908 4586 26920
rect 4801 26911 4859 26917
rect 4801 26908 4813 26911
rect 4580 26880 4813 26908
rect 4580 26868 4586 26880
rect 4801 26877 4813 26880
rect 4847 26877 4859 26911
rect 4801 26871 4859 26877
rect 12253 26911 12311 26917
rect 12253 26877 12265 26911
rect 12299 26908 12311 26911
rect 12526 26908 12532 26920
rect 12299 26880 12532 26908
rect 12299 26877 12311 26880
rect 12253 26871 12311 26877
rect 12526 26868 12532 26880
rect 12584 26868 12590 26920
rect 13354 26908 13360 26920
rect 13315 26880 13360 26908
rect 13354 26868 13360 26880
rect 13412 26868 13418 26920
rect 3142 26800 3148 26852
rect 3200 26800 3206 26852
rect 4709 26843 4767 26849
rect 4709 26809 4721 26843
rect 4755 26840 4767 26843
rect 5718 26840 5724 26852
rect 4755 26812 5724 26840
rect 4755 26809 4767 26812
rect 4709 26803 4767 26809
rect 5718 26800 5724 26812
rect 5776 26800 5782 26852
rect 13924 26840 13952 26939
rect 14274 26936 14280 26948
rect 14332 26936 14338 26988
rect 16853 26979 16911 26985
rect 16853 26945 16865 26979
rect 16899 26976 16911 26979
rect 16942 26976 16948 26988
rect 16899 26948 16948 26976
rect 16899 26945 16911 26948
rect 16853 26939 16911 26945
rect 16942 26936 16948 26948
rect 17000 26936 17006 26988
rect 17052 26976 17080 27016
rect 17120 27013 17132 27047
rect 17166 27044 17178 27047
rect 18046 27044 18052 27056
rect 17166 27016 18052 27044
rect 17166 27013 17178 27016
rect 17120 27007 17178 27013
rect 18046 27004 18052 27016
rect 18104 27004 18110 27056
rect 26237 27047 26295 27053
rect 26237 27044 26249 27047
rect 19168 27016 22508 27044
rect 19168 26976 19196 27016
rect 19426 26976 19432 26988
rect 17052 26948 19196 26976
rect 19387 26948 19432 26976
rect 19426 26936 19432 26948
rect 19484 26936 19490 26988
rect 19536 26948 20208 26976
rect 13998 26868 14004 26920
rect 14056 26908 14062 26920
rect 14182 26908 14188 26920
rect 14056 26880 14101 26908
rect 14143 26880 14188 26908
rect 14056 26868 14062 26880
rect 14182 26868 14188 26880
rect 14240 26868 14246 26920
rect 19536 26908 19564 26948
rect 19168 26880 19564 26908
rect 19168 26840 19196 26880
rect 19610 26868 19616 26920
rect 19668 26908 19674 26920
rect 19705 26911 19763 26917
rect 19705 26908 19717 26911
rect 19668 26880 19717 26908
rect 19668 26868 19674 26880
rect 19705 26877 19717 26880
rect 19751 26877 19763 26911
rect 19705 26871 19763 26877
rect 13924 26812 16574 26840
rect 4433 26775 4491 26781
rect 4433 26741 4445 26775
rect 4479 26772 4491 26775
rect 4614 26772 4620 26784
rect 4479 26744 4620 26772
rect 4479 26741 4491 26744
rect 4433 26735 4491 26741
rect 4614 26732 4620 26744
rect 4672 26732 4678 26784
rect 10594 26732 10600 26784
rect 10652 26772 10658 26784
rect 12621 26775 12679 26781
rect 12621 26772 12633 26775
rect 10652 26744 12633 26772
rect 10652 26732 10658 26744
rect 12621 26741 12633 26744
rect 12667 26741 12679 26775
rect 12621 26735 12679 26741
rect 13998 26732 14004 26784
rect 14056 26772 14062 26784
rect 14918 26772 14924 26784
rect 14056 26744 14924 26772
rect 14056 26732 14062 26744
rect 14918 26732 14924 26744
rect 14976 26772 14982 26784
rect 16025 26775 16083 26781
rect 16025 26772 16037 26775
rect 14976 26744 16037 26772
rect 14976 26732 14982 26744
rect 16025 26741 16037 26744
rect 16071 26772 16083 26775
rect 16114 26772 16120 26784
rect 16071 26744 16120 26772
rect 16071 26741 16083 26744
rect 16025 26735 16083 26741
rect 16114 26732 16120 26744
rect 16172 26732 16178 26784
rect 16209 26775 16267 26781
rect 16209 26741 16221 26775
rect 16255 26772 16267 26775
rect 16298 26772 16304 26784
rect 16255 26744 16304 26772
rect 16255 26741 16267 26744
rect 16209 26735 16267 26741
rect 16298 26732 16304 26744
rect 16356 26732 16362 26784
rect 16546 26772 16574 26812
rect 17788 26812 19196 26840
rect 19245 26843 19303 26849
rect 17788 26772 17816 26812
rect 19245 26809 19257 26843
rect 19291 26840 19303 26843
rect 20070 26840 20076 26852
rect 19291 26812 20076 26840
rect 19291 26809 19303 26812
rect 19245 26803 19303 26809
rect 20070 26800 20076 26812
rect 20128 26800 20134 26852
rect 16546 26744 17816 26772
rect 18414 26732 18420 26784
rect 18472 26772 18478 26784
rect 19613 26775 19671 26781
rect 19613 26772 19625 26775
rect 18472 26744 19625 26772
rect 18472 26732 18478 26744
rect 19613 26741 19625 26744
rect 19659 26741 19671 26775
rect 20180 26772 20208 26948
rect 22094 26936 22100 26988
rect 22152 26976 22158 26988
rect 22189 26979 22247 26985
rect 22189 26976 22201 26979
rect 22152 26948 22201 26976
rect 22152 26936 22158 26948
rect 22189 26945 22201 26948
rect 22235 26945 22247 26979
rect 22189 26939 22247 26945
rect 22370 26936 22376 26988
rect 22428 26976 22434 26988
rect 22480 26985 22508 27016
rect 24596 27016 26249 27044
rect 22465 26979 22523 26985
rect 22465 26976 22477 26979
rect 22428 26948 22477 26976
rect 22428 26936 22434 26948
rect 22465 26945 22477 26948
rect 22511 26976 22523 26979
rect 24210 26976 24216 26988
rect 22511 26948 24216 26976
rect 22511 26945 22523 26948
rect 22465 26939 22523 26945
rect 24210 26936 24216 26948
rect 24268 26936 24274 26988
rect 24596 26985 24624 27016
rect 26237 27013 26249 27016
rect 26283 27013 26295 27047
rect 26237 27007 26295 27013
rect 31757 27047 31815 27053
rect 31757 27013 31769 27047
rect 31803 27044 31815 27047
rect 32490 27044 32496 27056
rect 31803 27016 32496 27044
rect 31803 27013 31815 27016
rect 31757 27007 31815 27013
rect 32490 27004 32496 27016
rect 32548 27044 32554 27056
rect 32548 27016 33180 27044
rect 32548 27004 32554 27016
rect 24581 26979 24639 26985
rect 24581 26945 24593 26979
rect 24627 26945 24639 26979
rect 24762 26976 24768 26988
rect 24723 26948 24768 26976
rect 24581 26939 24639 26945
rect 24762 26936 24768 26948
rect 24820 26936 24826 26988
rect 24854 26936 24860 26988
rect 24912 26976 24918 26988
rect 25130 26976 25136 26988
rect 24912 26948 25136 26976
rect 24912 26936 24918 26948
rect 25130 26936 25136 26948
rect 25188 26936 25194 26988
rect 26053 26979 26111 26985
rect 26053 26945 26065 26979
rect 26099 26976 26111 26979
rect 27614 26976 27620 26988
rect 26099 26948 27620 26976
rect 26099 26945 26111 26948
rect 26053 26939 26111 26945
rect 27614 26936 27620 26948
rect 27672 26936 27678 26988
rect 27890 26976 27896 26988
rect 27851 26948 27896 26976
rect 27890 26936 27896 26948
rect 27948 26936 27954 26988
rect 27982 26936 27988 26988
rect 28040 26976 28046 26988
rect 28166 26976 28172 26988
rect 28040 26948 28085 26976
rect 28127 26948 28172 26976
rect 28040 26936 28046 26948
rect 28166 26936 28172 26948
rect 28224 26936 28230 26988
rect 28261 26979 28319 26985
rect 28261 26945 28273 26979
rect 28307 26976 28319 26979
rect 28626 26976 28632 26988
rect 28307 26948 28632 26976
rect 28307 26945 28319 26948
rect 28261 26939 28319 26945
rect 28626 26936 28632 26948
rect 28684 26936 28690 26988
rect 31386 26976 31392 26988
rect 31347 26948 31392 26976
rect 31386 26936 31392 26948
rect 31444 26936 31450 26988
rect 31665 26979 31723 26985
rect 31665 26945 31677 26979
rect 31711 26976 31723 26979
rect 31846 26976 31852 26988
rect 31711 26948 31852 26976
rect 31711 26945 31723 26948
rect 31665 26939 31723 26945
rect 31846 26936 31852 26948
rect 31904 26936 31910 26988
rect 32582 26976 32588 26988
rect 32543 26948 32588 26976
rect 32582 26936 32588 26948
rect 32640 26936 32646 26988
rect 33152 26985 33180 27016
rect 33137 26979 33195 26985
rect 33137 26945 33149 26979
rect 33183 26945 33195 26979
rect 33137 26939 33195 26945
rect 23474 26868 23480 26920
rect 23532 26908 23538 26920
rect 25961 26911 26019 26917
rect 25961 26908 25973 26911
rect 23532 26880 25973 26908
rect 23532 26868 23538 26880
rect 25961 26877 25973 26880
rect 26007 26908 26019 26911
rect 32858 26908 32864 26920
rect 26007 26880 32864 26908
rect 26007 26877 26019 26880
rect 25961 26871 26019 26877
rect 32858 26868 32864 26880
rect 32916 26868 32922 26920
rect 33410 26908 33416 26920
rect 33371 26880 33416 26908
rect 33410 26868 33416 26880
rect 33468 26868 33474 26920
rect 24854 26800 24860 26852
rect 24912 26840 24918 26852
rect 25041 26843 25099 26849
rect 25041 26840 25053 26843
rect 24912 26812 25053 26840
rect 24912 26800 24918 26812
rect 25041 26809 25053 26812
rect 25087 26809 25099 26843
rect 25041 26803 25099 26809
rect 25130 26800 25136 26852
rect 25188 26840 25194 26852
rect 27430 26840 27436 26852
rect 25188 26812 27436 26840
rect 25188 26800 25194 26812
rect 27430 26800 27436 26812
rect 27488 26800 27494 26852
rect 27709 26775 27767 26781
rect 27709 26772 27721 26775
rect 20180 26744 27721 26772
rect 19613 26735 19671 26741
rect 27709 26741 27721 26744
rect 27755 26741 27767 26775
rect 27709 26735 27767 26741
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 8478 26528 8484 26580
rect 8536 26568 8542 26580
rect 9125 26571 9183 26577
rect 9125 26568 9137 26571
rect 8536 26540 9137 26568
rect 8536 26528 8542 26540
rect 9125 26537 9137 26540
rect 9171 26537 9183 26571
rect 12526 26568 12532 26580
rect 9125 26531 9183 26537
rect 12360 26540 12532 26568
rect 5077 26503 5135 26509
rect 2792 26472 4752 26500
rect 2792 26441 2820 26472
rect 2777 26435 2835 26441
rect 2777 26401 2789 26435
rect 2823 26401 2835 26435
rect 4614 26432 4620 26444
rect 4575 26404 4620 26432
rect 2777 26395 2835 26401
rect 4614 26392 4620 26404
rect 4672 26392 4678 26444
rect 4724 26432 4752 26472
rect 5077 26469 5089 26503
rect 5123 26500 5135 26503
rect 5810 26500 5816 26512
rect 5123 26472 5816 26500
rect 5123 26469 5135 26472
rect 5077 26463 5135 26469
rect 5810 26460 5816 26472
rect 5868 26460 5874 26512
rect 10045 26503 10103 26509
rect 10045 26469 10057 26503
rect 10091 26469 10103 26503
rect 10045 26463 10103 26469
rect 10060 26432 10088 26463
rect 12161 26435 12219 26441
rect 12161 26432 12173 26435
rect 4724 26404 5396 26432
rect 5368 26376 5396 26404
rect 9324 26404 10088 26432
rect 10336 26404 12173 26432
rect 2685 26367 2743 26373
rect 2685 26333 2697 26367
rect 2731 26364 2743 26367
rect 4157 26367 4215 26373
rect 2731 26336 4108 26364
rect 2731 26333 2743 26336
rect 2685 26327 2743 26333
rect 3142 26256 3148 26308
rect 3200 26296 3206 26308
rect 3329 26299 3387 26305
rect 3329 26296 3341 26299
rect 3200 26268 3341 26296
rect 3200 26256 3206 26268
rect 3329 26265 3341 26268
rect 3375 26265 3387 26299
rect 3329 26259 3387 26265
rect 3970 26228 3976 26240
rect 3931 26200 3976 26228
rect 3970 26188 3976 26200
rect 4028 26188 4034 26240
rect 4080 26228 4108 26336
rect 4157 26333 4169 26367
rect 4203 26333 4215 26367
rect 4157 26327 4215 26333
rect 4172 26296 4200 26327
rect 4246 26324 4252 26376
rect 4304 26364 4310 26376
rect 4525 26367 4583 26373
rect 4304 26336 4349 26364
rect 4304 26324 4310 26336
rect 4525 26333 4537 26367
rect 4571 26364 4583 26367
rect 4706 26364 4712 26376
rect 4571 26336 4712 26364
rect 4571 26333 4583 26336
rect 4525 26327 4583 26333
rect 4706 26324 4712 26336
rect 4764 26324 4770 26376
rect 4982 26324 4988 26376
rect 5040 26364 5046 26376
rect 5350 26364 5356 26376
rect 5040 26336 5212 26364
rect 5311 26336 5356 26364
rect 5040 26324 5046 26336
rect 4614 26296 4620 26308
rect 4172 26268 4620 26296
rect 4614 26256 4620 26268
rect 4672 26256 4678 26308
rect 5074 26296 5080 26308
rect 5035 26268 5080 26296
rect 5074 26256 5080 26268
rect 5132 26256 5138 26308
rect 5184 26296 5212 26336
rect 5350 26324 5356 26336
rect 5408 26324 5414 26376
rect 8938 26324 8944 26376
rect 8996 26364 9002 26376
rect 9324 26373 9352 26404
rect 9309 26367 9367 26373
rect 9309 26364 9321 26367
rect 8996 26336 9321 26364
rect 8996 26324 9002 26336
rect 9309 26333 9321 26336
rect 9355 26333 9367 26367
rect 9582 26364 9588 26376
rect 9543 26336 9588 26364
rect 9309 26327 9367 26333
rect 9582 26324 9588 26336
rect 9640 26324 9646 26376
rect 10134 26324 10140 26376
rect 10192 26364 10198 26376
rect 10336 26373 10364 26404
rect 12161 26401 12173 26404
rect 12207 26401 12219 26435
rect 12161 26395 12219 26401
rect 10321 26367 10379 26373
rect 10321 26364 10333 26367
rect 10192 26336 10333 26364
rect 10192 26324 10198 26336
rect 10321 26333 10333 26336
rect 10367 26333 10379 26367
rect 12066 26364 12072 26376
rect 12027 26336 12072 26364
rect 10321 26327 10379 26333
rect 12066 26324 12072 26336
rect 12124 26324 12130 26376
rect 12360 26373 12388 26540
rect 12526 26528 12532 26540
rect 12584 26568 12590 26580
rect 26053 26571 26111 26577
rect 26053 26568 26065 26571
rect 12584 26540 26065 26568
rect 12584 26528 12590 26540
rect 26053 26537 26065 26540
rect 26099 26537 26111 26571
rect 26053 26531 26111 26537
rect 33873 26571 33931 26577
rect 33873 26537 33885 26571
rect 33919 26568 33931 26571
rect 34330 26568 34336 26580
rect 33919 26540 34336 26568
rect 33919 26537 33931 26540
rect 33873 26531 33931 26537
rect 34330 26528 34336 26540
rect 34388 26528 34394 26580
rect 20254 26460 20260 26512
rect 20312 26500 20318 26512
rect 20349 26503 20407 26509
rect 20349 26500 20361 26503
rect 20312 26472 20361 26500
rect 20312 26460 20318 26472
rect 20349 26469 20361 26472
rect 20395 26500 20407 26503
rect 20530 26500 20536 26512
rect 20395 26472 20536 26500
rect 20395 26469 20407 26472
rect 20349 26463 20407 26469
rect 20530 26460 20536 26472
rect 20588 26460 20594 26512
rect 22189 26503 22247 26509
rect 22189 26469 22201 26503
rect 22235 26500 22247 26503
rect 22235 26472 24164 26500
rect 22235 26469 22247 26472
rect 22189 26463 22247 26469
rect 14918 26432 14924 26444
rect 14879 26404 14924 26432
rect 14918 26392 14924 26404
rect 14976 26392 14982 26444
rect 20622 26432 20628 26444
rect 20548 26404 20628 26432
rect 12345 26367 12403 26373
rect 12345 26333 12357 26367
rect 12391 26364 12403 26367
rect 12434 26364 12440 26376
rect 12391 26336 12440 26364
rect 12391 26333 12403 26336
rect 12345 26327 12403 26333
rect 12434 26324 12440 26336
rect 12492 26324 12498 26376
rect 12713 26367 12771 26373
rect 12713 26333 12725 26367
rect 12759 26364 12771 26367
rect 13814 26364 13820 26376
rect 12759 26336 13820 26364
rect 12759 26333 12771 26336
rect 12713 26327 12771 26333
rect 13814 26324 13820 26336
rect 13872 26324 13878 26376
rect 14366 26364 14372 26376
rect 14327 26336 14372 26364
rect 14366 26324 14372 26336
rect 14424 26324 14430 26376
rect 16298 26364 16304 26376
rect 16259 26336 16304 26364
rect 16298 26324 16304 26336
rect 16356 26324 16362 26376
rect 20346 26324 20352 26376
rect 20404 26364 20410 26376
rect 20548 26373 20576 26404
rect 20622 26392 20628 26404
rect 20680 26392 20686 26444
rect 21453 26435 21511 26441
rect 21453 26401 21465 26435
rect 21499 26432 21511 26435
rect 21499 26404 22692 26432
rect 21499 26401 21511 26404
rect 21453 26395 21511 26401
rect 20533 26367 20591 26373
rect 20533 26364 20545 26367
rect 20404 26336 20545 26364
rect 20404 26324 20410 26336
rect 20533 26333 20545 26336
rect 20579 26333 20591 26367
rect 21358 26364 21364 26376
rect 21319 26336 21364 26364
rect 20533 26327 20591 26333
rect 21358 26324 21364 26336
rect 21416 26324 21422 26376
rect 21542 26364 21548 26376
rect 21503 26336 21548 26364
rect 21542 26324 21548 26336
rect 21600 26324 21606 26376
rect 22370 26364 22376 26376
rect 22331 26336 22376 26364
rect 22370 26324 22376 26336
rect 22428 26324 22434 26376
rect 22462 26324 22468 26376
rect 22520 26364 22526 26376
rect 22664 26373 22692 26404
rect 23474 26392 23480 26444
rect 23532 26432 23538 26444
rect 23661 26435 23719 26441
rect 23661 26432 23673 26435
rect 23532 26404 23673 26432
rect 23532 26392 23538 26404
rect 23661 26401 23673 26404
rect 23707 26432 23719 26435
rect 23750 26432 23756 26444
rect 23707 26404 23756 26432
rect 23707 26401 23719 26404
rect 23661 26395 23719 26401
rect 23750 26392 23756 26404
rect 23808 26392 23814 26444
rect 22649 26367 22707 26373
rect 22520 26336 22565 26364
rect 22520 26324 22526 26336
rect 22649 26333 22661 26367
rect 22695 26333 22707 26367
rect 22649 26327 22707 26333
rect 22741 26367 22799 26373
rect 22741 26333 22753 26367
rect 22787 26364 22799 26367
rect 23385 26367 23443 26373
rect 22787 26336 22876 26364
rect 22787 26333 22799 26336
rect 22741 26327 22799 26333
rect 5261 26299 5319 26305
rect 5261 26296 5273 26299
rect 5184 26268 5273 26296
rect 5261 26265 5273 26268
rect 5307 26296 5319 26299
rect 6914 26296 6920 26308
rect 5307 26268 6920 26296
rect 5307 26265 5319 26268
rect 5261 26259 5319 26265
rect 6914 26256 6920 26268
rect 6972 26256 6978 26308
rect 9858 26256 9864 26308
rect 9916 26296 9922 26308
rect 10045 26299 10103 26305
rect 10045 26296 10057 26299
rect 9916 26268 10057 26296
rect 9916 26256 9922 26268
rect 10045 26265 10057 26268
rect 10091 26265 10103 26299
rect 10045 26259 10103 26265
rect 19978 26256 19984 26308
rect 20036 26296 20042 26308
rect 20036 26268 20300 26296
rect 20036 26256 20042 26268
rect 4982 26228 4988 26240
rect 4080 26200 4988 26228
rect 4982 26188 4988 26200
rect 5040 26188 5046 26240
rect 9490 26228 9496 26240
rect 9451 26200 9496 26228
rect 9490 26188 9496 26200
rect 9548 26188 9554 26240
rect 10226 26228 10232 26240
rect 10187 26200 10232 26228
rect 10226 26188 10232 26200
rect 10284 26188 10290 26240
rect 17586 26228 17592 26240
rect 17547 26200 17592 26228
rect 17586 26188 17592 26200
rect 17644 26188 17650 26240
rect 20272 26234 20300 26268
rect 20530 26234 20536 26246
rect 20272 26206 20536 26234
rect 20530 26194 20536 26206
rect 20588 26194 20594 26246
rect 22002 26188 22008 26240
rect 22060 26228 22066 26240
rect 22848 26234 22876 26336
rect 23385 26333 23397 26367
rect 23431 26364 23443 26367
rect 24026 26364 24032 26376
rect 23431 26336 24032 26364
rect 23431 26333 23443 26336
rect 23385 26327 23443 26333
rect 24026 26324 24032 26336
rect 24084 26324 24090 26376
rect 24136 26296 24164 26472
rect 24210 26460 24216 26512
rect 24268 26500 24274 26512
rect 27890 26500 27896 26512
rect 24268 26472 27896 26500
rect 24268 26460 24274 26472
rect 27890 26460 27896 26472
rect 27948 26460 27954 26512
rect 27982 26460 27988 26512
rect 28040 26500 28046 26512
rect 32582 26500 32588 26512
rect 28040 26472 32260 26500
rect 32543 26472 32588 26500
rect 28040 26460 28046 26472
rect 25240 26404 25912 26432
rect 24854 26364 24860 26376
rect 24815 26336 24860 26364
rect 24854 26324 24860 26336
rect 24912 26324 24918 26376
rect 25240 26373 25268 26404
rect 25225 26367 25283 26373
rect 25225 26333 25237 26367
rect 25271 26333 25283 26367
rect 25225 26327 25283 26333
rect 25317 26367 25375 26373
rect 25317 26333 25329 26367
rect 25363 26333 25375 26367
rect 25317 26327 25375 26333
rect 25332 26296 25360 26327
rect 24136 26268 25360 26296
rect 25884 26296 25912 26404
rect 28074 26392 28080 26444
rect 28132 26432 28138 26444
rect 32232 26432 32260 26472
rect 32582 26460 32588 26472
rect 32640 26460 32646 26512
rect 33410 26500 33416 26512
rect 32968 26472 33416 26500
rect 32968 26441 32996 26472
rect 33410 26460 33416 26472
rect 33468 26460 33474 26512
rect 32953 26435 33011 26441
rect 32953 26432 32965 26435
rect 28132 26404 31800 26432
rect 32232 26404 32965 26432
rect 28132 26392 28138 26404
rect 26053 26367 26111 26373
rect 26053 26333 26065 26367
rect 26099 26364 26111 26367
rect 26234 26364 26240 26376
rect 26099 26336 26240 26364
rect 26099 26333 26111 26336
rect 26053 26327 26111 26333
rect 26234 26324 26240 26336
rect 26292 26364 26298 26376
rect 26602 26364 26608 26376
rect 26292 26336 26608 26364
rect 26292 26324 26298 26336
rect 26602 26324 26608 26336
rect 26660 26324 26666 26376
rect 31772 26373 31800 26404
rect 32953 26401 32965 26404
rect 32999 26401 33011 26435
rect 32953 26395 33011 26401
rect 33042 26392 33048 26444
rect 33100 26432 33106 26444
rect 33100 26404 33732 26432
rect 33100 26392 33106 26404
rect 31481 26367 31539 26373
rect 31481 26333 31493 26367
rect 31527 26364 31539 26367
rect 31757 26367 31815 26373
rect 31527 26336 31616 26364
rect 31527 26333 31539 26336
rect 31481 26327 31539 26333
rect 27522 26296 27528 26308
rect 25884 26268 27528 26296
rect 27522 26256 27528 26268
rect 27580 26256 27586 26308
rect 22756 26228 22876 26234
rect 31294 26228 31300 26240
rect 22060 26206 22876 26228
rect 22060 26200 22784 26206
rect 31255 26200 31300 26228
rect 22060 26188 22066 26200
rect 31294 26188 31300 26200
rect 31352 26188 31358 26240
rect 31588 26228 31616 26336
rect 31757 26333 31769 26367
rect 31803 26333 31815 26367
rect 32858 26364 32864 26376
rect 32819 26336 32864 26364
rect 31757 26327 31815 26333
rect 32858 26324 32864 26336
rect 32916 26324 32922 26376
rect 33704 26373 33732 26404
rect 33505 26367 33563 26373
rect 33505 26333 33517 26367
rect 33551 26333 33563 26367
rect 33505 26327 33563 26333
rect 33689 26367 33747 26373
rect 33689 26333 33701 26367
rect 33735 26333 33747 26367
rect 33689 26327 33747 26333
rect 31665 26299 31723 26305
rect 31665 26265 31677 26299
rect 31711 26296 31723 26299
rect 31846 26296 31852 26308
rect 31711 26268 31852 26296
rect 31711 26265 31723 26268
rect 31665 26259 31723 26265
rect 31846 26256 31852 26268
rect 31904 26296 31910 26308
rect 32309 26299 32367 26305
rect 32309 26296 32321 26299
rect 31904 26268 32321 26296
rect 31904 26256 31910 26268
rect 32309 26265 32321 26268
rect 32355 26265 32367 26299
rect 32309 26259 32367 26265
rect 32674 26256 32680 26308
rect 32732 26296 32738 26308
rect 33520 26296 33548 26327
rect 32732 26268 33548 26296
rect 32732 26256 32738 26268
rect 32582 26228 32588 26240
rect 31588 26200 32588 26228
rect 32582 26188 32588 26200
rect 32640 26188 32646 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 4246 25984 4252 26036
rect 4304 26024 4310 26036
rect 5169 26027 5227 26033
rect 5169 26024 5181 26027
rect 4304 25996 5181 26024
rect 4304 25984 4310 25996
rect 5169 25993 5181 25996
rect 5215 25993 5227 26027
rect 10778 26024 10784 26036
rect 5169 25987 5227 25993
rect 5552 25996 10784 26024
rect 3142 25956 3148 25968
rect 2424 25928 3148 25956
rect 2424 25897 2452 25928
rect 3142 25916 3148 25928
rect 3200 25916 3206 25968
rect 4709 25959 4767 25965
rect 4709 25925 4721 25959
rect 4755 25956 4767 25959
rect 5258 25956 5264 25968
rect 4755 25928 5264 25956
rect 4755 25925 4767 25928
rect 4709 25919 4767 25925
rect 5258 25916 5264 25928
rect 5316 25956 5322 25968
rect 5552 25965 5580 25996
rect 10778 25984 10784 25996
rect 10836 25984 10842 26036
rect 12434 26024 12440 26036
rect 12395 25996 12440 26024
rect 12434 25984 12440 25996
rect 12492 25984 12498 26036
rect 18417 26027 18475 26033
rect 18417 25993 18429 26027
rect 18463 26024 18475 26027
rect 19334 26024 19340 26036
rect 18463 25996 19340 26024
rect 18463 25993 18475 25996
rect 18417 25987 18475 25993
rect 19334 25984 19340 25996
rect 19392 26024 19398 26036
rect 20346 26024 20352 26036
rect 19392 25996 20352 26024
rect 19392 25984 19398 25996
rect 20346 25984 20352 25996
rect 20404 25984 20410 26036
rect 5445 25959 5503 25965
rect 5445 25956 5457 25959
rect 5316 25928 5457 25956
rect 5316 25916 5322 25928
rect 5445 25925 5457 25928
rect 5491 25925 5503 25959
rect 5445 25919 5503 25925
rect 5537 25959 5595 25965
rect 5537 25925 5549 25959
rect 5583 25925 5595 25959
rect 8938 25956 8944 25968
rect 8899 25928 8944 25956
rect 5537 25919 5595 25925
rect 8938 25916 8944 25928
rect 8996 25916 9002 25968
rect 9876 25928 10640 25956
rect 9876 25900 9904 25928
rect 2409 25891 2467 25897
rect 2409 25857 2421 25891
rect 2455 25857 2467 25891
rect 2409 25851 2467 25857
rect 2593 25891 2651 25897
rect 2593 25857 2605 25891
rect 2639 25888 2651 25891
rect 3329 25891 3387 25897
rect 2639 25860 3280 25888
rect 2639 25857 2651 25860
rect 2593 25851 2651 25857
rect 3050 25820 3056 25832
rect 3011 25792 3056 25820
rect 3050 25780 3056 25792
rect 3108 25780 3114 25832
rect 3252 25820 3280 25860
rect 3329 25857 3341 25891
rect 3375 25888 3387 25891
rect 3970 25888 3976 25900
rect 3375 25860 3976 25888
rect 3375 25857 3387 25860
rect 3329 25851 3387 25857
rect 3970 25848 3976 25860
rect 4028 25848 4034 25900
rect 5350 25888 5356 25900
rect 5311 25860 5356 25888
rect 5350 25848 5356 25860
rect 5408 25848 5414 25900
rect 5718 25888 5724 25900
rect 5679 25860 5724 25888
rect 5718 25848 5724 25860
rect 5776 25848 5782 25900
rect 5810 25848 5816 25900
rect 5868 25888 5874 25900
rect 5868 25860 5913 25888
rect 5868 25848 5874 25860
rect 7098 25848 7104 25900
rect 7156 25888 7162 25900
rect 7558 25888 7564 25900
rect 7156 25860 7564 25888
rect 7156 25848 7162 25860
rect 7558 25848 7564 25860
rect 7616 25888 7622 25900
rect 9858 25888 9864 25900
rect 7616 25860 9720 25888
rect 9819 25860 9864 25888
rect 7616 25848 7622 25860
rect 5074 25820 5080 25832
rect 3252 25792 5080 25820
rect 5074 25780 5080 25792
rect 5132 25780 5138 25832
rect 5736 25820 5764 25848
rect 8570 25820 8576 25832
rect 5736 25792 8576 25820
rect 8570 25780 8576 25792
rect 8628 25780 8634 25832
rect 9692 25820 9720 25860
rect 9858 25848 9864 25860
rect 9916 25848 9922 25900
rect 10042 25888 10048 25900
rect 10003 25860 10048 25888
rect 10042 25848 10048 25860
rect 10100 25848 10106 25900
rect 10612 25897 10640 25928
rect 16022 25916 16028 25968
rect 16080 25956 16086 25968
rect 16209 25959 16267 25965
rect 16209 25956 16221 25959
rect 16080 25928 16221 25956
rect 16080 25916 16086 25928
rect 16209 25925 16221 25928
rect 16255 25956 16267 25959
rect 17126 25956 17132 25968
rect 16255 25928 17132 25956
rect 16255 25925 16267 25928
rect 16209 25919 16267 25925
rect 17126 25916 17132 25928
rect 17184 25916 17190 25968
rect 10137 25891 10195 25897
rect 10137 25857 10149 25891
rect 10183 25857 10195 25891
rect 10137 25851 10195 25857
rect 10597 25891 10655 25897
rect 10597 25857 10609 25891
rect 10643 25857 10655 25891
rect 10597 25851 10655 25857
rect 10781 25891 10839 25897
rect 10781 25857 10793 25891
rect 10827 25888 10839 25891
rect 12069 25891 12127 25897
rect 12069 25888 12081 25891
rect 10827 25860 12081 25888
rect 10827 25857 10839 25860
rect 10781 25851 10839 25857
rect 12069 25857 12081 25860
rect 12115 25857 12127 25891
rect 12253 25891 12311 25897
rect 12253 25888 12265 25891
rect 12069 25851 12127 25857
rect 12176 25860 12265 25888
rect 10152 25820 10180 25851
rect 10226 25820 10232 25832
rect 9692 25792 10088 25820
rect 10139 25792 10232 25820
rect 9309 25755 9367 25761
rect 9309 25721 9321 25755
rect 9355 25752 9367 25755
rect 9490 25752 9496 25764
rect 9355 25724 9496 25752
rect 9355 25721 9367 25724
rect 9309 25715 9367 25721
rect 9490 25712 9496 25724
rect 9548 25752 9554 25764
rect 9953 25755 10011 25761
rect 9953 25752 9965 25755
rect 9548 25724 9965 25752
rect 9548 25712 9554 25724
rect 9953 25721 9965 25724
rect 9999 25721 10011 25755
rect 10060 25752 10088 25792
rect 10226 25780 10232 25792
rect 10284 25820 10290 25832
rect 10796 25820 10824 25851
rect 10284 25792 10824 25820
rect 10284 25780 10290 25792
rect 12176 25752 12204 25860
rect 12253 25857 12265 25860
rect 12299 25857 12311 25891
rect 12253 25851 12311 25857
rect 12529 25891 12587 25897
rect 12529 25857 12541 25891
rect 12575 25888 12587 25891
rect 13814 25888 13820 25900
rect 12575 25860 13820 25888
rect 12575 25857 12587 25860
rect 12529 25851 12587 25857
rect 13814 25848 13820 25860
rect 13872 25848 13878 25900
rect 15654 25888 15660 25900
rect 15615 25860 15660 25888
rect 15654 25848 15660 25860
rect 15712 25848 15718 25900
rect 17304 25891 17362 25897
rect 17304 25857 17316 25891
rect 17350 25888 17362 25891
rect 17862 25888 17868 25900
rect 17350 25860 17868 25888
rect 17350 25857 17362 25860
rect 17304 25851 17362 25857
rect 17862 25848 17868 25860
rect 17920 25848 17926 25900
rect 23845 25891 23903 25897
rect 23845 25857 23857 25891
rect 23891 25888 23903 25891
rect 24854 25888 24860 25900
rect 23891 25860 24860 25888
rect 23891 25857 23903 25860
rect 23845 25851 23903 25857
rect 24854 25848 24860 25860
rect 24912 25848 24918 25900
rect 28629 25891 28687 25897
rect 28629 25857 28641 25891
rect 28675 25888 28687 25891
rect 30926 25888 30932 25900
rect 28675 25860 30932 25888
rect 28675 25857 28687 25860
rect 28629 25851 28687 25857
rect 30926 25848 30932 25860
rect 30984 25848 30990 25900
rect 31018 25848 31024 25900
rect 31076 25888 31082 25900
rect 31202 25888 31208 25900
rect 31076 25860 31121 25888
rect 31163 25860 31208 25888
rect 31076 25848 31082 25860
rect 31202 25848 31208 25860
rect 31260 25848 31266 25900
rect 31297 25891 31355 25897
rect 31297 25857 31309 25891
rect 31343 25888 31355 25891
rect 32306 25888 32312 25900
rect 31343 25860 32312 25888
rect 31343 25857 31355 25860
rect 31297 25851 31355 25857
rect 32306 25848 32312 25860
rect 32364 25848 32370 25900
rect 16942 25780 16948 25832
rect 17000 25820 17006 25832
rect 17037 25823 17095 25829
rect 17037 25820 17049 25823
rect 17000 25792 17049 25820
rect 17000 25780 17006 25792
rect 17037 25789 17049 25792
rect 17083 25789 17095 25823
rect 17037 25783 17095 25789
rect 21266 25780 21272 25832
rect 21324 25820 21330 25832
rect 23566 25820 23572 25832
rect 21324 25792 23572 25820
rect 21324 25780 21330 25792
rect 23566 25780 23572 25792
rect 23624 25820 23630 25832
rect 24029 25823 24087 25829
rect 24029 25820 24041 25823
rect 23624 25792 24041 25820
rect 23624 25780 23630 25792
rect 24029 25789 24041 25792
rect 24075 25789 24087 25823
rect 24029 25783 24087 25789
rect 10060 25724 12204 25752
rect 9953 25715 10011 25721
rect 2501 25687 2559 25693
rect 2501 25653 2513 25687
rect 2547 25684 2559 25687
rect 4062 25684 4068 25696
rect 2547 25656 4068 25684
rect 2547 25653 2559 25656
rect 2501 25647 2559 25653
rect 4062 25644 4068 25656
rect 4120 25644 4126 25696
rect 8294 25644 8300 25696
rect 8352 25684 8358 25696
rect 9401 25687 9459 25693
rect 9401 25684 9413 25687
rect 8352 25656 9413 25684
rect 8352 25644 8358 25656
rect 9401 25653 9413 25656
rect 9447 25653 9459 25687
rect 9401 25647 9459 25653
rect 9674 25644 9680 25696
rect 9732 25684 9738 25696
rect 10689 25687 10747 25693
rect 10689 25684 10701 25687
rect 9732 25656 10701 25684
rect 9732 25644 9738 25656
rect 10689 25653 10701 25656
rect 10735 25653 10747 25687
rect 10689 25647 10747 25653
rect 20254 25644 20260 25696
rect 20312 25684 20318 25696
rect 21284 25684 21312 25780
rect 29914 25684 29920 25696
rect 20312 25656 21312 25684
rect 29875 25656 29920 25684
rect 20312 25644 20318 25656
rect 29914 25644 29920 25656
rect 29972 25644 29978 25696
rect 30834 25684 30840 25696
rect 30795 25656 30840 25684
rect 30834 25644 30840 25656
rect 30892 25644 30898 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 3237 25483 3295 25489
rect 3237 25449 3249 25483
rect 3283 25480 3295 25483
rect 4614 25480 4620 25492
rect 3283 25452 4620 25480
rect 3283 25449 3295 25452
rect 3237 25443 3295 25449
rect 4614 25440 4620 25452
rect 4672 25440 4678 25492
rect 5074 25440 5080 25492
rect 5132 25480 5138 25492
rect 5353 25483 5411 25489
rect 5353 25480 5365 25483
rect 5132 25452 5365 25480
rect 5132 25440 5138 25452
rect 5353 25449 5365 25452
rect 5399 25449 5411 25483
rect 5353 25443 5411 25449
rect 7834 25440 7840 25492
rect 7892 25480 7898 25492
rect 8389 25483 8447 25489
rect 8389 25480 8401 25483
rect 7892 25452 8401 25480
rect 7892 25440 7898 25452
rect 8389 25449 8401 25452
rect 8435 25480 8447 25483
rect 9582 25480 9588 25492
rect 8435 25452 9588 25480
rect 8435 25449 8447 25452
rect 8389 25443 8447 25449
rect 9582 25440 9588 25452
rect 9640 25440 9646 25492
rect 10502 25440 10508 25492
rect 10560 25480 10566 25492
rect 10689 25483 10747 25489
rect 10689 25480 10701 25483
rect 10560 25452 10701 25480
rect 10560 25440 10566 25452
rect 10689 25449 10701 25452
rect 10735 25480 10747 25483
rect 16482 25480 16488 25492
rect 10735 25452 12388 25480
rect 10735 25449 10747 25452
rect 10689 25443 10747 25449
rect 3510 25372 3516 25424
rect 3568 25412 3574 25424
rect 3973 25415 4031 25421
rect 3973 25412 3985 25415
rect 3568 25384 3985 25412
rect 3568 25372 3574 25384
rect 3973 25381 3985 25384
rect 4019 25381 4031 25415
rect 3973 25375 4031 25381
rect 4154 25372 4160 25424
rect 4212 25412 4218 25424
rect 4982 25412 4988 25424
rect 4212 25384 4988 25412
rect 4212 25372 4218 25384
rect 4982 25372 4988 25384
rect 5040 25372 5046 25424
rect 7561 25415 7619 25421
rect 7561 25381 7573 25415
rect 7607 25412 7619 25415
rect 10873 25415 10931 25421
rect 7607 25384 9352 25412
rect 7607 25381 7619 25384
rect 7561 25375 7619 25381
rect 5350 25344 5356 25356
rect 3252 25316 5356 25344
rect 3252 25285 3280 25316
rect 5350 25304 5356 25316
rect 5408 25304 5414 25356
rect 8570 25344 8576 25356
rect 7760 25316 8340 25344
rect 8531 25316 8576 25344
rect 3237 25279 3295 25285
rect 3237 25245 3249 25279
rect 3283 25245 3295 25279
rect 3237 25239 3295 25245
rect 3421 25279 3479 25285
rect 3421 25245 3433 25279
rect 3467 25245 3479 25279
rect 3421 25239 3479 25245
rect 3436 25140 3464 25239
rect 4062 25236 4068 25288
rect 4120 25276 4126 25288
rect 4157 25279 4215 25285
rect 4157 25276 4169 25279
rect 4120 25248 4169 25276
rect 4120 25236 4126 25248
rect 4157 25245 4169 25248
rect 4203 25245 4215 25279
rect 4157 25239 4215 25245
rect 4249 25279 4307 25285
rect 4249 25245 4261 25279
rect 4295 25276 4307 25279
rect 4706 25276 4712 25288
rect 4295 25248 4712 25276
rect 4295 25245 4307 25248
rect 4249 25239 4307 25245
rect 4706 25236 4712 25248
rect 4764 25236 4770 25288
rect 5077 25279 5135 25285
rect 5077 25245 5089 25279
rect 5123 25245 5135 25279
rect 5077 25239 5135 25245
rect 3973 25211 4031 25217
rect 3973 25177 3985 25211
rect 4019 25208 4031 25211
rect 4614 25208 4620 25220
rect 4019 25180 4620 25208
rect 4019 25177 4031 25180
rect 3973 25171 4031 25177
rect 4614 25168 4620 25180
rect 4672 25168 4678 25220
rect 5092 25208 5120 25239
rect 5166 25236 5172 25288
rect 5224 25276 5230 25288
rect 7760 25285 7788 25316
rect 8312 25288 8340 25316
rect 8570 25304 8576 25316
rect 8628 25304 8634 25356
rect 9324 25353 9352 25384
rect 10873 25381 10885 25415
rect 10919 25381 10931 25415
rect 10873 25375 10931 25381
rect 9309 25347 9367 25353
rect 9309 25313 9321 25347
rect 9355 25313 9367 25347
rect 9674 25344 9680 25356
rect 9635 25316 9680 25344
rect 9309 25307 9367 25313
rect 9674 25304 9680 25316
rect 9732 25304 9738 25356
rect 9769 25347 9827 25353
rect 9769 25313 9781 25347
rect 9815 25344 9827 25347
rect 10888 25344 10916 25375
rect 9815 25316 10916 25344
rect 9815 25313 9827 25316
rect 9769 25307 9827 25313
rect 7745 25279 7803 25285
rect 5224 25248 5269 25276
rect 5224 25236 5230 25248
rect 7745 25245 7757 25279
rect 7791 25245 7803 25279
rect 7745 25239 7803 25245
rect 7834 25236 7840 25288
rect 7892 25276 7898 25288
rect 8294 25276 8300 25288
rect 7892 25248 7937 25276
rect 8255 25248 8300 25276
rect 7892 25236 7898 25248
rect 8294 25236 8300 25248
rect 8352 25236 8358 25288
rect 9401 25279 9459 25285
rect 9401 25245 9413 25279
rect 9447 25276 9459 25279
rect 10042 25276 10048 25288
rect 9447 25248 10048 25276
rect 9447 25245 9459 25248
rect 9401 25239 9459 25245
rect 10042 25236 10048 25248
rect 10100 25236 10106 25288
rect 10321 25279 10379 25285
rect 10321 25245 10333 25279
rect 10367 25245 10379 25279
rect 10594 25276 10600 25288
rect 10555 25248 10600 25276
rect 10321 25239 10379 25245
rect 5258 25208 5264 25220
rect 5092 25180 5264 25208
rect 5258 25168 5264 25180
rect 5316 25168 5322 25220
rect 7561 25211 7619 25217
rect 7561 25177 7573 25211
rect 7607 25208 7619 25211
rect 8573 25211 8631 25217
rect 8573 25208 8585 25211
rect 7607 25180 8585 25208
rect 7607 25177 7619 25180
rect 7561 25171 7619 25177
rect 8573 25177 8585 25180
rect 8619 25177 8631 25211
rect 8573 25171 8631 25177
rect 8680 25180 9536 25208
rect 4154 25140 4160 25152
rect 3436 25112 4160 25140
rect 4154 25100 4160 25112
rect 4212 25100 4218 25152
rect 4632 25140 4660 25168
rect 7742 25140 7748 25152
rect 4632 25112 7748 25140
rect 7742 25100 7748 25112
rect 7800 25140 7806 25152
rect 8680 25140 8708 25180
rect 9122 25140 9128 25152
rect 7800 25112 8708 25140
rect 9083 25112 9128 25140
rect 7800 25100 7806 25112
rect 9122 25100 9128 25112
rect 9180 25100 9186 25152
rect 9508 25149 9536 25180
rect 9674 25168 9680 25220
rect 9732 25208 9738 25220
rect 10336 25208 10364 25239
rect 10594 25236 10600 25248
rect 10652 25236 10658 25288
rect 10686 25236 10692 25288
rect 10744 25276 10750 25288
rect 12360 25285 12388 25452
rect 12544 25452 16488 25480
rect 12544 25285 12572 25452
rect 16482 25440 16488 25452
rect 16540 25440 16546 25492
rect 16942 25480 16948 25492
rect 16903 25452 16948 25480
rect 16942 25440 16948 25452
rect 17000 25440 17006 25492
rect 17862 25480 17868 25492
rect 17823 25452 17868 25480
rect 17862 25440 17868 25452
rect 17920 25440 17926 25492
rect 20180 25452 20484 25480
rect 13449 25415 13507 25421
rect 13449 25381 13461 25415
rect 13495 25412 13507 25415
rect 14458 25412 14464 25424
rect 13495 25384 14464 25412
rect 13495 25381 13507 25384
rect 13449 25375 13507 25381
rect 14458 25372 14464 25384
rect 14516 25412 14522 25424
rect 20180 25412 20208 25452
rect 14516 25384 20208 25412
rect 20456 25412 20484 25452
rect 26206 25452 31616 25480
rect 26206 25412 26234 25452
rect 20456 25384 26234 25412
rect 14516 25372 14522 25384
rect 14642 25304 14648 25356
rect 14700 25344 14706 25356
rect 16758 25344 16764 25356
rect 14700 25316 16764 25344
rect 14700 25304 14706 25316
rect 16758 25304 16764 25316
rect 16816 25304 16822 25356
rect 20162 25344 20168 25356
rect 17972 25316 18368 25344
rect 11701 25279 11759 25285
rect 11701 25276 11713 25279
rect 10744 25248 11713 25276
rect 10744 25236 10750 25248
rect 11701 25245 11713 25248
rect 11747 25245 11759 25279
rect 11701 25239 11759 25245
rect 12345 25279 12403 25285
rect 12345 25245 12357 25279
rect 12391 25245 12403 25279
rect 12345 25239 12403 25245
rect 12529 25279 12587 25285
rect 12529 25245 12541 25279
rect 12575 25245 12587 25279
rect 12529 25239 12587 25245
rect 12618 25236 12624 25288
rect 12676 25276 12682 25288
rect 13173 25279 13231 25285
rect 13173 25276 13185 25279
rect 12676 25248 13185 25276
rect 12676 25236 12682 25248
rect 13173 25245 13185 25248
rect 13219 25245 13231 25279
rect 13446 25276 13452 25288
rect 13359 25248 13452 25276
rect 13173 25239 13231 25245
rect 13446 25236 13452 25248
rect 13504 25276 13510 25288
rect 17972 25276 18000 25316
rect 13504 25248 18000 25276
rect 13504 25236 13510 25248
rect 18046 25236 18052 25288
rect 18104 25276 18110 25288
rect 18340 25285 18368 25316
rect 19444 25316 20168 25344
rect 18325 25279 18383 25285
rect 18104 25248 18149 25276
rect 18104 25236 18110 25248
rect 18325 25245 18337 25279
rect 18371 25276 18383 25279
rect 18506 25276 18512 25288
rect 18371 25248 18512 25276
rect 18371 25245 18383 25248
rect 18325 25239 18383 25245
rect 18506 25236 18512 25248
rect 18564 25276 18570 25288
rect 19242 25276 19248 25288
rect 18564 25248 19248 25276
rect 18564 25236 18570 25248
rect 19242 25236 19248 25248
rect 19300 25236 19306 25288
rect 19444 25285 19472 25316
rect 20162 25304 20168 25316
rect 20220 25304 20226 25356
rect 20441 25347 20499 25353
rect 20441 25313 20453 25347
rect 20487 25344 20499 25347
rect 20622 25344 20628 25356
rect 20487 25316 20628 25344
rect 20487 25313 20499 25316
rect 20441 25307 20499 25313
rect 20622 25304 20628 25316
rect 20680 25304 20686 25356
rect 23750 25304 23756 25356
rect 23808 25304 23814 25356
rect 19429 25279 19487 25285
rect 19429 25245 19441 25279
rect 19475 25245 19487 25279
rect 19429 25239 19487 25245
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25245 19671 25279
rect 19613 25239 19671 25245
rect 20073 25279 20131 25285
rect 20073 25245 20085 25279
rect 20119 25276 20131 25279
rect 20254 25276 20260 25288
rect 20119 25248 20260 25276
rect 20119 25245 20131 25248
rect 20073 25239 20131 25245
rect 10778 25208 10784 25220
rect 9732 25180 10784 25208
rect 9732 25168 9738 25180
rect 10778 25168 10784 25180
rect 10836 25168 10842 25220
rect 11793 25211 11851 25217
rect 11793 25177 11805 25211
rect 11839 25208 11851 25211
rect 12894 25208 12900 25220
rect 11839 25180 12900 25208
rect 11839 25177 11851 25180
rect 11793 25171 11851 25177
rect 12894 25168 12900 25180
rect 12952 25168 12958 25220
rect 15657 25211 15715 25217
rect 15657 25177 15669 25211
rect 15703 25208 15715 25211
rect 16574 25208 16580 25220
rect 15703 25180 16580 25208
rect 15703 25177 15715 25180
rect 15657 25171 15715 25177
rect 16574 25168 16580 25180
rect 16632 25208 16638 25220
rect 17586 25208 17592 25220
rect 16632 25180 17592 25208
rect 16632 25168 16638 25180
rect 17586 25168 17592 25180
rect 17644 25168 17650 25220
rect 18233 25211 18291 25217
rect 18233 25177 18245 25211
rect 18279 25208 18291 25211
rect 19334 25208 19340 25220
rect 18279 25180 19340 25208
rect 18279 25177 18291 25180
rect 18233 25171 18291 25177
rect 19334 25168 19340 25180
rect 19392 25168 19398 25220
rect 19628 25208 19656 25239
rect 20254 25236 20260 25248
rect 20312 25236 20318 25288
rect 20349 25279 20407 25285
rect 20349 25245 20361 25279
rect 20395 25276 20407 25279
rect 22278 25276 22284 25288
rect 20395 25248 22284 25276
rect 20395 25245 20407 25248
rect 20349 25239 20407 25245
rect 22278 25236 22284 25248
rect 22336 25236 22342 25288
rect 23201 25279 23259 25285
rect 23201 25245 23213 25279
rect 23247 25276 23259 25279
rect 23768 25276 23796 25304
rect 23247 25248 23796 25276
rect 27341 25279 27399 25285
rect 23247 25245 23259 25248
rect 23201 25239 23259 25245
rect 27341 25245 27353 25279
rect 27387 25276 27399 25279
rect 29914 25276 29920 25288
rect 27387 25248 29920 25276
rect 27387 25245 27399 25248
rect 27341 25239 27399 25245
rect 29914 25236 29920 25248
rect 29972 25276 29978 25288
rect 30561 25279 30619 25285
rect 30561 25276 30573 25279
rect 29972 25248 30573 25276
rect 29972 25236 29978 25248
rect 30561 25245 30573 25248
rect 30607 25245 30619 25279
rect 30561 25239 30619 25245
rect 30828 25279 30886 25285
rect 30828 25245 30840 25279
rect 30874 25276 30886 25279
rect 31294 25276 31300 25288
rect 30874 25248 31300 25276
rect 30874 25245 30886 25248
rect 30828 25239 30886 25245
rect 31294 25236 31300 25248
rect 31352 25236 31358 25288
rect 31588 25276 31616 25452
rect 31846 25440 31852 25492
rect 31904 25480 31910 25492
rect 31941 25483 31999 25489
rect 31941 25480 31953 25483
rect 31904 25452 31953 25480
rect 31904 25440 31910 25452
rect 31941 25449 31953 25452
rect 31987 25449 31999 25483
rect 31941 25443 31999 25449
rect 32493 25279 32551 25285
rect 32493 25276 32505 25279
rect 31588 25248 32505 25276
rect 32493 25245 32505 25248
rect 32539 25245 32551 25279
rect 32493 25239 32551 25245
rect 23474 25208 23480 25220
rect 19628 25180 23480 25208
rect 23474 25168 23480 25180
rect 23532 25208 23538 25220
rect 23569 25211 23627 25217
rect 23569 25208 23581 25211
rect 23532 25180 23581 25208
rect 23532 25168 23538 25180
rect 23569 25177 23581 25180
rect 23615 25208 23627 25211
rect 23658 25208 23664 25220
rect 23615 25180 23664 25208
rect 23615 25177 23627 25180
rect 23569 25171 23627 25177
rect 23658 25168 23664 25180
rect 23716 25168 23722 25220
rect 27614 25217 27620 25220
rect 27608 25171 27620 25217
rect 27672 25208 27678 25220
rect 27672 25180 27708 25208
rect 27614 25168 27620 25171
rect 27672 25168 27678 25180
rect 9493 25143 9551 25149
rect 9493 25109 9505 25143
rect 9539 25109 9551 25143
rect 9493 25103 9551 25109
rect 12621 25143 12679 25149
rect 12621 25109 12633 25143
rect 12667 25140 12679 25143
rect 14642 25140 14648 25152
rect 12667 25112 14648 25140
rect 12667 25109 12679 25112
rect 12621 25103 12679 25109
rect 14642 25100 14648 25112
rect 14700 25100 14706 25152
rect 19613 25143 19671 25149
rect 19613 25109 19625 25143
rect 19659 25140 19671 25143
rect 20070 25140 20076 25152
rect 19659 25112 20076 25140
rect 19659 25109 19671 25112
rect 19613 25103 19671 25109
rect 20070 25100 20076 25112
rect 20128 25100 20134 25152
rect 28718 25140 28724 25152
rect 28679 25112 28724 25140
rect 28718 25100 28724 25112
rect 28776 25100 28782 25152
rect 32582 25140 32588 25152
rect 32543 25112 32588 25140
rect 32582 25100 32588 25112
rect 32640 25100 32646 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 9858 24936 9864 24948
rect 9819 24908 9864 24936
rect 9858 24896 9864 24908
rect 9916 24896 9922 24948
rect 10502 24936 10508 24948
rect 10463 24908 10508 24936
rect 10502 24896 10508 24908
rect 10560 24896 10566 24948
rect 17126 24896 17132 24948
rect 17184 24936 17190 24948
rect 24765 24939 24823 24945
rect 17184 24908 24716 24936
rect 17184 24896 17190 24908
rect 3050 24828 3056 24880
rect 3108 24868 3114 24880
rect 13265 24871 13323 24877
rect 3108 24840 4200 24868
rect 3108 24828 3114 24840
rect 4172 24800 4200 24840
rect 13265 24837 13277 24871
rect 13311 24868 13323 24871
rect 15654 24868 15660 24880
rect 13311 24840 15660 24868
rect 13311 24837 13323 24840
rect 13265 24831 13323 24837
rect 15654 24828 15660 24840
rect 15712 24828 15718 24880
rect 16482 24828 16488 24880
rect 16540 24868 16546 24880
rect 16540 24840 16620 24868
rect 16540 24828 16546 24840
rect 4706 24800 4712 24812
rect 4172 24772 4712 24800
rect 4706 24760 4712 24772
rect 4764 24800 4770 24812
rect 7837 24803 7895 24809
rect 7837 24800 7849 24803
rect 4764 24772 7849 24800
rect 4764 24760 4770 24772
rect 7837 24769 7849 24772
rect 7883 24800 7895 24803
rect 7926 24800 7932 24812
rect 7883 24772 7932 24800
rect 7883 24769 7895 24772
rect 7837 24763 7895 24769
rect 7926 24760 7932 24772
rect 7984 24760 7990 24812
rect 8104 24803 8162 24809
rect 8104 24769 8116 24803
rect 8150 24800 8162 24803
rect 9122 24800 9128 24812
rect 8150 24772 9128 24800
rect 8150 24769 8162 24772
rect 8104 24763 8162 24769
rect 9122 24760 9128 24772
rect 9180 24760 9186 24812
rect 9769 24803 9827 24809
rect 9769 24800 9781 24803
rect 9232 24772 9781 24800
rect 9232 24732 9260 24772
rect 9769 24769 9781 24772
rect 9815 24769 9827 24803
rect 9769 24763 9827 24769
rect 9953 24803 10011 24809
rect 9953 24769 9965 24803
rect 9999 24800 10011 24803
rect 10413 24803 10471 24809
rect 10413 24800 10425 24803
rect 9999 24772 10425 24800
rect 9999 24769 10011 24772
rect 9953 24763 10011 24769
rect 10413 24769 10425 24772
rect 10459 24769 10471 24803
rect 10413 24763 10471 24769
rect 12253 24803 12311 24809
rect 12253 24769 12265 24803
rect 12299 24769 12311 24803
rect 12253 24763 12311 24769
rect 12345 24803 12403 24809
rect 12345 24769 12357 24803
rect 12391 24800 12403 24803
rect 12618 24800 12624 24812
rect 12391 24772 12624 24800
rect 12391 24769 12403 24772
rect 12345 24763 12403 24769
rect 9048 24704 9260 24732
rect 5166 24556 5172 24608
rect 5224 24596 5230 24608
rect 8202 24596 8208 24608
rect 5224 24568 8208 24596
rect 5224 24556 5230 24568
rect 8202 24556 8208 24568
rect 8260 24596 8266 24608
rect 9048 24596 9076 24704
rect 9582 24692 9588 24744
rect 9640 24732 9646 24744
rect 9968 24732 9996 24763
rect 9640 24704 9996 24732
rect 9640 24692 9646 24704
rect 9122 24624 9128 24676
rect 9180 24664 9186 24676
rect 12268 24664 12296 24763
rect 12618 24760 12624 24772
rect 12676 24760 12682 24812
rect 12894 24800 12900 24812
rect 12855 24772 12900 24800
rect 12894 24760 12900 24772
rect 12952 24760 12958 24812
rect 13173 24803 13231 24809
rect 13173 24769 13185 24803
rect 13219 24800 13231 24803
rect 13446 24800 13452 24812
rect 13219 24772 13452 24800
rect 13219 24769 13231 24772
rect 13173 24763 13231 24769
rect 13446 24760 13452 24772
rect 13504 24760 13510 24812
rect 16592 24732 16620 24840
rect 19334 24828 19340 24880
rect 19392 24868 19398 24880
rect 20438 24868 20444 24880
rect 19392 24840 20444 24868
rect 19392 24828 19398 24840
rect 20438 24828 20444 24840
rect 20496 24828 20502 24880
rect 22278 24828 22284 24880
rect 22336 24868 22342 24880
rect 24688 24868 24716 24908
rect 24765 24905 24777 24939
rect 24811 24936 24823 24939
rect 24854 24936 24860 24948
rect 24811 24908 24860 24936
rect 24811 24905 24823 24908
rect 24765 24899 24823 24905
rect 24854 24896 24860 24908
rect 24912 24896 24918 24948
rect 25774 24868 25780 24880
rect 22336 24840 22876 24868
rect 24688 24840 25780 24868
rect 22336 24828 22342 24840
rect 22848 24812 22876 24840
rect 25774 24828 25780 24840
rect 25832 24828 25838 24880
rect 32306 24828 32312 24880
rect 32364 24868 32370 24880
rect 32364 24840 32812 24868
rect 32364 24828 32370 24840
rect 16850 24800 16856 24812
rect 16811 24772 16856 24800
rect 16850 24760 16856 24772
rect 16908 24760 16914 24812
rect 17034 24800 17040 24812
rect 16995 24772 17040 24800
rect 17034 24760 17040 24772
rect 17092 24760 17098 24812
rect 17218 24800 17224 24812
rect 17179 24772 17224 24800
rect 17218 24760 17224 24772
rect 17276 24760 17282 24812
rect 17313 24803 17371 24809
rect 17313 24769 17325 24803
rect 17359 24769 17371 24803
rect 17313 24763 17371 24769
rect 17328 24732 17356 24763
rect 18690 24760 18696 24812
rect 18748 24800 18754 24812
rect 22370 24800 22376 24812
rect 18748 24772 22376 24800
rect 18748 24760 18754 24772
rect 22370 24760 22376 24772
rect 22428 24800 22434 24812
rect 22649 24803 22707 24809
rect 22649 24800 22661 24803
rect 22428 24772 22661 24800
rect 22428 24760 22434 24772
rect 22649 24769 22661 24772
rect 22695 24769 22707 24803
rect 22830 24800 22836 24812
rect 22791 24772 22836 24800
rect 22649 24763 22707 24769
rect 22830 24760 22836 24772
rect 22888 24760 22894 24812
rect 22922 24760 22928 24812
rect 22980 24800 22986 24812
rect 23385 24803 23443 24809
rect 22980 24772 23025 24800
rect 22980 24760 22986 24772
rect 23385 24769 23397 24803
rect 23431 24800 23443 24803
rect 24578 24800 24584 24812
rect 23431 24772 24584 24800
rect 23431 24769 23443 24772
rect 23385 24763 23443 24769
rect 24578 24760 24584 24772
rect 24636 24760 24642 24812
rect 29730 24800 29736 24812
rect 29691 24772 29736 24800
rect 29730 24760 29736 24772
rect 29788 24760 29794 24812
rect 32398 24760 32404 24812
rect 32456 24800 32462 24812
rect 32784 24809 32812 24840
rect 32493 24803 32551 24809
rect 32493 24800 32505 24803
rect 32456 24772 32505 24800
rect 32456 24760 32462 24772
rect 32493 24769 32505 24772
rect 32539 24769 32551 24803
rect 32493 24763 32551 24769
rect 32677 24803 32735 24809
rect 32677 24769 32689 24803
rect 32723 24769 32735 24803
rect 32677 24763 32735 24769
rect 32769 24803 32827 24809
rect 32769 24769 32781 24803
rect 32815 24769 32827 24803
rect 32769 24763 32827 24769
rect 23658 24732 23664 24744
rect 16592 24704 17356 24732
rect 23619 24704 23664 24732
rect 23658 24692 23664 24704
rect 23716 24692 23722 24744
rect 27617 24735 27675 24741
rect 27617 24701 27629 24735
rect 27663 24732 27675 24735
rect 27798 24732 27804 24744
rect 27663 24704 27804 24732
rect 27663 24701 27675 24704
rect 27617 24695 27675 24701
rect 27798 24692 27804 24704
rect 27856 24692 27862 24744
rect 27893 24735 27951 24741
rect 27893 24701 27905 24735
rect 27939 24732 27951 24735
rect 32309 24735 32367 24741
rect 32309 24732 32321 24735
rect 27939 24704 32321 24732
rect 27939 24701 27951 24704
rect 27893 24695 27951 24701
rect 32309 24701 32321 24704
rect 32355 24701 32367 24735
rect 32309 24695 32367 24701
rect 9180 24636 12296 24664
rect 9180 24624 9186 24636
rect 30926 24624 30932 24676
rect 30984 24664 30990 24676
rect 31021 24667 31079 24673
rect 31021 24664 31033 24667
rect 30984 24636 31033 24664
rect 30984 24624 30990 24636
rect 31021 24633 31033 24636
rect 31067 24633 31079 24667
rect 31021 24627 31079 24633
rect 9214 24596 9220 24608
rect 8260 24568 9076 24596
rect 9175 24568 9220 24596
rect 8260 24556 8266 24568
rect 9214 24556 9220 24568
rect 9272 24596 9278 24608
rect 9582 24596 9588 24608
rect 9272 24568 9588 24596
rect 9272 24556 9278 24568
rect 9582 24556 9588 24568
rect 9640 24556 9646 24608
rect 22465 24599 22523 24605
rect 22465 24565 22477 24599
rect 22511 24596 22523 24599
rect 23382 24596 23388 24608
rect 22511 24568 23388 24596
rect 22511 24565 22523 24568
rect 22465 24559 22523 24565
rect 23382 24556 23388 24568
rect 23440 24556 23446 24608
rect 28902 24556 28908 24608
rect 28960 24596 28966 24608
rect 29181 24599 29239 24605
rect 29181 24596 29193 24599
rect 28960 24568 29193 24596
rect 28960 24556 28966 24568
rect 29181 24565 29193 24568
rect 29227 24596 29239 24599
rect 32692 24596 32720 24763
rect 29227 24568 32720 24596
rect 29227 24565 29239 24568
rect 29181 24559 29239 24565
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 16666 24352 16672 24404
rect 16724 24392 16730 24404
rect 16853 24395 16911 24401
rect 16853 24392 16865 24395
rect 16724 24364 16865 24392
rect 16724 24352 16730 24364
rect 16853 24361 16865 24364
rect 16899 24361 16911 24395
rect 16853 24355 16911 24361
rect 22830 24352 22836 24404
rect 22888 24392 22894 24404
rect 24026 24392 24032 24404
rect 22888 24364 23704 24392
rect 23987 24364 24032 24392
rect 22888 24352 22894 24364
rect 23676 24256 23704 24364
rect 24026 24352 24032 24364
rect 24084 24352 24090 24404
rect 27249 24395 27307 24401
rect 27249 24361 27261 24395
rect 27295 24392 27307 24395
rect 27614 24392 27620 24404
rect 27295 24364 27620 24392
rect 27295 24361 27307 24364
rect 27249 24355 27307 24361
rect 27614 24352 27620 24364
rect 27672 24352 27678 24404
rect 31202 24352 31208 24404
rect 31260 24392 31266 24404
rect 31389 24395 31447 24401
rect 31389 24392 31401 24395
rect 31260 24364 31401 24392
rect 31260 24352 31266 24364
rect 31389 24361 31401 24364
rect 31435 24361 31447 24395
rect 31389 24355 31447 24361
rect 24854 24284 24860 24336
rect 24912 24324 24918 24336
rect 29822 24324 29828 24336
rect 24912 24296 29828 24324
rect 24912 24284 24918 24296
rect 29822 24284 29828 24296
rect 29880 24284 29886 24336
rect 24949 24259 25007 24265
rect 24949 24256 24961 24259
rect 23676 24228 24961 24256
rect 24949 24225 24961 24228
rect 24995 24225 25007 24259
rect 26418 24256 26424 24268
rect 26331 24228 26424 24256
rect 24949 24219 25007 24225
rect 26418 24216 26424 24228
rect 26476 24256 26482 24268
rect 27338 24256 27344 24268
rect 26476 24228 27344 24256
rect 26476 24216 26482 24228
rect 27338 24216 27344 24228
rect 27396 24216 27402 24268
rect 27614 24216 27620 24268
rect 27672 24256 27678 24268
rect 28074 24256 28080 24268
rect 27672 24228 28080 24256
rect 27672 24216 27678 24228
rect 15470 24188 15476 24200
rect 15431 24160 15476 24188
rect 15470 24148 15476 24160
rect 15528 24148 15534 24200
rect 15746 24197 15752 24200
rect 15740 24151 15752 24197
rect 15804 24188 15810 24200
rect 22646 24188 22652 24200
rect 15804 24160 15840 24188
rect 22607 24160 22652 24188
rect 15746 24148 15752 24151
rect 15804 24148 15810 24160
rect 22646 24148 22652 24160
rect 22704 24148 22710 24200
rect 24486 24148 24492 24200
rect 24544 24188 24550 24200
rect 24670 24188 24676 24200
rect 24544 24160 24676 24188
rect 24544 24148 24550 24160
rect 24670 24148 24676 24160
rect 24728 24148 24734 24200
rect 25869 24191 25927 24197
rect 25869 24157 25881 24191
rect 25915 24188 25927 24191
rect 25958 24188 25964 24200
rect 25915 24160 25964 24188
rect 25915 24157 25927 24160
rect 25869 24151 25927 24157
rect 25958 24148 25964 24160
rect 26016 24148 26022 24200
rect 27724 24197 27752 24228
rect 28074 24216 28080 24228
rect 28132 24216 28138 24268
rect 27433 24191 27491 24197
rect 27433 24188 27445 24191
rect 26068 24160 27445 24188
rect 20714 24080 20720 24132
rect 20772 24120 20778 24132
rect 21821 24123 21879 24129
rect 21821 24120 21833 24123
rect 20772 24092 21833 24120
rect 20772 24080 20778 24092
rect 21821 24089 21833 24092
rect 21867 24089 21879 24123
rect 22186 24120 22192 24132
rect 22147 24092 22192 24120
rect 21821 24083 21879 24089
rect 22186 24080 22192 24092
rect 22244 24080 22250 24132
rect 22462 24080 22468 24132
rect 22520 24120 22526 24132
rect 22894 24123 22952 24129
rect 22894 24120 22906 24123
rect 22520 24092 22906 24120
rect 22520 24080 22526 24092
rect 22894 24089 22906 24092
rect 22940 24089 22952 24123
rect 22894 24083 22952 24089
rect 22738 24012 22744 24064
rect 22796 24052 22802 24064
rect 26068 24052 26096 24160
rect 27433 24157 27445 24160
rect 27479 24157 27491 24191
rect 27433 24151 27491 24157
rect 27709 24191 27767 24197
rect 27709 24157 27721 24191
rect 27755 24157 27767 24191
rect 27709 24151 27767 24157
rect 27798 24148 27804 24200
rect 27856 24188 27862 24200
rect 30009 24191 30067 24197
rect 30009 24188 30021 24191
rect 27856 24160 30021 24188
rect 27856 24148 27862 24160
rect 30009 24157 30021 24160
rect 30055 24188 30067 24191
rect 32490 24188 32496 24200
rect 30055 24160 32496 24188
rect 30055 24157 30067 24160
rect 30009 24151 30067 24157
rect 32490 24148 32496 24160
rect 32548 24148 32554 24200
rect 26142 24080 26148 24132
rect 26200 24120 26206 24132
rect 27617 24123 27675 24129
rect 26200 24080 26234 24120
rect 27617 24089 27629 24123
rect 27663 24120 27675 24123
rect 28718 24120 28724 24132
rect 27663 24092 28724 24120
rect 27663 24089 27675 24092
rect 27617 24083 27675 24089
rect 28718 24080 28724 24092
rect 28776 24080 28782 24132
rect 30276 24123 30334 24129
rect 30276 24089 30288 24123
rect 30322 24120 30334 24123
rect 30834 24120 30840 24132
rect 30322 24092 30840 24120
rect 30322 24089 30334 24092
rect 30276 24083 30334 24089
rect 30834 24080 30840 24092
rect 30892 24080 30898 24132
rect 22796 24024 26096 24052
rect 26206 24052 26234 24080
rect 31754 24052 31760 24064
rect 26206 24024 31760 24052
rect 22796 24012 22802 24024
rect 31754 24012 31760 24024
rect 31812 24052 31818 24064
rect 32398 24052 32404 24064
rect 31812 24024 32404 24052
rect 31812 24012 31818 24024
rect 32398 24012 32404 24024
rect 32456 24012 32462 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 22462 23848 22468 23860
rect 22423 23820 22468 23848
rect 22462 23808 22468 23820
rect 22520 23808 22526 23860
rect 22833 23851 22891 23857
rect 22833 23817 22845 23851
rect 22879 23848 22891 23851
rect 23474 23848 23480 23860
rect 22879 23820 23480 23848
rect 22879 23817 22891 23820
rect 22833 23811 22891 23817
rect 23474 23808 23480 23820
rect 23532 23808 23538 23860
rect 27801 23851 27859 23857
rect 27801 23817 27813 23851
rect 27847 23848 27859 23851
rect 29730 23848 29736 23860
rect 27847 23820 29736 23848
rect 27847 23817 27859 23820
rect 27801 23811 27859 23817
rect 29730 23808 29736 23820
rect 29788 23808 29794 23860
rect 14366 23780 14372 23792
rect 14214 23752 14372 23780
rect 14366 23740 14372 23752
rect 14424 23740 14430 23792
rect 21358 23780 21364 23792
rect 20272 23752 21364 23780
rect 20272 23724 20300 23752
rect 21358 23740 21364 23752
rect 21416 23740 21422 23792
rect 22572 23752 22876 23780
rect 12710 23712 12716 23724
rect 12671 23684 12716 23712
rect 12710 23672 12716 23684
rect 12768 23672 12774 23724
rect 19705 23715 19763 23721
rect 19705 23681 19717 23715
rect 19751 23712 19763 23715
rect 20254 23712 20260 23724
rect 19751 23684 20260 23712
rect 19751 23681 19763 23684
rect 19705 23675 19763 23681
rect 20254 23672 20260 23684
rect 20312 23672 20318 23724
rect 20349 23715 20407 23721
rect 20349 23681 20361 23715
rect 20395 23712 20407 23715
rect 20530 23712 20536 23724
rect 20395 23684 20536 23712
rect 20395 23681 20407 23684
rect 20349 23675 20407 23681
rect 20530 23672 20536 23684
rect 20588 23712 20594 23724
rect 22572 23712 22600 23752
rect 20588 23684 22600 23712
rect 22649 23715 22707 23721
rect 20588 23672 20594 23684
rect 22649 23681 22661 23715
rect 22695 23681 22707 23715
rect 22649 23675 22707 23681
rect 12989 23647 13047 23653
rect 12989 23613 13001 23647
rect 13035 23644 13047 23647
rect 14182 23644 14188 23656
rect 13035 23616 14188 23644
rect 13035 23613 13047 23616
rect 12989 23607 13047 23613
rect 14182 23604 14188 23616
rect 14240 23604 14246 23656
rect 19794 23604 19800 23656
rect 19852 23644 19858 23656
rect 20441 23647 20499 23653
rect 20441 23644 20453 23647
rect 19852 23616 20453 23644
rect 19852 23604 19858 23616
rect 20441 23613 20453 23616
rect 20487 23613 20499 23647
rect 22664 23644 22692 23675
rect 22738 23644 22744 23656
rect 20441 23607 20499 23613
rect 20548 23616 22744 23644
rect 20548 23588 20576 23616
rect 22738 23604 22744 23616
rect 22796 23604 22802 23656
rect 22848 23644 22876 23752
rect 24670 23740 24676 23792
rect 24728 23780 24734 23792
rect 25133 23783 25191 23789
rect 25133 23780 25145 23783
rect 24728 23752 25145 23780
rect 24728 23740 24734 23752
rect 25133 23749 25145 23752
rect 25179 23780 25191 23783
rect 25179 23752 27752 23780
rect 25179 23749 25191 23752
rect 25133 23743 25191 23749
rect 22922 23672 22928 23724
rect 22980 23712 22986 23724
rect 23385 23715 23443 23721
rect 22980 23684 23022 23712
rect 22980 23672 22986 23684
rect 23385 23681 23397 23715
rect 23431 23712 23443 23715
rect 25222 23712 25228 23724
rect 23431 23684 25228 23712
rect 23431 23681 23443 23684
rect 23385 23675 23443 23681
rect 25222 23672 25228 23684
rect 25280 23672 25286 23724
rect 25685 23715 25743 23721
rect 25685 23681 25697 23715
rect 25731 23712 25743 23715
rect 26418 23712 26424 23724
rect 25731 23684 26424 23712
rect 25731 23681 25743 23684
rect 25685 23675 25743 23681
rect 26418 23672 26424 23684
rect 26476 23672 26482 23724
rect 27430 23672 27436 23724
rect 27488 23712 27494 23724
rect 27724 23721 27752 23752
rect 34532 23752 36124 23780
rect 27525 23715 27583 23721
rect 27525 23712 27537 23715
rect 27488 23684 27537 23712
rect 27488 23672 27494 23684
rect 27525 23681 27537 23684
rect 27571 23681 27583 23715
rect 27525 23675 27583 23681
rect 27709 23715 27767 23721
rect 27709 23681 27721 23715
rect 27755 23681 27767 23715
rect 27709 23675 27767 23681
rect 25961 23647 26019 23653
rect 25961 23644 25973 23647
rect 22848 23616 25973 23644
rect 25961 23613 25973 23616
rect 26007 23644 26019 23647
rect 26234 23644 26240 23656
rect 26007 23616 26240 23644
rect 26007 23613 26019 23616
rect 25961 23607 26019 23613
rect 26234 23604 26240 23616
rect 26292 23604 26298 23656
rect 32950 23604 32956 23656
rect 33008 23644 33014 23656
rect 34532 23653 34560 23752
rect 34793 23715 34851 23721
rect 34793 23681 34805 23715
rect 34839 23712 34851 23715
rect 35986 23712 35992 23724
rect 34839 23684 35992 23712
rect 34839 23681 34851 23684
rect 34793 23675 34851 23681
rect 35986 23672 35992 23684
rect 36044 23672 36050 23724
rect 36096 23721 36124 23752
rect 36081 23715 36139 23721
rect 36081 23681 36093 23715
rect 36127 23681 36139 23715
rect 36081 23675 36139 23681
rect 34517 23647 34575 23653
rect 34517 23644 34529 23647
rect 33008 23616 34529 23644
rect 33008 23604 33014 23616
rect 34517 23613 34529 23616
rect 34563 23613 34575 23647
rect 34517 23607 34575 23613
rect 34606 23604 34612 23656
rect 34664 23644 34670 23656
rect 35345 23647 35403 23653
rect 35345 23644 35357 23647
rect 34664 23616 35357 23644
rect 34664 23604 34670 23616
rect 35345 23613 35357 23616
rect 35391 23613 35403 23647
rect 35345 23607 35403 23613
rect 17034 23536 17040 23588
rect 17092 23576 17098 23588
rect 20530 23576 20536 23588
rect 17092 23548 20536 23576
rect 17092 23536 17098 23548
rect 20530 23536 20536 23548
rect 20588 23536 20594 23588
rect 8018 23468 8024 23520
rect 8076 23508 8082 23520
rect 14461 23511 14519 23517
rect 14461 23508 14473 23511
rect 8076 23480 14473 23508
rect 8076 23468 8082 23480
rect 14461 23477 14473 23480
rect 14507 23477 14519 23511
rect 14461 23471 14519 23477
rect 19797 23511 19855 23517
rect 19797 23477 19809 23511
rect 19843 23508 19855 23511
rect 19978 23508 19984 23520
rect 19843 23480 19984 23508
rect 19843 23477 19855 23480
rect 19797 23471 19855 23477
rect 19978 23468 19984 23480
rect 20036 23468 20042 23520
rect 36078 23468 36084 23520
rect 36136 23508 36142 23520
rect 36265 23511 36323 23517
rect 36265 23508 36277 23511
rect 36136 23480 36277 23508
rect 36136 23468 36142 23480
rect 36265 23477 36277 23480
rect 36311 23477 36323 23511
rect 36265 23471 36323 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 4154 23264 4160 23316
rect 4212 23304 4218 23316
rect 4614 23304 4620 23316
rect 4212 23276 4620 23304
rect 4212 23264 4218 23276
rect 4614 23264 4620 23276
rect 4672 23264 4678 23316
rect 7377 23307 7435 23313
rect 7377 23273 7389 23307
rect 7423 23304 7435 23307
rect 7834 23304 7840 23316
rect 7423 23276 7840 23304
rect 7423 23273 7435 23276
rect 7377 23267 7435 23273
rect 7834 23264 7840 23276
rect 7892 23264 7898 23316
rect 14366 23304 14372 23316
rect 14327 23276 14372 23304
rect 14366 23264 14372 23276
rect 14424 23264 14430 23316
rect 19429 23307 19487 23313
rect 19429 23273 19441 23307
rect 19475 23304 19487 23307
rect 20346 23304 20352 23316
rect 19475 23276 20352 23304
rect 19475 23273 19487 23276
rect 19429 23267 19487 23273
rect 20346 23264 20352 23276
rect 20404 23264 20410 23316
rect 20622 23264 20628 23316
rect 20680 23304 20686 23316
rect 23201 23307 23259 23313
rect 20680 23276 20944 23304
rect 20680 23264 20686 23276
rect 3973 23239 4031 23245
rect 3973 23205 3985 23239
rect 4019 23236 4031 23239
rect 4706 23236 4712 23248
rect 4019 23208 4712 23236
rect 4019 23205 4031 23208
rect 3973 23199 4031 23205
rect 4706 23196 4712 23208
rect 4764 23196 4770 23248
rect 4798 23196 4804 23248
rect 4856 23236 4862 23248
rect 11882 23236 11888 23248
rect 4856 23208 11888 23236
rect 4856 23196 4862 23208
rect 11882 23196 11888 23208
rect 11940 23196 11946 23248
rect 17770 23236 17776 23248
rect 16546 23208 17776 23236
rect 3602 23128 3608 23180
rect 3660 23168 3666 23180
rect 3660 23140 4568 23168
rect 3660 23128 3666 23140
rect 3234 23060 3240 23112
rect 3292 23100 3298 23112
rect 4540 23109 4568 23140
rect 10962 23128 10968 23180
rect 11020 23168 11026 23180
rect 13449 23171 13507 23177
rect 13449 23168 13461 23171
rect 11020 23140 13461 23168
rect 11020 23128 11026 23140
rect 13449 23137 13461 23140
rect 13495 23168 13507 23171
rect 16546 23168 16574 23208
rect 17770 23196 17776 23208
rect 17828 23196 17834 23248
rect 20162 23196 20168 23248
rect 20220 23236 20226 23248
rect 20220 23208 20852 23236
rect 20220 23196 20226 23208
rect 13495 23140 16574 23168
rect 19705 23171 19763 23177
rect 13495 23137 13507 23140
rect 13449 23131 13507 23137
rect 19705 23137 19717 23171
rect 19751 23168 19763 23171
rect 19794 23168 19800 23180
rect 19751 23140 19800 23168
rect 19751 23137 19763 23140
rect 19705 23131 19763 23137
rect 19794 23128 19800 23140
rect 19852 23128 19858 23180
rect 20070 23128 20076 23180
rect 20128 23168 20134 23180
rect 20824 23177 20852 23208
rect 20916 23177 20944 23276
rect 23201 23273 23213 23307
rect 23247 23304 23259 23307
rect 23658 23304 23664 23316
rect 23247 23276 23664 23304
rect 23247 23273 23259 23276
rect 23201 23267 23259 23273
rect 23658 23264 23664 23276
rect 23716 23264 23722 23316
rect 25222 23264 25228 23316
rect 25280 23304 25286 23316
rect 26050 23304 26056 23316
rect 25280 23276 26056 23304
rect 25280 23264 25286 23276
rect 26050 23264 26056 23276
rect 26108 23304 26114 23316
rect 27801 23307 27859 23313
rect 27801 23304 27813 23307
rect 26108 23276 27813 23304
rect 26108 23264 26114 23276
rect 27801 23273 27813 23276
rect 27847 23273 27859 23307
rect 32490 23304 32496 23316
rect 32451 23276 32496 23304
rect 27801 23267 27859 23273
rect 32490 23264 32496 23276
rect 32548 23264 32554 23316
rect 25958 23236 25964 23248
rect 25919 23208 25964 23236
rect 25958 23196 25964 23208
rect 26016 23196 26022 23248
rect 36170 23236 36176 23248
rect 35820 23208 36176 23236
rect 20809 23171 20867 23177
rect 20128 23140 20173 23168
rect 20128 23128 20134 23140
rect 20809 23137 20821 23171
rect 20855 23137 20867 23171
rect 20809 23131 20867 23137
rect 20901 23171 20959 23177
rect 20901 23137 20913 23171
rect 20947 23137 20959 23171
rect 20901 23131 20959 23137
rect 22922 23128 22928 23180
rect 22980 23168 22986 23180
rect 35820 23177 35848 23208
rect 36170 23196 36176 23208
rect 36228 23196 36234 23248
rect 35805 23171 35863 23177
rect 22980 23140 23704 23168
rect 22980 23128 22986 23140
rect 4525 23103 4583 23109
rect 3292 23072 4292 23100
rect 3292 23060 3298 23072
rect 4154 23032 4160 23044
rect 4115 23004 4160 23032
rect 4154 22992 4160 23004
rect 4212 22992 4218 23044
rect 4264 22973 4292 23072
rect 4525 23069 4537 23103
rect 4571 23069 4583 23103
rect 4525 23063 4583 23069
rect 5350 23060 5356 23112
rect 5408 23100 5414 23112
rect 12529 23103 12587 23109
rect 12529 23100 12541 23103
rect 5408 23072 12541 23100
rect 5408 23060 5414 23072
rect 12529 23069 12541 23072
rect 12575 23069 12587 23103
rect 12986 23100 12992 23112
rect 12947 23072 12992 23100
rect 12529 23063 12587 23069
rect 12986 23060 12992 23072
rect 13044 23060 13050 23112
rect 13170 23100 13176 23112
rect 13131 23072 13176 23100
rect 13170 23060 13176 23072
rect 13228 23060 13234 23112
rect 13541 23103 13599 23109
rect 13541 23069 13553 23103
rect 13587 23069 13599 23103
rect 14274 23100 14280 23112
rect 14235 23072 14280 23100
rect 13541 23063 13599 23069
rect 7650 23032 7656 23044
rect 7611 23004 7656 23032
rect 7650 22992 7656 23004
rect 7708 22992 7714 23044
rect 7926 23032 7932 23044
rect 7887 23004 7932 23032
rect 7926 22992 7932 23004
rect 7984 22992 7990 23044
rect 12802 22992 12808 23044
rect 12860 23032 12866 23044
rect 13556 23032 13584 23063
rect 14274 23060 14280 23072
rect 14332 23060 14338 23112
rect 14366 23060 14372 23112
rect 14424 23100 14430 23112
rect 14461 23103 14519 23109
rect 14461 23100 14473 23103
rect 14424 23072 14473 23100
rect 14424 23060 14430 23072
rect 14461 23069 14473 23072
rect 14507 23100 14519 23103
rect 14550 23100 14556 23112
rect 14507 23072 14556 23100
rect 14507 23069 14519 23072
rect 14461 23063 14519 23069
rect 14550 23060 14556 23072
rect 14608 23060 14614 23112
rect 19334 23060 19340 23112
rect 19392 23100 19398 23112
rect 19613 23103 19671 23109
rect 19613 23100 19625 23103
rect 19392 23072 19625 23100
rect 19392 23060 19398 23072
rect 19613 23069 19625 23072
rect 19659 23069 19671 23103
rect 20622 23100 20628 23112
rect 19613 23063 19671 23069
rect 19904 23072 20628 23100
rect 14182 23032 14188 23044
rect 12860 23004 14188 23032
rect 12860 22992 12866 23004
rect 14182 22992 14188 23004
rect 14240 22992 14246 23044
rect 14292 23032 14320 23060
rect 15838 23032 15844 23044
rect 14292 23004 15844 23032
rect 15838 22992 15844 23004
rect 15896 23032 15902 23044
rect 17586 23032 17592 23044
rect 15896 23004 17592 23032
rect 15896 22992 15902 23004
rect 17586 22992 17592 23004
rect 17644 22992 17650 23044
rect 19904 23032 19932 23072
rect 20622 23060 20628 23072
rect 20680 23060 20686 23112
rect 20717 23103 20775 23109
rect 20717 23069 20729 23103
rect 20763 23069 20775 23103
rect 20717 23063 20775 23069
rect 20732 23032 20760 23063
rect 20990 23060 20996 23112
rect 21048 23100 21054 23112
rect 21048 23072 21093 23100
rect 21048 23060 21054 23072
rect 22186 23060 22192 23112
rect 22244 23100 22250 23112
rect 23385 23103 23443 23109
rect 23385 23100 23397 23103
rect 22244 23072 23397 23100
rect 22244 23060 22250 23072
rect 23385 23069 23397 23072
rect 23431 23069 23443 23103
rect 23566 23100 23572 23112
rect 23527 23072 23572 23100
rect 23385 23063 23443 23069
rect 19812 23004 19932 23032
rect 19996 23004 20760 23032
rect 4249 22967 4307 22973
rect 4249 22933 4261 22967
rect 4295 22933 4307 22967
rect 4249 22927 4307 22933
rect 4338 22924 4344 22976
rect 4396 22964 4402 22976
rect 4396 22936 4441 22964
rect 4396 22924 4402 22936
rect 7558 22924 7564 22976
rect 7616 22964 7622 22976
rect 7742 22964 7748 22976
rect 7616 22936 7748 22964
rect 7616 22924 7622 22936
rect 7742 22924 7748 22936
rect 7800 22964 7806 22976
rect 19812 22973 19840 23004
rect 19996 22976 20024 23004
rect 7837 22967 7895 22973
rect 7837 22964 7849 22967
rect 7800 22936 7849 22964
rect 7800 22924 7806 22936
rect 7837 22933 7849 22936
rect 7883 22933 7895 22967
rect 7837 22927 7895 22933
rect 19797 22967 19855 22973
rect 19797 22933 19809 22967
rect 19843 22933 19855 22967
rect 19978 22964 19984 22976
rect 19939 22936 19984 22964
rect 19797 22927 19855 22933
rect 19978 22924 19984 22936
rect 20036 22924 20042 22976
rect 20533 22967 20591 22973
rect 20533 22933 20545 22967
rect 20579 22964 20591 22967
rect 22554 22964 22560 22976
rect 20579 22936 22560 22964
rect 20579 22933 20591 22936
rect 20533 22927 20591 22933
rect 22554 22924 22560 22936
rect 22612 22924 22618 22976
rect 23400 22964 23428 23063
rect 23566 23060 23572 23072
rect 23624 23060 23630 23112
rect 23676 23109 23704 23140
rect 35805 23137 35817 23171
rect 35851 23137 35863 23171
rect 35805 23131 35863 23137
rect 35986 23128 35992 23180
rect 36044 23168 36050 23180
rect 36449 23171 36507 23177
rect 36449 23168 36461 23171
rect 36044 23140 36461 23168
rect 36044 23128 36050 23140
rect 36449 23137 36461 23140
rect 36495 23137 36507 23171
rect 36449 23131 36507 23137
rect 23661 23103 23719 23109
rect 23661 23069 23673 23103
rect 23707 23100 23719 23103
rect 24026 23100 24032 23112
rect 23707 23072 24032 23100
rect 23707 23069 23719 23072
rect 23661 23063 23719 23069
rect 24026 23060 24032 23072
rect 24084 23060 24090 23112
rect 24578 23100 24584 23112
rect 24539 23072 24584 23100
rect 24578 23060 24584 23072
rect 24636 23060 24642 23112
rect 30926 23060 30932 23112
rect 30984 23100 30990 23112
rect 31205 23103 31263 23109
rect 31205 23100 31217 23103
rect 30984 23072 31217 23100
rect 30984 23060 30990 23072
rect 31205 23069 31217 23072
rect 31251 23069 31263 23103
rect 31205 23063 31263 23069
rect 35897 23103 35955 23109
rect 35897 23069 35909 23103
rect 35943 23100 35955 23103
rect 36354 23100 36360 23112
rect 35943 23072 36360 23100
rect 35943 23069 35955 23072
rect 35897 23063 35955 23069
rect 36354 23060 36360 23072
rect 36412 23060 36418 23112
rect 24848 23035 24906 23041
rect 24848 23001 24860 23035
rect 24894 23032 24906 23035
rect 25866 23032 25872 23044
rect 24894 23004 25872 23032
rect 24894 23001 24906 23004
rect 24848 22995 24906 23001
rect 25866 22992 25872 23004
rect 25924 22992 25930 23044
rect 26510 23032 26516 23044
rect 26471 23004 26516 23032
rect 26510 22992 26516 23004
rect 26568 22992 26574 23044
rect 26142 22964 26148 22976
rect 23400 22936 26148 22964
rect 26142 22924 26148 22936
rect 26200 22924 26206 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 2958 22720 2964 22772
rect 3016 22760 3022 22772
rect 4338 22760 4344 22772
rect 3016 22732 4344 22760
rect 3016 22720 3022 22732
rect 4338 22720 4344 22732
rect 4396 22720 4402 22772
rect 4985 22763 5043 22769
rect 4985 22729 4997 22763
rect 5031 22760 5043 22763
rect 7650 22760 7656 22772
rect 5031 22732 7656 22760
rect 5031 22729 5043 22732
rect 4985 22723 5043 22729
rect 7650 22720 7656 22732
rect 7708 22760 7714 22772
rect 8294 22760 8300 22772
rect 7708 22732 8300 22760
rect 7708 22720 7714 22732
rect 8294 22720 8300 22732
rect 8352 22720 8358 22772
rect 8386 22720 8392 22772
rect 8444 22760 8450 22772
rect 8665 22763 8723 22769
rect 8665 22760 8677 22763
rect 8444 22732 8677 22760
rect 8444 22720 8450 22732
rect 8665 22729 8677 22732
rect 8711 22729 8723 22763
rect 8665 22723 8723 22729
rect 11882 22720 11888 22772
rect 11940 22760 11946 22772
rect 14366 22760 14372 22772
rect 11940 22732 14372 22760
rect 11940 22720 11946 22732
rect 14366 22720 14372 22732
rect 14424 22720 14430 22772
rect 16850 22720 16856 22772
rect 16908 22760 16914 22772
rect 17773 22763 17831 22769
rect 17773 22760 17785 22763
rect 16908 22732 17785 22760
rect 16908 22720 16914 22732
rect 17773 22729 17785 22732
rect 17819 22729 17831 22763
rect 20622 22760 20628 22772
rect 17773 22723 17831 22729
rect 20180 22732 20628 22760
rect 3510 22692 3516 22704
rect 3471 22664 3516 22692
rect 3510 22652 3516 22664
rect 3568 22652 3574 22704
rect 8018 22692 8024 22704
rect 7979 22664 8024 22692
rect 8018 22652 8024 22664
rect 8076 22652 8082 22704
rect 4614 22584 4620 22636
rect 4672 22584 4678 22636
rect 5718 22584 5724 22636
rect 5776 22624 5782 22636
rect 6549 22627 6607 22633
rect 6549 22624 6561 22627
rect 5776 22596 6561 22624
rect 5776 22584 5782 22596
rect 6549 22593 6561 22596
rect 6595 22593 6607 22627
rect 7006 22624 7012 22636
rect 6967 22596 7012 22624
rect 6549 22587 6607 22593
rect 7006 22584 7012 22596
rect 7064 22584 7070 22636
rect 7374 22624 7380 22636
rect 7335 22596 7380 22624
rect 7374 22584 7380 22596
rect 7432 22584 7438 22636
rect 8202 22633 8208 22636
rect 8168 22627 8208 22633
rect 8168 22593 8180 22627
rect 8168 22587 8208 22593
rect 8202 22584 8208 22587
rect 8260 22584 8266 22636
rect 8404 22624 8432 22720
rect 14274 22692 14280 22704
rect 11808 22664 14280 22692
rect 11808 22633 11836 22664
rect 14274 22652 14280 22664
rect 14332 22652 14338 22704
rect 14737 22695 14795 22701
rect 14737 22661 14749 22695
rect 14783 22692 14795 22695
rect 15470 22692 15476 22704
rect 14783 22664 15476 22692
rect 14783 22661 14795 22664
rect 14737 22655 14795 22661
rect 15470 22652 15476 22664
rect 15528 22652 15534 22704
rect 17586 22692 17592 22704
rect 17547 22664 17592 22692
rect 17586 22652 17592 22664
rect 17644 22652 17650 22704
rect 18874 22652 18880 22704
rect 18932 22692 18938 22704
rect 19337 22695 19395 22701
rect 19337 22692 19349 22695
rect 18932 22664 19349 22692
rect 18932 22652 18938 22664
rect 19337 22661 19349 22664
rect 19383 22661 19395 22695
rect 19337 22655 19395 22661
rect 19429 22695 19487 22701
rect 19429 22661 19441 22695
rect 19475 22692 19487 22695
rect 19978 22692 19984 22704
rect 19475 22664 19984 22692
rect 19475 22661 19487 22664
rect 19429 22655 19487 22661
rect 19978 22652 19984 22664
rect 20036 22652 20042 22704
rect 8312 22596 8432 22624
rect 9677 22627 9735 22633
rect 3237 22559 3295 22565
rect 3237 22525 3249 22559
rect 3283 22556 3295 22559
rect 3602 22556 3608 22568
rect 3283 22528 3608 22556
rect 3283 22525 3295 22528
rect 3237 22519 3295 22525
rect 3602 22516 3608 22528
rect 3660 22516 3666 22568
rect 7469 22559 7527 22565
rect 7469 22525 7481 22559
rect 7515 22556 7527 22559
rect 8312 22556 8340 22596
rect 9677 22593 9689 22627
rect 9723 22593 9735 22627
rect 9677 22587 9735 22593
rect 11793 22627 11851 22633
rect 11793 22593 11805 22627
rect 11839 22593 11851 22627
rect 11793 22587 11851 22593
rect 7515 22528 8340 22556
rect 7515 22525 7527 22528
rect 7469 22519 7527 22525
rect 8386 22516 8392 22568
rect 8444 22556 8450 22568
rect 9582 22556 9588 22568
rect 8444 22528 9588 22556
rect 8444 22516 8450 22528
rect 9582 22516 9588 22528
rect 9640 22516 9646 22568
rect 7098 22448 7104 22500
rect 7156 22488 7162 22500
rect 9692 22488 9720 22587
rect 11882 22584 11888 22636
rect 11940 22624 11946 22636
rect 12989 22627 13047 22633
rect 11940 22596 11985 22624
rect 11940 22584 11946 22596
rect 12989 22593 13001 22627
rect 13035 22624 13047 22627
rect 16574 22624 16580 22636
rect 13035 22596 16580 22624
rect 13035 22593 13047 22596
rect 12989 22587 13047 22593
rect 16574 22584 16580 22596
rect 16632 22584 16638 22636
rect 18509 22627 18567 22633
rect 18509 22593 18521 22627
rect 18555 22624 18567 22627
rect 19058 22624 19064 22636
rect 18555 22596 19064 22624
rect 18555 22593 18567 22596
rect 18509 22587 18567 22593
rect 19058 22584 19064 22596
rect 19116 22584 19122 22636
rect 20180 22633 20208 22732
rect 20622 22720 20628 22732
rect 20680 22720 20686 22772
rect 25866 22760 25872 22772
rect 25827 22732 25872 22760
rect 25866 22720 25872 22732
rect 25924 22720 25930 22772
rect 26234 22720 26240 22772
rect 26292 22760 26298 22772
rect 26292 22732 26337 22760
rect 26292 22720 26298 22732
rect 27522 22720 27528 22772
rect 27580 22760 27586 22772
rect 29825 22763 29883 22769
rect 29825 22760 29837 22763
rect 27580 22732 29837 22760
rect 27580 22720 27586 22732
rect 29825 22729 29837 22732
rect 29871 22729 29883 22763
rect 36354 22760 36360 22772
rect 36315 22732 36360 22760
rect 29825 22723 29883 22729
rect 36354 22720 36360 22732
rect 36412 22720 36418 22772
rect 20349 22695 20407 22701
rect 20349 22661 20361 22695
rect 20395 22692 20407 22695
rect 21082 22692 21088 22704
rect 20395 22664 21088 22692
rect 20395 22661 20407 22664
rect 20349 22655 20407 22661
rect 21082 22652 21088 22664
rect 21140 22652 21146 22704
rect 31018 22692 31024 22704
rect 26068 22664 31024 22692
rect 20165 22627 20223 22633
rect 20165 22593 20177 22627
rect 20211 22593 20223 22627
rect 20438 22624 20444 22636
rect 20399 22596 20444 22624
rect 20165 22587 20223 22593
rect 20438 22584 20444 22596
rect 20496 22584 20502 22636
rect 23661 22627 23719 22633
rect 23661 22593 23673 22627
rect 23707 22624 23719 22627
rect 24854 22624 24860 22636
rect 23707 22596 24860 22624
rect 23707 22593 23719 22596
rect 23661 22587 23719 22593
rect 24854 22584 24860 22596
rect 24912 22584 24918 22636
rect 25774 22584 25780 22636
rect 25832 22624 25838 22636
rect 26068 22633 26096 22664
rect 31018 22652 31024 22664
rect 31076 22652 31082 22704
rect 35544 22664 36308 22692
rect 26053 22627 26111 22633
rect 26053 22624 26065 22627
rect 25832 22596 26065 22624
rect 25832 22584 25838 22596
rect 26053 22593 26065 22596
rect 26099 22593 26111 22627
rect 26326 22624 26332 22636
rect 26239 22596 26332 22624
rect 26053 22587 26111 22593
rect 26326 22584 26332 22596
rect 26384 22624 26390 22636
rect 27614 22624 27620 22636
rect 26384 22596 27620 22624
rect 26384 22584 26390 22596
rect 27614 22584 27620 22596
rect 27672 22584 27678 22636
rect 27801 22627 27859 22633
rect 27801 22593 27813 22627
rect 27847 22593 27859 22627
rect 27801 22587 27859 22593
rect 12066 22556 12072 22568
rect 12027 22528 12072 22556
rect 12066 22516 12072 22528
rect 12124 22516 12130 22568
rect 18969 22559 19027 22565
rect 18969 22525 18981 22559
rect 19015 22525 19027 22559
rect 18969 22519 19027 22525
rect 27709 22559 27767 22565
rect 27709 22525 27721 22559
rect 27755 22525 27767 22559
rect 27816 22556 27844 22587
rect 27890 22584 27896 22636
rect 27948 22624 27954 22636
rect 28077 22627 28135 22633
rect 28077 22624 28089 22627
rect 27948 22596 28089 22624
rect 27948 22584 27954 22596
rect 28077 22593 28089 22596
rect 28123 22593 28135 22627
rect 28077 22587 28135 22593
rect 28166 22584 28172 22636
rect 28224 22624 28230 22636
rect 29914 22624 29920 22636
rect 28224 22596 28269 22624
rect 29875 22596 29920 22624
rect 28224 22584 28230 22596
rect 29914 22584 29920 22596
rect 29972 22584 29978 22636
rect 30469 22627 30527 22633
rect 30469 22593 30481 22627
rect 30515 22624 30527 22627
rect 30926 22624 30932 22636
rect 30515 22596 30932 22624
rect 30515 22593 30527 22596
rect 30469 22587 30527 22593
rect 30926 22584 30932 22596
rect 30984 22584 30990 22636
rect 33318 22624 33324 22636
rect 33279 22596 33324 22624
rect 33318 22584 33324 22596
rect 33376 22584 33382 22636
rect 33410 22584 33416 22636
rect 33468 22624 33474 22636
rect 35544 22633 35572 22664
rect 36280 22636 36308 22664
rect 35529 22627 35587 22633
rect 33468 22596 33513 22624
rect 33468 22584 33474 22596
rect 35529 22593 35541 22627
rect 35575 22593 35587 22627
rect 35529 22587 35587 22593
rect 35621 22627 35679 22633
rect 35621 22593 35633 22627
rect 35667 22593 35679 22627
rect 35621 22587 35679 22593
rect 35713 22627 35771 22633
rect 35713 22593 35725 22627
rect 35759 22624 35771 22627
rect 36078 22624 36084 22636
rect 35759 22596 36084 22624
rect 35759 22593 35771 22596
rect 35713 22587 35771 22593
rect 29546 22556 29552 22568
rect 27816 22528 29552 22556
rect 27709 22519 27767 22525
rect 7156 22460 9720 22488
rect 7156 22448 7162 22460
rect 18874 22448 18880 22500
rect 18932 22488 18938 22500
rect 18984 22488 19012 22519
rect 27724 22488 27752 22519
rect 29546 22516 29552 22528
rect 29604 22516 29610 22568
rect 30653 22559 30711 22565
rect 30653 22525 30665 22559
rect 30699 22525 30711 22559
rect 30653 22519 30711 22525
rect 35437 22559 35495 22565
rect 35437 22525 35449 22559
rect 35483 22525 35495 22559
rect 35636 22556 35664 22587
rect 36078 22584 36084 22596
rect 36136 22584 36142 22636
rect 36262 22624 36268 22636
rect 36223 22596 36268 22624
rect 36262 22584 36268 22596
rect 36320 22584 36326 22636
rect 36449 22627 36507 22633
rect 36449 22593 36461 22627
rect 36495 22593 36507 22627
rect 36449 22587 36507 22593
rect 35894 22556 35900 22568
rect 35636 22528 35900 22556
rect 35437 22519 35495 22525
rect 27982 22488 27988 22500
rect 18932 22460 27988 22488
rect 18932 22448 18938 22460
rect 27982 22448 27988 22460
rect 28040 22448 28046 22500
rect 30668 22488 30696 22519
rect 30742 22488 30748 22500
rect 30655 22460 30748 22488
rect 30742 22448 30748 22460
rect 30800 22488 30806 22500
rect 33597 22491 33655 22497
rect 33597 22488 33609 22491
rect 30800 22460 33609 22488
rect 30800 22448 30806 22460
rect 33597 22457 33609 22460
rect 33643 22457 33655 22491
rect 35452 22488 35480 22519
rect 35894 22516 35900 22528
rect 35952 22556 35958 22568
rect 36464 22556 36492 22587
rect 35952 22528 36492 22556
rect 35952 22516 35958 22528
rect 35986 22488 35992 22500
rect 35452 22460 35992 22488
rect 33597 22451 33655 22457
rect 35986 22448 35992 22460
rect 36044 22448 36050 22500
rect 7742 22380 7748 22432
rect 7800 22420 7806 22432
rect 8297 22423 8355 22429
rect 8297 22420 8309 22423
rect 7800 22392 8309 22420
rect 7800 22380 7806 22392
rect 8297 22389 8309 22392
rect 8343 22420 8355 22423
rect 8570 22420 8576 22432
rect 8343 22392 8576 22420
rect 8343 22389 8355 22392
rect 8297 22383 8355 22389
rect 8570 22380 8576 22392
rect 8628 22380 8634 22432
rect 9766 22420 9772 22432
rect 9727 22392 9772 22420
rect 9766 22380 9772 22392
rect 9824 22380 9830 22432
rect 12986 22380 12992 22432
rect 13044 22420 13050 22432
rect 13998 22420 14004 22432
rect 13044 22392 14004 22420
rect 13044 22380 13050 22392
rect 13998 22380 14004 22392
rect 14056 22420 14062 22432
rect 17773 22423 17831 22429
rect 17773 22420 17785 22423
rect 14056 22392 17785 22420
rect 14056 22380 14062 22392
rect 17773 22389 17785 22392
rect 17819 22389 17831 22423
rect 17954 22420 17960 22432
rect 17915 22392 17960 22420
rect 17773 22383 17831 22389
rect 17954 22380 17960 22392
rect 18012 22380 18018 22432
rect 18782 22420 18788 22432
rect 18743 22392 18788 22420
rect 18782 22380 18788 22392
rect 18840 22380 18846 22432
rect 19978 22420 19984 22432
rect 19939 22392 19984 22420
rect 19978 22380 19984 22392
rect 20036 22380 20042 22432
rect 24762 22380 24768 22432
rect 24820 22420 24826 22432
rect 24949 22423 25007 22429
rect 24949 22420 24961 22423
rect 24820 22392 24961 22420
rect 24820 22380 24826 22392
rect 24949 22389 24961 22392
rect 24995 22389 25007 22423
rect 24949 22383 25007 22389
rect 27525 22423 27583 22429
rect 27525 22389 27537 22423
rect 27571 22420 27583 22423
rect 27614 22420 27620 22432
rect 27571 22392 27620 22420
rect 27571 22389 27583 22392
rect 27525 22383 27583 22389
rect 27614 22380 27620 22392
rect 27672 22380 27678 22432
rect 34514 22380 34520 22432
rect 34572 22420 34578 22432
rect 35253 22423 35311 22429
rect 35253 22420 35265 22423
rect 34572 22392 35265 22420
rect 34572 22380 34578 22392
rect 35253 22389 35265 22392
rect 35299 22389 35311 22423
rect 35253 22383 35311 22389
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 3234 22216 3240 22228
rect 3195 22188 3240 22216
rect 3234 22176 3240 22188
rect 3292 22176 3298 22228
rect 3421 22219 3479 22225
rect 3421 22185 3433 22219
rect 3467 22216 3479 22219
rect 3602 22216 3608 22228
rect 3467 22188 3608 22216
rect 3467 22185 3479 22188
rect 3421 22179 3479 22185
rect 3602 22176 3608 22188
rect 3660 22176 3666 22228
rect 7193 22219 7251 22225
rect 7193 22185 7205 22219
rect 7239 22216 7251 22219
rect 7926 22216 7932 22228
rect 7239 22188 7932 22216
rect 7239 22185 7251 22188
rect 7193 22179 7251 22185
rect 7926 22176 7932 22188
rect 7984 22176 7990 22228
rect 12710 22216 12716 22228
rect 10796 22188 12716 22216
rect 6549 22151 6607 22157
rect 6549 22117 6561 22151
rect 6595 22148 6607 22151
rect 7558 22148 7564 22160
rect 6595 22120 7564 22148
rect 6595 22117 6607 22120
rect 6549 22111 6607 22117
rect 7558 22108 7564 22120
rect 7616 22108 7622 22160
rect 8386 22148 8392 22160
rect 8312 22120 8392 22148
rect 4341 22083 4399 22089
rect 4341 22049 4353 22083
rect 4387 22080 4399 22083
rect 4614 22080 4620 22092
rect 4387 22052 4620 22080
rect 4387 22049 4399 22052
rect 4341 22043 4399 22049
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 8312 22080 8340 22120
rect 8386 22108 8392 22120
rect 8444 22108 8450 22160
rect 9766 22108 9772 22160
rect 9824 22148 9830 22160
rect 10796 22148 10824 22188
rect 12710 22176 12716 22188
rect 12768 22176 12774 22228
rect 16206 22176 16212 22228
rect 16264 22216 16270 22228
rect 16264 22188 16574 22216
rect 16264 22176 16270 22188
rect 9824 22120 10824 22148
rect 16546 22148 16574 22188
rect 19058 22176 19064 22228
rect 19116 22216 19122 22228
rect 26329 22219 26387 22225
rect 19116 22188 26234 22216
rect 19116 22176 19122 22188
rect 16850 22148 16856 22160
rect 16546 22120 16856 22148
rect 9824 22108 9830 22120
rect 7300 22052 8340 22080
rect 7300 22024 7328 22052
rect 8570 22040 8576 22092
rect 8628 22080 8634 22092
rect 9585 22083 9643 22089
rect 8628 22052 9444 22080
rect 8628 22040 8634 22052
rect 2409 22015 2467 22021
rect 2409 21981 2421 22015
rect 2455 22012 2467 22015
rect 4065 22015 4123 22021
rect 2455 21984 2774 22012
rect 2455 21981 2467 21984
rect 2409 21975 2467 21981
rect 2746 21944 2774 21984
rect 4065 21981 4077 22015
rect 4111 21981 4123 22015
rect 4065 21975 4123 21981
rect 4157 22015 4215 22021
rect 4157 21981 4169 22015
rect 4203 22012 4215 22015
rect 4430 22012 4436 22024
rect 4203 21984 4436 22012
rect 4203 21981 4215 21984
rect 4157 21975 4215 21981
rect 2958 21944 2964 21956
rect 2746 21916 2964 21944
rect 2958 21904 2964 21916
rect 3016 21944 3022 21956
rect 3053 21947 3111 21953
rect 3053 21944 3065 21947
rect 3016 21916 3065 21944
rect 3016 21904 3022 21916
rect 3053 21913 3065 21916
rect 3099 21913 3111 21947
rect 4080 21944 4108 21975
rect 4430 21972 4436 21984
rect 4488 22012 4494 22024
rect 4798 22012 4804 22024
rect 4488 21984 4804 22012
rect 4488 21972 4494 21984
rect 4798 21972 4804 21984
rect 4856 21972 4862 22024
rect 7101 22015 7159 22021
rect 7101 22012 7113 22015
rect 6104 21984 7113 22012
rect 4246 21944 4252 21956
rect 4080 21916 4252 21944
rect 3053 21907 3111 21913
rect 4246 21904 4252 21916
rect 4304 21904 4310 21956
rect 1854 21836 1860 21888
rect 1912 21876 1918 21888
rect 2501 21879 2559 21885
rect 2501 21876 2513 21879
rect 1912 21848 2513 21876
rect 1912 21836 1918 21848
rect 2501 21845 2513 21848
rect 2547 21845 2559 21879
rect 2501 21839 2559 21845
rect 3263 21879 3321 21885
rect 3263 21845 3275 21879
rect 3309 21876 3321 21879
rect 6104 21876 6132 21984
rect 7101 21981 7113 21984
rect 7147 21981 7159 22015
rect 7282 22012 7288 22024
rect 7243 21984 7288 22012
rect 7101 21975 7159 21981
rect 7282 21972 7288 21984
rect 7340 21972 7346 22024
rect 8294 22012 8300 22024
rect 8255 21984 8300 22012
rect 8294 21972 8300 21984
rect 8352 21972 8358 22024
rect 8478 22012 8484 22024
rect 8439 21984 8484 22012
rect 8478 21972 8484 21984
rect 8536 21972 8542 22024
rect 9306 22012 9312 22024
rect 9267 21984 9312 22012
rect 9306 21972 9312 21984
rect 9364 21972 9370 22024
rect 9416 22021 9444 22052
rect 9585 22049 9597 22083
rect 9631 22049 9643 22083
rect 9585 22043 9643 22049
rect 10689 22083 10747 22089
rect 10689 22049 10701 22083
rect 10735 22080 10747 22083
rect 10796 22080 10824 22120
rect 16850 22108 16856 22120
rect 16908 22108 16914 22160
rect 24854 22148 24860 22160
rect 24815 22120 24860 22148
rect 24854 22108 24860 22120
rect 24912 22108 24918 22160
rect 26206 22148 26234 22188
rect 26329 22185 26341 22219
rect 26375 22216 26387 22219
rect 26510 22216 26516 22228
rect 26375 22188 26516 22216
rect 26375 22185 26387 22188
rect 26329 22179 26387 22185
rect 26510 22176 26516 22188
rect 26568 22176 26574 22228
rect 27798 22216 27804 22228
rect 27759 22188 27804 22216
rect 27798 22176 27804 22188
rect 27856 22176 27862 22228
rect 29914 22176 29920 22228
rect 29972 22216 29978 22228
rect 30193 22219 30251 22225
rect 30193 22216 30205 22219
rect 29972 22188 30205 22216
rect 29972 22176 29978 22188
rect 30193 22185 30205 22188
rect 30239 22185 30251 22219
rect 30193 22179 30251 22185
rect 33318 22176 33324 22228
rect 33376 22216 33382 22228
rect 33781 22219 33839 22225
rect 33781 22216 33793 22219
rect 33376 22188 33793 22216
rect 33376 22176 33382 22188
rect 33781 22185 33793 22188
rect 33827 22216 33839 22219
rect 37093 22219 37151 22225
rect 37093 22216 37105 22219
rect 33827 22188 37105 22216
rect 33827 22185 33839 22188
rect 33781 22179 33839 22185
rect 37093 22185 37105 22188
rect 37139 22185 37151 22219
rect 37093 22179 37151 22185
rect 34606 22148 34612 22160
rect 26206 22120 34612 22148
rect 34606 22108 34612 22120
rect 34664 22108 34670 22160
rect 34885 22151 34943 22157
rect 34885 22117 34897 22151
rect 34931 22117 34943 22151
rect 34885 22111 34943 22117
rect 10962 22080 10968 22092
rect 10735 22052 10824 22080
rect 10923 22052 10968 22080
rect 10735 22049 10747 22052
rect 10689 22043 10747 22049
rect 9401 22015 9459 22021
rect 9401 21981 9413 22015
rect 9447 21981 9459 22015
rect 9401 21975 9459 21981
rect 6181 21947 6239 21953
rect 6181 21913 6193 21947
rect 6227 21944 6239 21947
rect 7466 21944 7472 21956
rect 6227 21916 7472 21944
rect 6227 21913 6239 21916
rect 6181 21907 6239 21913
rect 7466 21904 7472 21916
rect 7524 21944 7530 21956
rect 8018 21944 8024 21956
rect 7524 21916 8024 21944
rect 7524 21904 7530 21916
rect 8018 21904 8024 21916
rect 8076 21904 8082 21956
rect 8389 21947 8447 21953
rect 8389 21913 8401 21947
rect 8435 21944 8447 21947
rect 9600 21944 9628 22043
rect 10962 22040 10968 22052
rect 11020 22040 11026 22092
rect 16666 22080 16672 22092
rect 16040 22052 16672 22080
rect 9674 21972 9680 22024
rect 9732 22012 9738 22024
rect 9732 21984 9777 22012
rect 9732 21972 9738 21984
rect 12066 21972 12072 22024
rect 12124 21972 12130 22024
rect 14366 22012 14372 22024
rect 14327 21984 14372 22012
rect 14366 21972 14372 21984
rect 14424 21972 14430 22024
rect 15562 21972 15568 22024
rect 15620 22012 15626 22024
rect 16040 22021 16068 22052
rect 16666 22040 16672 22052
rect 16724 22040 16730 22092
rect 19334 22080 19340 22092
rect 17880 22052 19340 22080
rect 15841 22015 15899 22021
rect 15841 22012 15853 22015
rect 15620 21984 15853 22012
rect 15620 21972 15626 21984
rect 15841 21981 15853 21984
rect 15887 21981 15899 22015
rect 15841 21975 15899 21981
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 21981 16083 22015
rect 16206 22012 16212 22024
rect 16167 21984 16212 22012
rect 16025 21975 16083 21981
rect 16206 21972 16212 21984
rect 16264 21972 16270 22024
rect 16298 21972 16304 22024
rect 16356 22012 16362 22024
rect 16853 22015 16911 22021
rect 16853 22012 16865 22015
rect 16356 21984 16865 22012
rect 16356 21972 16362 21984
rect 16853 21981 16865 21984
rect 16899 21981 16911 22015
rect 17880 22012 17908 22052
rect 19334 22040 19340 22052
rect 19392 22040 19398 22092
rect 26602 22080 26608 22092
rect 26252 22052 26608 22080
rect 26252 22024 26280 22052
rect 26602 22040 26608 22052
rect 26660 22040 26666 22092
rect 27706 22080 27712 22092
rect 27667 22052 27712 22080
rect 27706 22040 27712 22052
rect 27764 22040 27770 22092
rect 29546 22040 29552 22092
rect 29604 22080 29610 22092
rect 32950 22080 32956 22092
rect 29604 22052 32812 22080
rect 32911 22052 32956 22080
rect 29604 22040 29610 22052
rect 19426 22012 19432 22024
rect 16853 21975 16911 21981
rect 17512 21984 17908 22012
rect 19387 21984 19432 22012
rect 14826 21944 14832 21956
rect 8435 21916 9628 21944
rect 14787 21916 14832 21944
rect 8435 21913 8447 21916
rect 8389 21907 8447 21913
rect 14826 21904 14832 21916
rect 14884 21904 14890 21956
rect 16117 21947 16175 21953
rect 16117 21913 16129 21947
rect 16163 21944 16175 21947
rect 16574 21944 16580 21956
rect 16163 21916 16580 21944
rect 16163 21913 16175 21916
rect 16117 21907 16175 21913
rect 16574 21904 16580 21916
rect 16632 21904 16638 21956
rect 16942 21904 16948 21956
rect 17000 21944 17006 21956
rect 17098 21947 17156 21953
rect 17098 21944 17110 21947
rect 17000 21916 17110 21944
rect 17000 21904 17006 21916
rect 17098 21913 17110 21916
rect 17144 21913 17156 21947
rect 17098 21907 17156 21913
rect 6641 21879 6699 21885
rect 6641 21876 6653 21879
rect 3309 21848 6653 21876
rect 3309 21845 3321 21848
rect 3263 21839 3321 21845
rect 6641 21845 6653 21848
rect 6687 21845 6699 21879
rect 6641 21839 6699 21845
rect 6914 21836 6920 21888
rect 6972 21876 6978 21888
rect 8202 21876 8208 21888
rect 6972 21848 8208 21876
rect 6972 21836 6978 21848
rect 8202 21836 8208 21848
rect 8260 21836 8266 21888
rect 9125 21879 9183 21885
rect 9125 21845 9137 21879
rect 9171 21876 9183 21879
rect 9766 21876 9772 21888
rect 9171 21848 9772 21876
rect 9171 21845 9183 21848
rect 9125 21839 9183 21845
rect 9766 21836 9772 21848
rect 9824 21836 9830 21888
rect 9858 21836 9864 21888
rect 9916 21876 9922 21888
rect 12437 21879 12495 21885
rect 12437 21876 12449 21879
rect 9916 21848 12449 21876
rect 9916 21836 9922 21848
rect 12437 21845 12449 21848
rect 12483 21845 12495 21879
rect 12437 21839 12495 21845
rect 16393 21879 16451 21885
rect 16393 21845 16405 21879
rect 16439 21876 16451 21879
rect 17512 21876 17540 21984
rect 19426 21972 19432 21984
rect 19484 21972 19490 22024
rect 19696 22015 19754 22021
rect 19696 21981 19708 22015
rect 19742 22012 19754 22015
rect 19978 22012 19984 22024
rect 19742 21984 19984 22012
rect 19742 21981 19754 21984
rect 19696 21975 19754 21981
rect 19978 21972 19984 21984
rect 20036 21972 20042 22024
rect 20254 21972 20260 22024
rect 20312 22012 20318 22024
rect 24581 22015 24639 22021
rect 24581 22012 24593 22015
rect 20312 21984 24593 22012
rect 20312 21972 20318 21984
rect 24581 21981 24593 21984
rect 24627 21981 24639 22015
rect 24581 21975 24639 21981
rect 24670 21972 24676 22024
rect 24728 22012 24734 22024
rect 24765 22015 24823 22021
rect 24765 22012 24777 22015
rect 24728 21984 24777 22012
rect 24728 21972 24734 21984
rect 24765 21981 24777 21984
rect 24811 21981 24823 22015
rect 26234 22012 26240 22024
rect 26195 21984 26240 22012
rect 24765 21975 24823 21981
rect 26234 21972 26240 21984
rect 26292 21972 26298 22024
rect 26421 22015 26479 22021
rect 26421 21981 26433 22015
rect 26467 21981 26479 22015
rect 27614 22012 27620 22024
rect 27575 21984 27620 22012
rect 26421 21975 26479 21981
rect 17586 21904 17592 21956
rect 17644 21944 17650 21956
rect 21910 21944 21916 21956
rect 17644 21916 19656 21944
rect 17644 21904 17650 21916
rect 16439 21848 17540 21876
rect 18233 21879 18291 21885
rect 16439 21845 16451 21848
rect 16393 21839 16451 21845
rect 18233 21845 18245 21879
rect 18279 21876 18291 21879
rect 18322 21876 18328 21888
rect 18279 21848 18328 21876
rect 18279 21845 18291 21848
rect 18233 21839 18291 21845
rect 18322 21836 18328 21848
rect 18380 21836 18386 21888
rect 19628 21876 19656 21916
rect 20180 21916 21916 21944
rect 20180 21876 20208 21916
rect 21910 21904 21916 21916
rect 21968 21944 21974 21956
rect 26436 21944 26464 21975
rect 27614 21972 27620 21984
rect 27672 21972 27678 22024
rect 29917 22015 29975 22021
rect 29917 21981 29929 22015
rect 29963 22012 29975 22015
rect 30742 22012 30748 22024
rect 29963 21984 30604 22012
rect 30703 21984 30748 22012
rect 29963 21981 29975 21984
rect 29917 21975 29975 21981
rect 21968 21916 26464 21944
rect 21968 21904 21974 21916
rect 28074 21904 28080 21956
rect 28132 21944 28138 21956
rect 28902 21944 28908 21956
rect 28132 21916 28908 21944
rect 28132 21904 28138 21916
rect 28902 21904 28908 21916
rect 28960 21944 28966 21956
rect 30101 21947 30159 21953
rect 30101 21944 30113 21947
rect 28960 21916 30113 21944
rect 28960 21904 28966 21916
rect 30101 21913 30113 21916
rect 30147 21913 30159 21947
rect 30576 21944 30604 21984
rect 30742 21972 30748 21984
rect 30800 21972 30806 22024
rect 30926 22012 30932 22024
rect 30887 21984 30932 22012
rect 30926 21972 30932 21984
rect 30984 21972 30990 22024
rect 32493 22015 32551 22021
rect 32493 22012 32505 22015
rect 31726 21984 32505 22012
rect 30837 21947 30895 21953
rect 30837 21944 30849 21947
rect 30576 21916 30849 21944
rect 30101 21907 30159 21913
rect 30837 21913 30849 21916
rect 30883 21944 30895 21947
rect 31726 21944 31754 21984
rect 32493 21981 32505 21984
rect 32539 21981 32551 22015
rect 32784 22012 32812 22052
rect 32950 22040 32956 22052
rect 33008 22040 33014 22092
rect 34900 22080 34928 22111
rect 33244 22052 34928 22080
rect 35989 22083 36047 22089
rect 33244 22012 33272 22052
rect 35989 22049 36001 22083
rect 36035 22080 36047 22083
rect 36035 22052 38056 22080
rect 36035 22049 36047 22052
rect 35989 22043 36047 22049
rect 38028 22024 38056 22052
rect 32784 21984 33272 22012
rect 33321 22015 33379 22021
rect 32493 21975 32551 21981
rect 33321 21981 33333 22015
rect 33367 22012 33379 22015
rect 33410 22012 33416 22024
rect 33367 21984 33416 22012
rect 33367 21981 33379 21984
rect 33321 21975 33379 21981
rect 33410 21972 33416 21984
rect 33468 21972 33474 22024
rect 34514 21972 34520 22024
rect 34572 22012 34578 22024
rect 35161 22015 35219 22021
rect 35161 22012 35173 22015
rect 34572 21984 35173 22012
rect 34572 21972 34578 21984
rect 35161 21981 35173 21984
rect 35207 21981 35219 22015
rect 35161 21975 35219 21981
rect 36173 22015 36231 22021
rect 36173 21981 36185 22015
rect 36219 21981 36231 22015
rect 36173 21975 36231 21981
rect 36357 22015 36415 22021
rect 36357 21981 36369 22015
rect 36403 22012 36415 22015
rect 37001 22015 37059 22021
rect 37001 22012 37013 22015
rect 36403 21984 37013 22012
rect 36403 21981 36415 21984
rect 36357 21975 36415 21981
rect 37001 21981 37013 21984
rect 37047 21981 37059 22015
rect 37001 21975 37059 21981
rect 30883 21916 31754 21944
rect 34885 21947 34943 21953
rect 30883 21913 30895 21916
rect 30837 21907 30895 21913
rect 34885 21913 34897 21947
rect 34931 21944 34943 21947
rect 35342 21944 35348 21956
rect 34931 21916 35348 21944
rect 34931 21913 34943 21916
rect 34885 21907 34943 21913
rect 35342 21904 35348 21916
rect 35400 21904 35406 21956
rect 36188 21944 36216 21975
rect 37182 21972 37188 22024
rect 37240 22012 37246 22024
rect 37829 22015 37887 22021
rect 37829 22012 37841 22015
rect 37240 21984 37841 22012
rect 37240 21972 37246 21984
rect 37829 21981 37841 21984
rect 37875 21981 37887 22015
rect 38010 22012 38016 22024
rect 37971 21984 38016 22012
rect 37829 21975 37887 21981
rect 38010 21972 38016 21984
rect 38068 21972 38074 22024
rect 36722 21944 36728 21956
rect 36188 21916 36728 21944
rect 36722 21904 36728 21916
rect 36780 21904 36786 21956
rect 36817 21947 36875 21953
rect 36817 21913 36829 21947
rect 36863 21944 36875 21947
rect 37921 21947 37979 21953
rect 37921 21944 37933 21947
rect 36863 21916 37933 21944
rect 36863 21913 36875 21916
rect 36817 21907 36875 21913
rect 37921 21913 37933 21916
rect 37967 21913 37979 21947
rect 37921 21907 37979 21913
rect 19628 21848 20208 21876
rect 20809 21879 20867 21885
rect 20809 21845 20821 21879
rect 20855 21876 20867 21879
rect 21082 21876 21088 21888
rect 20855 21848 21088 21876
rect 20855 21845 20867 21848
rect 20809 21839 20867 21845
rect 21082 21836 21088 21848
rect 21140 21876 21146 21888
rect 21358 21876 21364 21888
rect 21140 21848 21364 21876
rect 21140 21836 21146 21848
rect 21358 21836 21364 21848
rect 21416 21836 21422 21888
rect 21450 21836 21456 21888
rect 21508 21876 21514 21888
rect 27985 21879 28043 21885
rect 27985 21876 27997 21879
rect 21508 21848 27997 21876
rect 21508 21836 21514 21848
rect 27985 21845 27997 21848
rect 28031 21845 28043 21879
rect 35066 21876 35072 21888
rect 35027 21848 35072 21876
rect 27985 21839 28043 21845
rect 35066 21836 35072 21848
rect 35124 21836 35130 21888
rect 36740 21876 36768 21904
rect 37182 21876 37188 21888
rect 36740 21848 37188 21876
rect 37182 21836 37188 21848
rect 37240 21836 37246 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 6917 21675 6975 21681
rect 6917 21641 6929 21675
rect 6963 21672 6975 21675
rect 7006 21672 7012 21684
rect 6963 21644 7012 21672
rect 6963 21641 6975 21644
rect 6917 21635 6975 21641
rect 7006 21632 7012 21644
rect 7064 21632 7070 21684
rect 7374 21632 7380 21684
rect 7432 21672 7438 21684
rect 7561 21675 7619 21681
rect 7561 21672 7573 21675
rect 7432 21644 7573 21672
rect 7432 21632 7438 21644
rect 7561 21641 7573 21644
rect 7607 21641 7619 21675
rect 7561 21635 7619 21641
rect 9306 21632 9312 21684
rect 9364 21672 9370 21684
rect 9677 21675 9735 21681
rect 9677 21672 9689 21675
rect 9364 21644 9689 21672
rect 9364 21632 9370 21644
rect 9677 21641 9689 21644
rect 9723 21641 9735 21675
rect 9677 21635 9735 21641
rect 11057 21675 11115 21681
rect 11057 21641 11069 21675
rect 11103 21672 11115 21675
rect 14366 21672 14372 21684
rect 11103 21644 14372 21672
rect 11103 21641 11115 21644
rect 11057 21635 11115 21641
rect 14366 21632 14372 21644
rect 14424 21672 14430 21684
rect 20714 21672 20720 21684
rect 14424 21644 20720 21672
rect 14424 21632 14430 21644
rect 20714 21632 20720 21644
rect 20772 21632 20778 21684
rect 20806 21632 20812 21684
rect 20864 21672 20870 21684
rect 21450 21672 21456 21684
rect 20864 21644 21456 21672
rect 20864 21632 20870 21644
rect 21450 21632 21456 21644
rect 21508 21632 21514 21684
rect 24486 21672 24492 21684
rect 24447 21644 24492 21672
rect 24486 21632 24492 21644
rect 24544 21632 24550 21684
rect 34609 21675 34667 21681
rect 34609 21672 34621 21675
rect 33244 21644 34621 21672
rect 4525 21607 4583 21613
rect 4525 21604 4537 21607
rect 3358 21576 4537 21604
rect 4525 21573 4537 21576
rect 4571 21573 4583 21607
rect 7742 21604 7748 21616
rect 4525 21567 4583 21573
rect 6748 21576 7748 21604
rect 1854 21536 1860 21548
rect 1815 21508 1860 21536
rect 1854 21496 1860 21508
rect 1912 21496 1918 21548
rect 4246 21536 4252 21548
rect 4207 21508 4252 21536
rect 4246 21496 4252 21508
rect 4304 21496 4310 21548
rect 4430 21496 4436 21548
rect 4488 21536 4494 21548
rect 5074 21536 5080 21548
rect 4488 21508 5080 21536
rect 4488 21496 4494 21508
rect 5074 21496 5080 21508
rect 5132 21496 5138 21548
rect 6748 21545 6776 21576
rect 7742 21564 7748 21576
rect 7800 21564 7806 21616
rect 8110 21564 8116 21616
rect 8168 21604 8174 21616
rect 9858 21604 9864 21616
rect 8168 21576 9864 21604
rect 8168 21564 8174 21576
rect 9858 21564 9864 21576
rect 9916 21564 9922 21616
rect 15654 21564 15660 21616
rect 15712 21604 15718 21616
rect 16209 21607 16267 21613
rect 15712 21576 16160 21604
rect 15712 21564 15718 21576
rect 6733 21539 6791 21545
rect 6733 21505 6745 21539
rect 6779 21505 6791 21539
rect 7466 21536 7472 21548
rect 7427 21508 7472 21536
rect 6733 21499 6791 21505
rect 7466 21496 7472 21508
rect 7524 21496 7530 21548
rect 7558 21496 7564 21548
rect 7616 21536 7622 21548
rect 7653 21539 7711 21545
rect 7653 21536 7665 21539
rect 7616 21508 7665 21536
rect 7616 21496 7622 21508
rect 7653 21505 7665 21508
rect 7699 21536 7711 21539
rect 8128 21536 8156 21564
rect 7699 21508 8156 21536
rect 7699 21505 7711 21508
rect 7653 21499 7711 21505
rect 9122 21496 9128 21548
rect 9180 21536 9186 21548
rect 9217 21539 9275 21545
rect 9217 21536 9229 21539
rect 9180 21508 9229 21536
rect 9180 21496 9186 21508
rect 9217 21505 9229 21508
rect 9263 21505 9275 21539
rect 9217 21499 9275 21505
rect 9493 21539 9551 21545
rect 9493 21505 9505 21539
rect 9539 21536 9551 21539
rect 10226 21536 10232 21548
rect 9539 21508 10232 21536
rect 9539 21505 9551 21508
rect 9493 21499 9551 21505
rect 10226 21496 10232 21508
rect 10284 21536 10290 21548
rect 10686 21536 10692 21548
rect 10284 21508 10692 21536
rect 10284 21496 10290 21508
rect 10686 21496 10692 21508
rect 10744 21496 10750 21548
rect 10870 21536 10876 21548
rect 10831 21508 10876 21536
rect 10870 21496 10876 21508
rect 10928 21496 10934 21548
rect 10965 21539 11023 21545
rect 10965 21505 10977 21539
rect 11011 21505 11023 21539
rect 12066 21536 12072 21548
rect 12027 21508 12072 21536
rect 10965 21499 11023 21505
rect 2133 21471 2191 21477
rect 2133 21437 2145 21471
rect 2179 21468 2191 21471
rect 2774 21468 2780 21480
rect 2179 21440 2780 21468
rect 2179 21437 2191 21440
rect 2133 21431 2191 21437
rect 2774 21428 2780 21440
rect 2832 21428 2838 21480
rect 4264 21468 4292 21496
rect 4798 21468 4804 21480
rect 4264 21440 4804 21468
rect 4798 21428 4804 21440
rect 4856 21428 4862 21480
rect 5442 21428 5448 21480
rect 5500 21468 5506 21480
rect 6549 21471 6607 21477
rect 6549 21468 6561 21471
rect 5500 21440 6561 21468
rect 5500 21428 5506 21440
rect 6549 21437 6561 21440
rect 6595 21468 6607 21471
rect 7282 21468 7288 21480
rect 6595 21440 7288 21468
rect 6595 21437 6607 21440
rect 6549 21431 6607 21437
rect 7282 21428 7288 21440
rect 7340 21428 7346 21480
rect 9398 21468 9404 21480
rect 9359 21440 9404 21468
rect 9398 21428 9404 21440
rect 9456 21428 9462 21480
rect 10980 21468 11008 21499
rect 12066 21496 12072 21508
rect 12124 21496 12130 21548
rect 12989 21539 13047 21545
rect 12989 21505 13001 21539
rect 13035 21536 13047 21539
rect 13998 21536 14004 21548
rect 13035 21508 14004 21536
rect 13035 21505 13047 21508
rect 12989 21499 13047 21505
rect 13998 21496 14004 21508
rect 14056 21496 14062 21548
rect 14826 21496 14832 21548
rect 14884 21536 14890 21548
rect 16022 21536 16028 21548
rect 14884 21508 16028 21536
rect 14884 21496 14890 21508
rect 16022 21496 16028 21508
rect 16080 21496 16086 21548
rect 16132 21536 16160 21576
rect 16209 21573 16221 21607
rect 16255 21604 16267 21607
rect 16574 21604 16580 21616
rect 16255 21576 16580 21604
rect 16255 21573 16267 21576
rect 16209 21567 16267 21573
rect 16574 21564 16580 21576
rect 16632 21604 16638 21616
rect 17218 21604 17224 21616
rect 16632 21576 17224 21604
rect 16632 21564 16638 21576
rect 17218 21564 17224 21576
rect 17276 21564 17282 21616
rect 17954 21564 17960 21616
rect 18012 21604 18018 21616
rect 18233 21607 18291 21613
rect 18233 21604 18245 21607
rect 18012 21576 18245 21604
rect 18012 21564 18018 21576
rect 18233 21573 18245 21576
rect 18279 21573 18291 21607
rect 18233 21567 18291 21573
rect 20438 21564 20444 21616
rect 20496 21604 20502 21616
rect 23382 21613 23388 21616
rect 23376 21604 23388 21613
rect 20496 21576 21404 21604
rect 23343 21576 23388 21604
rect 20496 21564 20502 21576
rect 16301 21539 16359 21545
rect 16301 21536 16313 21539
rect 16132 21508 16313 21536
rect 16301 21505 16313 21508
rect 16347 21536 16359 21539
rect 16482 21536 16488 21548
rect 16347 21508 16488 21536
rect 16347 21505 16359 21508
rect 16301 21499 16359 21505
rect 16482 21496 16488 21508
rect 16540 21496 16546 21548
rect 21085 21539 21143 21545
rect 21085 21505 21097 21539
rect 21131 21505 21143 21539
rect 21266 21536 21272 21548
rect 21227 21508 21272 21536
rect 21085 21499 21143 21505
rect 12526 21468 12532 21480
rect 10980 21440 12532 21468
rect 12526 21428 12532 21440
rect 12584 21428 12590 21480
rect 13170 21428 13176 21480
rect 13228 21468 13234 21480
rect 20806 21468 20812 21480
rect 13228 21440 20812 21468
rect 13228 21428 13234 21440
rect 20806 21428 20812 21440
rect 20864 21428 20870 21480
rect 21100 21468 21128 21499
rect 21266 21496 21272 21508
rect 21324 21496 21330 21548
rect 21376 21545 21404 21576
rect 23376 21567 23388 21576
rect 23382 21564 23388 21567
rect 23440 21564 23446 21616
rect 21361 21539 21419 21545
rect 21361 21505 21373 21539
rect 21407 21536 21419 21539
rect 21542 21536 21548 21548
rect 21407 21508 21548 21536
rect 21407 21505 21419 21508
rect 21361 21499 21419 21505
rect 21542 21496 21548 21508
rect 21600 21496 21606 21548
rect 27982 21536 27988 21548
rect 27943 21508 27988 21536
rect 27982 21496 27988 21508
rect 28040 21496 28046 21548
rect 28166 21536 28172 21548
rect 28127 21508 28172 21536
rect 28166 21496 28172 21508
rect 28224 21496 28230 21548
rect 33244 21545 33272 21644
rect 34609 21641 34621 21644
rect 34655 21672 34667 21675
rect 35066 21672 35072 21684
rect 34655 21644 35072 21672
rect 34655 21641 34667 21644
rect 34609 21635 34667 21641
rect 35066 21632 35072 21644
rect 35124 21632 35130 21684
rect 36630 21564 36636 21616
rect 36688 21604 36694 21616
rect 36909 21607 36967 21613
rect 36909 21604 36921 21607
rect 36688 21576 36921 21604
rect 36688 21564 36694 21576
rect 36909 21573 36921 21576
rect 36955 21604 36967 21607
rect 38010 21604 38016 21616
rect 36955 21576 38016 21604
rect 36955 21573 36967 21576
rect 36909 21567 36967 21573
rect 38010 21564 38016 21576
rect 38068 21564 38074 21616
rect 33229 21539 33287 21545
rect 33229 21505 33241 21539
rect 33275 21505 33287 21539
rect 33229 21499 33287 21505
rect 34609 21539 34667 21545
rect 34609 21505 34621 21539
rect 34655 21536 34667 21539
rect 35894 21536 35900 21548
rect 34655 21508 35900 21536
rect 34655 21505 34667 21508
rect 34609 21499 34667 21505
rect 35894 21496 35900 21508
rect 35952 21496 35958 21548
rect 22370 21468 22376 21480
rect 21100 21440 22376 21468
rect 14918 21360 14924 21412
rect 14976 21400 14982 21412
rect 21100 21400 21128 21440
rect 22370 21428 22376 21440
rect 22428 21428 22434 21480
rect 22554 21428 22560 21480
rect 22612 21468 22618 21480
rect 23109 21471 23167 21477
rect 23109 21468 23121 21471
rect 22612 21440 23121 21468
rect 22612 21428 22618 21440
rect 23109 21437 23121 21440
rect 23155 21437 23167 21471
rect 23109 21431 23167 21437
rect 28353 21471 28411 21477
rect 28353 21437 28365 21471
rect 28399 21468 28411 21471
rect 29730 21468 29736 21480
rect 28399 21440 29736 21468
rect 28399 21437 28411 21440
rect 28353 21431 28411 21437
rect 29730 21428 29736 21440
rect 29788 21428 29794 21480
rect 33321 21471 33379 21477
rect 33321 21437 33333 21471
rect 33367 21468 33379 21471
rect 34514 21468 34520 21480
rect 33367 21440 34520 21468
rect 33367 21437 33379 21440
rect 33321 21431 33379 21437
rect 34514 21428 34520 21440
rect 34572 21428 34578 21480
rect 34790 21477 34796 21480
rect 34747 21471 34796 21477
rect 34747 21437 34759 21471
rect 34793 21437 34796 21471
rect 34747 21431 34796 21437
rect 34790 21428 34796 21431
rect 34848 21428 34854 21480
rect 34977 21471 35035 21477
rect 34977 21437 34989 21471
rect 35023 21468 35035 21471
rect 35342 21468 35348 21480
rect 35023 21440 35348 21468
rect 35023 21437 35035 21440
rect 34977 21431 35035 21437
rect 35342 21428 35348 21440
rect 35400 21428 35406 21480
rect 35802 21428 35808 21480
rect 35860 21468 35866 21480
rect 36004 21468 36032 21522
rect 35860 21440 36032 21468
rect 36081 21471 36139 21477
rect 35860 21428 35866 21440
rect 36081 21437 36093 21471
rect 36127 21468 36139 21471
rect 36170 21468 36176 21480
rect 36127 21440 36176 21468
rect 36127 21437 36139 21440
rect 36081 21431 36139 21437
rect 36170 21428 36176 21440
rect 36228 21428 36234 21480
rect 14976 21372 21128 21400
rect 14976 21360 14982 21372
rect 2866 21292 2872 21344
rect 2924 21332 2930 21344
rect 3142 21332 3148 21344
rect 2924 21304 3148 21332
rect 2924 21292 2930 21304
rect 3142 21292 3148 21304
rect 3200 21332 3206 21344
rect 3605 21335 3663 21341
rect 3605 21332 3617 21335
rect 3200 21304 3617 21332
rect 3200 21292 3206 21304
rect 3605 21301 3617 21304
rect 3651 21301 3663 21335
rect 3605 21295 3663 21301
rect 8294 21292 8300 21344
rect 8352 21332 8358 21344
rect 9214 21332 9220 21344
rect 8352 21304 9220 21332
rect 8352 21292 8358 21304
rect 9214 21292 9220 21304
rect 9272 21292 9278 21344
rect 11974 21292 11980 21344
rect 12032 21332 12038 21344
rect 12161 21335 12219 21341
rect 12161 21332 12173 21335
rect 12032 21304 12173 21332
rect 12032 21292 12038 21304
rect 12161 21301 12173 21304
rect 12207 21301 12219 21335
rect 12161 21295 12219 21301
rect 13170 21292 13176 21344
rect 13228 21332 13234 21344
rect 14277 21335 14335 21341
rect 14277 21332 14289 21335
rect 13228 21304 14289 21332
rect 13228 21292 13234 21304
rect 14277 21301 14289 21304
rect 14323 21301 14335 21335
rect 14277 21295 14335 21301
rect 15841 21335 15899 21341
rect 15841 21301 15853 21335
rect 15887 21332 15899 21335
rect 16114 21332 16120 21344
rect 15887 21304 16120 21332
rect 15887 21301 15899 21304
rect 15841 21295 15899 21301
rect 16114 21292 16120 21304
rect 16172 21292 16178 21344
rect 16206 21292 16212 21344
rect 16264 21332 16270 21344
rect 18046 21332 18052 21344
rect 16264 21304 18052 21332
rect 16264 21292 16270 21304
rect 18046 21292 18052 21304
rect 18104 21292 18110 21344
rect 19334 21292 19340 21344
rect 19392 21332 19398 21344
rect 19521 21335 19579 21341
rect 19521 21332 19533 21335
rect 19392 21304 19533 21332
rect 19392 21292 19398 21304
rect 19521 21301 19533 21304
rect 19567 21301 19579 21335
rect 20898 21332 20904 21344
rect 20859 21304 20904 21332
rect 19521 21295 19579 21301
rect 20898 21292 20904 21304
rect 20956 21292 20962 21344
rect 29822 21292 29828 21344
rect 29880 21332 29886 21344
rect 33505 21335 33563 21341
rect 33505 21332 33517 21335
rect 29880 21304 33517 21332
rect 29880 21292 29886 21304
rect 33505 21301 33517 21304
rect 33551 21301 33563 21335
rect 33505 21295 33563 21301
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 5537 21131 5595 21137
rect 5537 21097 5549 21131
rect 5583 21128 5595 21131
rect 6914 21128 6920 21140
rect 5583 21100 6920 21128
rect 5583 21097 5595 21100
rect 5537 21091 5595 21097
rect 6914 21088 6920 21100
rect 6972 21088 6978 21140
rect 10870 21088 10876 21140
rect 10928 21128 10934 21140
rect 10965 21131 11023 21137
rect 10965 21128 10977 21131
rect 10928 21100 10977 21128
rect 10928 21088 10934 21100
rect 10965 21097 10977 21100
rect 11011 21097 11023 21131
rect 10965 21091 11023 21097
rect 12066 21088 12072 21140
rect 12124 21128 12130 21140
rect 23658 21128 23664 21140
rect 12124 21100 23664 21128
rect 12124 21088 12130 21100
rect 23658 21088 23664 21100
rect 23716 21088 23722 21140
rect 24578 21088 24584 21140
rect 24636 21128 24642 21140
rect 27341 21131 27399 21137
rect 27341 21128 27353 21131
rect 24636 21100 27353 21128
rect 24636 21088 24642 21100
rect 27341 21097 27353 21100
rect 27387 21097 27399 21131
rect 27341 21091 27399 21097
rect 35989 21131 36047 21137
rect 35989 21097 36001 21131
rect 36035 21128 36047 21131
rect 36078 21128 36084 21140
rect 36035 21100 36084 21128
rect 36035 21097 36047 21100
rect 35989 21091 36047 21097
rect 36078 21088 36084 21100
rect 36136 21088 36142 21140
rect 4614 21020 4620 21072
rect 4672 21060 4678 21072
rect 5721 21063 5779 21069
rect 5721 21060 5733 21063
rect 4672 21032 5733 21060
rect 4672 21020 4678 21032
rect 5721 21029 5733 21032
rect 5767 21029 5779 21063
rect 35342 21060 35348 21072
rect 35303 21032 35348 21060
rect 5721 21023 5779 21029
rect 35342 21020 35348 21032
rect 35400 21020 35406 21072
rect 3053 20995 3111 21001
rect 3053 20961 3065 20995
rect 3099 20992 3111 20995
rect 7098 20992 7104 21004
rect 3099 20964 7104 20992
rect 3099 20961 3111 20964
rect 3053 20955 3111 20961
rect 7098 20952 7104 20964
rect 7156 20952 7162 21004
rect 7466 20992 7472 21004
rect 7392 20964 7472 20992
rect 2774 20884 2780 20936
rect 2832 20924 2838 20936
rect 7392 20933 7420 20964
rect 7466 20952 7472 20964
rect 7524 20992 7530 21004
rect 9858 20992 9864 21004
rect 7524 20964 9168 20992
rect 7524 20952 7530 20964
rect 3237 20927 3295 20933
rect 2832 20896 2877 20924
rect 2832 20884 2838 20896
rect 3237 20893 3249 20927
rect 3283 20893 3295 20927
rect 3237 20887 3295 20893
rect 7377 20927 7435 20933
rect 7377 20893 7389 20927
rect 7423 20893 7435 20927
rect 7558 20924 7564 20936
rect 7519 20896 7564 20924
rect 7377 20887 7435 20893
rect 2958 20816 2964 20868
rect 3016 20856 3022 20868
rect 3252 20856 3280 20887
rect 7558 20884 7564 20896
rect 7616 20884 7622 20936
rect 9140 20933 9168 20964
rect 9600 20964 9864 20992
rect 9600 20933 9628 20964
rect 9858 20952 9864 20964
rect 9916 20952 9922 21004
rect 12253 20995 12311 21001
rect 12253 20961 12265 20995
rect 12299 20992 12311 20995
rect 12434 20992 12440 21004
rect 12299 20964 12440 20992
rect 12299 20961 12311 20964
rect 12253 20955 12311 20961
rect 12434 20952 12440 20964
rect 12492 20992 12498 21004
rect 13446 20992 13452 21004
rect 12492 20964 13452 20992
rect 12492 20952 12498 20964
rect 13446 20952 13452 20964
rect 13504 20952 13510 21004
rect 14550 20952 14556 21004
rect 14608 20992 14614 21004
rect 14918 20992 14924 21004
rect 14608 20964 14924 20992
rect 14608 20952 14614 20964
rect 14918 20952 14924 20964
rect 14976 20952 14982 21004
rect 17405 20995 17463 21001
rect 17405 20961 17417 20995
rect 17451 20992 17463 20995
rect 17586 20992 17592 21004
rect 17451 20964 17592 20992
rect 17451 20961 17463 20964
rect 17405 20955 17463 20961
rect 17586 20952 17592 20964
rect 17644 20952 17650 21004
rect 22554 20992 22560 21004
rect 22515 20964 22560 20992
rect 22554 20952 22560 20964
rect 22612 20952 22618 21004
rect 28902 20952 28908 21004
rect 28960 20992 28966 21004
rect 28960 20964 29960 20992
rect 28960 20952 28966 20964
rect 9125 20927 9183 20933
rect 9125 20893 9137 20927
rect 9171 20893 9183 20927
rect 9125 20887 9183 20893
rect 9585 20927 9643 20933
rect 9585 20893 9597 20927
rect 9631 20893 9643 20927
rect 9766 20924 9772 20936
rect 9727 20896 9772 20924
rect 9585 20887 9643 20893
rect 9766 20884 9772 20896
rect 9824 20884 9830 20936
rect 10873 20927 10931 20933
rect 10873 20893 10885 20927
rect 10919 20893 10931 20927
rect 11974 20924 11980 20936
rect 11935 20896 11980 20924
rect 10873 20887 10931 20893
rect 3016 20828 3280 20856
rect 5353 20859 5411 20865
rect 3016 20816 3022 20828
rect 5353 20825 5365 20859
rect 5399 20856 5411 20859
rect 5442 20856 5448 20868
rect 5399 20828 5448 20856
rect 5399 20825 5411 20828
rect 5353 20819 5411 20825
rect 5442 20816 5448 20828
rect 5500 20816 5506 20868
rect 5569 20859 5627 20865
rect 5569 20825 5581 20859
rect 5615 20856 5627 20859
rect 7006 20856 7012 20868
rect 5615 20828 7012 20856
rect 5615 20825 5627 20828
rect 5569 20819 5627 20825
rect 7006 20816 7012 20828
rect 7064 20856 7070 20868
rect 7469 20859 7527 20865
rect 7469 20856 7481 20859
rect 7064 20828 7481 20856
rect 7064 20816 7070 20828
rect 7469 20825 7481 20828
rect 7515 20856 7527 20859
rect 9030 20856 9036 20868
rect 7515 20828 9036 20856
rect 7515 20825 7527 20828
rect 7469 20819 7527 20825
rect 9030 20816 9036 20828
rect 9088 20816 9094 20868
rect 10888 20856 10916 20887
rect 11974 20884 11980 20896
rect 12032 20924 12038 20936
rect 13906 20924 13912 20936
rect 12032 20896 13912 20924
rect 12032 20884 12038 20896
rect 13906 20884 13912 20896
rect 13964 20884 13970 20936
rect 14369 20927 14427 20933
rect 14369 20893 14381 20927
rect 14415 20924 14427 20927
rect 14458 20924 14464 20936
rect 14415 20896 14464 20924
rect 14415 20893 14427 20896
rect 14369 20887 14427 20893
rect 14458 20884 14464 20896
rect 14516 20884 14522 20936
rect 20809 20927 20867 20933
rect 20809 20893 20821 20927
rect 20855 20924 20867 20927
rect 24762 20924 24768 20936
rect 20855 20896 24768 20924
rect 20855 20893 20867 20896
rect 20809 20887 20867 20893
rect 24762 20884 24768 20896
rect 24820 20924 24826 20936
rect 26053 20927 26111 20933
rect 26053 20924 26065 20927
rect 24820 20896 26065 20924
rect 24820 20884 24826 20896
rect 26053 20893 26065 20896
rect 26099 20893 26111 20927
rect 26053 20887 26111 20893
rect 29733 20927 29791 20933
rect 29733 20893 29745 20927
rect 29779 20924 29791 20927
rect 29822 20924 29828 20936
rect 29779 20896 29828 20924
rect 29779 20893 29791 20896
rect 29733 20887 29791 20893
rect 29822 20884 29828 20896
rect 29880 20884 29886 20936
rect 29932 20933 29960 20964
rect 34790 20952 34796 21004
rect 34848 20992 34854 21004
rect 35437 20995 35495 21001
rect 35437 20992 35449 20995
rect 34848 20964 35449 20992
rect 34848 20952 34854 20964
rect 35437 20961 35449 20964
rect 35483 20961 35495 20995
rect 35437 20955 35495 20961
rect 35802 20952 35808 21004
rect 35860 20992 35866 21004
rect 36630 20992 36636 21004
rect 35860 20964 36308 20992
rect 36591 20964 36636 20992
rect 35860 20952 35866 20964
rect 36170 20933 36176 20936
rect 29917 20927 29975 20933
rect 29917 20893 29929 20927
rect 29963 20893 29975 20927
rect 29917 20887 29975 20893
rect 34885 20927 34943 20933
rect 34885 20893 34897 20927
rect 34931 20893 34943 20927
rect 34885 20887 34943 20893
rect 35069 20927 35127 20933
rect 35069 20893 35081 20927
rect 35115 20924 35127 20927
rect 36153 20927 36176 20933
rect 36153 20924 36165 20927
rect 35115 20896 36165 20924
rect 35115 20893 35127 20896
rect 35069 20887 35127 20893
rect 36153 20893 36165 20896
rect 36153 20887 36176 20893
rect 9646 20828 10916 20856
rect 15657 20859 15715 20865
rect 5258 20748 5264 20800
rect 5316 20788 5322 20800
rect 9398 20788 9404 20800
rect 5316 20760 9404 20788
rect 5316 20748 5322 20760
rect 9398 20748 9404 20760
rect 9456 20788 9462 20800
rect 9646 20788 9674 20828
rect 15657 20825 15669 20859
rect 15703 20856 15715 20859
rect 16482 20856 16488 20868
rect 15703 20828 16488 20856
rect 15703 20825 15715 20828
rect 15657 20819 15715 20825
rect 16482 20816 16488 20828
rect 16540 20816 16546 20868
rect 34900 20856 34928 20887
rect 36170 20884 36176 20887
rect 36228 20884 36234 20936
rect 36280 20933 36308 20964
rect 36630 20952 36636 20964
rect 36688 20952 36694 21004
rect 36265 20927 36323 20933
rect 36265 20893 36277 20927
rect 36311 20893 36323 20927
rect 36265 20887 36323 20893
rect 35894 20856 35900 20868
rect 34900 20828 35900 20856
rect 35894 20816 35900 20828
rect 35952 20816 35958 20868
rect 36541 20859 36599 20865
rect 36541 20825 36553 20859
rect 36587 20856 36599 20859
rect 36722 20856 36728 20868
rect 36587 20828 36728 20856
rect 36587 20825 36599 20828
rect 36541 20819 36599 20825
rect 36722 20816 36728 20828
rect 36780 20816 36786 20868
rect 10410 20788 10416 20800
rect 9456 20760 9674 20788
rect 10371 20760 10416 20788
rect 9456 20748 9462 20760
rect 10410 20748 10416 20760
rect 10468 20748 10474 20800
rect 28994 20748 29000 20800
rect 29052 20788 29058 20800
rect 29825 20791 29883 20797
rect 29825 20788 29837 20791
rect 29052 20760 29837 20788
rect 29052 20748 29058 20760
rect 29825 20757 29837 20760
rect 29871 20757 29883 20791
rect 29825 20751 29883 20757
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 2774 20544 2780 20596
rect 2832 20584 2838 20596
rect 2832 20556 2877 20584
rect 2832 20544 2838 20556
rect 6914 20544 6920 20596
rect 6972 20593 6978 20596
rect 6972 20584 6984 20593
rect 9217 20587 9275 20593
rect 6972 20556 7017 20584
rect 6972 20547 6984 20556
rect 9217 20553 9229 20587
rect 9263 20584 9275 20587
rect 12066 20584 12072 20596
rect 9263 20556 12072 20584
rect 9263 20553 9275 20556
rect 9217 20547 9275 20553
rect 6972 20544 6978 20547
rect 12066 20544 12072 20556
rect 12124 20544 12130 20596
rect 16853 20587 16911 20593
rect 16853 20553 16865 20587
rect 16899 20584 16911 20587
rect 16942 20584 16948 20596
rect 16899 20556 16948 20584
rect 16899 20553 16911 20556
rect 16853 20547 16911 20553
rect 16942 20544 16948 20556
rect 17000 20544 17006 20596
rect 17221 20587 17279 20593
rect 17221 20553 17233 20587
rect 17267 20584 17279 20587
rect 18322 20584 18328 20596
rect 17267 20556 18328 20584
rect 17267 20553 17279 20556
rect 17221 20547 17279 20553
rect 18322 20544 18328 20556
rect 18380 20544 18386 20596
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 19521 20587 19579 20593
rect 19521 20584 19533 20587
rect 19484 20556 19533 20584
rect 19484 20544 19490 20556
rect 19521 20553 19533 20556
rect 19567 20553 19579 20587
rect 19521 20547 19579 20553
rect 20990 20544 20996 20596
rect 21048 20584 21054 20596
rect 21085 20587 21143 20593
rect 21085 20584 21097 20587
rect 21048 20556 21097 20584
rect 21048 20544 21054 20556
rect 21085 20553 21097 20556
rect 21131 20553 21143 20587
rect 21085 20547 21143 20553
rect 6549 20519 6607 20525
rect 6549 20485 6561 20519
rect 6595 20516 6607 20519
rect 7558 20516 7564 20528
rect 6595 20488 7564 20516
rect 6595 20485 6607 20488
rect 6549 20479 6607 20485
rect 7558 20476 7564 20488
rect 7616 20476 7622 20528
rect 12989 20519 13047 20525
rect 12989 20485 13001 20519
rect 13035 20516 13047 20519
rect 18233 20519 18291 20525
rect 18233 20516 18245 20519
rect 13035 20488 18245 20516
rect 13035 20485 13047 20488
rect 12989 20479 13047 20485
rect 18233 20485 18245 20488
rect 18279 20516 18291 20519
rect 19334 20516 19340 20528
rect 18279 20488 19340 20516
rect 18279 20485 18291 20488
rect 18233 20479 18291 20485
rect 19334 20476 19340 20488
rect 19392 20476 19398 20528
rect 20806 20516 20812 20528
rect 20719 20488 20812 20516
rect 20806 20476 20812 20488
rect 20864 20516 20870 20528
rect 21266 20516 21272 20528
rect 20864 20488 21272 20516
rect 20864 20476 20870 20488
rect 21266 20476 21272 20488
rect 21324 20476 21330 20528
rect 21634 20476 21640 20528
rect 21692 20516 21698 20528
rect 26237 20519 26295 20525
rect 26237 20516 26249 20519
rect 21692 20488 26249 20516
rect 21692 20476 21698 20488
rect 26237 20485 26249 20488
rect 26283 20516 26295 20519
rect 26602 20516 26608 20528
rect 26283 20488 26608 20516
rect 26283 20485 26295 20488
rect 26237 20479 26295 20485
rect 26602 20476 26608 20488
rect 26660 20476 26666 20528
rect 29546 20476 29552 20528
rect 29604 20516 29610 20528
rect 31754 20516 31760 20528
rect 29604 20488 30880 20516
rect 29604 20476 29610 20488
rect 2685 20451 2743 20457
rect 2685 20417 2697 20451
rect 2731 20448 2743 20451
rect 2866 20448 2872 20460
rect 2731 20420 2872 20448
rect 2731 20417 2743 20420
rect 2685 20411 2743 20417
rect 2866 20408 2872 20420
rect 2924 20408 2930 20460
rect 4706 20408 4712 20460
rect 4764 20448 4770 20460
rect 7193 20451 7251 20457
rect 7193 20448 7205 20451
rect 4764 20420 7205 20448
rect 4764 20408 4770 20420
rect 7193 20417 7205 20420
rect 7239 20417 7251 20451
rect 7193 20411 7251 20417
rect 7374 20408 7380 20460
rect 7432 20448 7438 20460
rect 7653 20451 7711 20457
rect 7653 20448 7665 20451
rect 7432 20420 7665 20448
rect 7432 20408 7438 20420
rect 7653 20417 7665 20420
rect 7699 20417 7711 20451
rect 9030 20448 9036 20460
rect 8991 20420 9036 20448
rect 7653 20411 7711 20417
rect 9030 20408 9036 20420
rect 9088 20408 9094 20460
rect 9674 20448 9680 20460
rect 9508 20420 9680 20448
rect 9508 20389 9536 20420
rect 9674 20408 9680 20420
rect 9732 20408 9738 20460
rect 11885 20451 11943 20457
rect 11885 20417 11897 20451
rect 11931 20448 11943 20451
rect 12434 20448 12440 20460
rect 11931 20420 12440 20448
rect 11931 20417 11943 20420
rect 11885 20411 11943 20417
rect 12434 20408 12440 20420
rect 12492 20408 12498 20460
rect 14826 20408 14832 20460
rect 14884 20448 14890 20460
rect 15381 20451 15439 20457
rect 15381 20448 15393 20451
rect 14884 20420 15393 20448
rect 14884 20408 14890 20420
rect 15381 20417 15393 20420
rect 15427 20417 15439 20451
rect 15562 20448 15568 20460
rect 15523 20420 15568 20448
rect 15381 20411 15439 20417
rect 15562 20408 15568 20420
rect 15620 20408 15626 20460
rect 15654 20408 15660 20460
rect 15712 20448 15718 20460
rect 15712 20420 16988 20448
rect 15712 20408 15718 20420
rect 9493 20383 9551 20389
rect 9493 20349 9505 20383
rect 9539 20349 9551 20383
rect 9493 20343 9551 20349
rect 9585 20383 9643 20389
rect 9585 20349 9597 20383
rect 9631 20349 9643 20383
rect 9585 20343 9643 20349
rect 12161 20383 12219 20389
rect 12161 20349 12173 20383
rect 12207 20380 12219 20383
rect 12526 20380 12532 20392
rect 12207 20352 12532 20380
rect 12207 20349 12219 20352
rect 12161 20343 12219 20349
rect 8202 20272 8208 20324
rect 8260 20312 8266 20324
rect 9600 20312 9628 20343
rect 12526 20340 12532 20352
rect 12584 20380 12590 20392
rect 13630 20380 13636 20392
rect 12584 20352 13636 20380
rect 12584 20340 12590 20352
rect 13630 20340 13636 20352
rect 13688 20340 13694 20392
rect 14737 20383 14795 20389
rect 14737 20349 14749 20383
rect 14783 20380 14795 20383
rect 16298 20380 16304 20392
rect 14783 20352 16304 20380
rect 14783 20349 14795 20352
rect 14737 20343 14795 20349
rect 16298 20340 16304 20352
rect 16356 20340 16362 20392
rect 16960 20380 16988 20420
rect 17034 20408 17040 20460
rect 17092 20448 17098 20460
rect 17313 20451 17371 20457
rect 17092 20420 17137 20448
rect 17092 20408 17098 20420
rect 17313 20417 17325 20451
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 17328 20380 17356 20411
rect 20162 20408 20168 20460
rect 20220 20448 20226 20460
rect 20441 20451 20499 20457
rect 20441 20448 20453 20451
rect 20220 20420 20453 20448
rect 20220 20408 20226 20420
rect 20441 20417 20453 20420
rect 20487 20417 20499 20451
rect 20441 20411 20499 20417
rect 20530 20408 20536 20460
rect 20588 20448 20594 20460
rect 20714 20448 20720 20460
rect 20588 20420 20633 20448
rect 20675 20420 20720 20448
rect 20588 20408 20594 20420
rect 20714 20408 20720 20420
rect 20772 20408 20778 20460
rect 20906 20451 20964 20457
rect 20906 20448 20918 20451
rect 20824 20420 20918 20448
rect 20824 20380 20852 20420
rect 20906 20417 20918 20420
rect 20952 20448 20964 20451
rect 21450 20448 21456 20460
rect 20952 20420 21456 20448
rect 20952 20417 20964 20420
rect 20906 20411 20964 20417
rect 21450 20408 21456 20420
rect 21508 20408 21514 20460
rect 23382 20408 23388 20460
rect 23440 20448 23446 20460
rect 23753 20451 23811 20457
rect 23753 20448 23765 20451
rect 23440 20420 23765 20448
rect 23440 20408 23446 20420
rect 16960 20352 17356 20380
rect 17972 20352 20852 20380
rect 8260 20284 9628 20312
rect 8260 20272 8266 20284
rect 16850 20272 16856 20324
rect 16908 20312 16914 20324
rect 17972 20312 18000 20352
rect 16908 20284 18000 20312
rect 16908 20272 16914 20284
rect 6917 20247 6975 20253
rect 6917 20213 6929 20247
rect 6963 20244 6975 20247
rect 7466 20244 7472 20256
rect 6963 20216 7472 20244
rect 6963 20213 6975 20216
rect 6917 20207 6975 20213
rect 7466 20204 7472 20216
rect 7524 20204 7530 20256
rect 7742 20244 7748 20256
rect 7703 20216 7748 20244
rect 7742 20204 7748 20216
rect 7800 20204 7806 20256
rect 13814 20204 13820 20256
rect 13872 20244 13878 20256
rect 15197 20247 15255 20253
rect 15197 20244 15209 20247
rect 13872 20216 15209 20244
rect 13872 20204 13878 20216
rect 15197 20213 15209 20216
rect 15243 20213 15255 20247
rect 15197 20207 15255 20213
rect 18046 20204 18052 20256
rect 18104 20244 18110 20256
rect 23566 20244 23572 20256
rect 18104 20216 23572 20244
rect 18104 20204 18110 20216
rect 23566 20204 23572 20216
rect 23624 20204 23630 20256
rect 23676 20244 23704 20420
rect 23753 20417 23765 20420
rect 23799 20417 23811 20451
rect 23753 20411 23811 20417
rect 25958 20408 25964 20460
rect 26016 20448 26022 20460
rect 26053 20451 26111 20457
rect 26053 20448 26065 20451
rect 26016 20420 26065 20448
rect 26016 20408 26022 20420
rect 26053 20417 26065 20420
rect 26099 20417 26111 20451
rect 26326 20448 26332 20460
rect 26287 20420 26332 20448
rect 26053 20411 26111 20417
rect 26326 20408 26332 20420
rect 26384 20448 26390 20460
rect 27614 20448 27620 20460
rect 26384 20420 27620 20448
rect 26384 20408 26390 20420
rect 27614 20408 27620 20420
rect 27672 20408 27678 20460
rect 24026 20380 24032 20392
rect 23939 20352 24032 20380
rect 24026 20340 24032 20352
rect 24084 20380 24090 20392
rect 26344 20380 26372 20408
rect 24084 20352 26372 20380
rect 24084 20340 24090 20352
rect 23750 20272 23756 20324
rect 23808 20312 23814 20324
rect 24044 20312 24072 20340
rect 29546 20312 29552 20324
rect 23808 20284 24072 20312
rect 25700 20284 29552 20312
rect 23808 20272 23814 20284
rect 25700 20244 25728 20284
rect 29546 20272 29552 20284
rect 29604 20272 29610 20324
rect 30484 20312 30512 20488
rect 30561 20451 30619 20457
rect 30561 20417 30573 20451
rect 30607 20417 30619 20451
rect 30742 20448 30748 20460
rect 30703 20420 30748 20448
rect 30561 20411 30619 20417
rect 30576 20380 30604 20411
rect 30742 20408 30748 20420
rect 30800 20408 30806 20460
rect 30852 20457 30880 20488
rect 31128 20488 31760 20516
rect 30837 20451 30895 20457
rect 30837 20417 30849 20451
rect 30883 20417 30895 20451
rect 30837 20411 30895 20417
rect 31128 20392 31156 20488
rect 31754 20476 31760 20488
rect 31812 20476 31818 20528
rect 31110 20380 31116 20392
rect 30576 20352 31116 20380
rect 31110 20340 31116 20352
rect 31168 20340 31174 20392
rect 32306 20380 32312 20392
rect 31726 20352 32312 20380
rect 31726 20312 31754 20352
rect 32306 20340 32312 20352
rect 32364 20340 32370 20392
rect 38102 20380 38108 20392
rect 38063 20352 38108 20380
rect 38102 20340 38108 20352
rect 38160 20340 38166 20392
rect 30484 20284 31754 20312
rect 25866 20244 25872 20256
rect 23676 20216 25728 20244
rect 25827 20216 25872 20244
rect 25866 20204 25872 20216
rect 25924 20204 25930 20256
rect 30006 20204 30012 20256
rect 30064 20244 30070 20256
rect 30377 20247 30435 20253
rect 30377 20244 30389 20247
rect 30064 20216 30389 20244
rect 30064 20204 30070 20216
rect 30377 20213 30389 20216
rect 30423 20213 30435 20247
rect 30377 20207 30435 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 17218 20040 17224 20052
rect 14660 20012 16804 20040
rect 17179 20012 17224 20040
rect 13725 19975 13783 19981
rect 13725 19941 13737 19975
rect 13771 19972 13783 19975
rect 14660 19972 14688 20012
rect 13771 19944 14688 19972
rect 16776 19972 16804 20012
rect 17218 20000 17224 20012
rect 17276 20000 17282 20052
rect 20530 20040 20536 20052
rect 17328 20012 20536 20040
rect 17328 19972 17356 20012
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 20806 20040 20812 20052
rect 20767 20012 20812 20040
rect 20806 20000 20812 20012
rect 20864 20000 20870 20052
rect 21913 20043 21971 20049
rect 21913 20009 21925 20043
rect 21959 20040 21971 20043
rect 22002 20040 22008 20052
rect 21959 20012 22008 20040
rect 21959 20009 21971 20012
rect 21913 20003 21971 20009
rect 22002 20000 22008 20012
rect 22060 20000 22066 20052
rect 24854 20040 24860 20052
rect 22112 20012 24860 20040
rect 16776 19944 17356 19972
rect 13771 19941 13783 19944
rect 13725 19935 13783 19941
rect 12345 19839 12403 19845
rect 12345 19805 12357 19839
rect 12391 19836 12403 19839
rect 12894 19836 12900 19848
rect 12391 19808 12900 19836
rect 12391 19805 12403 19808
rect 12345 19799 12403 19805
rect 12894 19796 12900 19808
rect 12952 19836 12958 19848
rect 13170 19836 13176 19848
rect 12952 19808 13176 19836
rect 12952 19796 12958 19808
rect 13170 19796 13176 19808
rect 13228 19796 13234 19848
rect 14461 19839 14519 19845
rect 14461 19805 14473 19839
rect 14507 19836 14519 19839
rect 14550 19836 14556 19848
rect 14507 19808 14556 19836
rect 14507 19805 14519 19808
rect 14461 19799 14519 19805
rect 14550 19796 14556 19808
rect 14608 19796 14614 19848
rect 14660 19845 14688 19944
rect 19426 19904 19432 19916
rect 19387 19876 19432 19904
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 22112 19904 22140 20012
rect 24854 20000 24860 20012
rect 24912 20040 24918 20052
rect 27525 20043 27583 20049
rect 24912 20012 25176 20040
rect 24912 20000 24918 20012
rect 22186 19932 22192 19984
rect 22244 19972 22250 19984
rect 22244 19944 25084 19972
rect 22244 19932 22250 19944
rect 22066 19876 22140 19904
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19805 14703 19839
rect 14645 19799 14703 19805
rect 14737 19839 14795 19845
rect 14737 19805 14749 19839
rect 14783 19836 14795 19839
rect 15654 19836 15660 19848
rect 14783 19808 15660 19836
rect 14783 19805 14795 19808
rect 14737 19799 14795 19805
rect 12612 19771 12670 19777
rect 12612 19737 12624 19771
rect 12658 19768 12670 19771
rect 14277 19771 14335 19777
rect 14277 19768 14289 19771
rect 12658 19740 14289 19768
rect 12658 19737 12670 19740
rect 12612 19731 12670 19737
rect 14277 19737 14289 19740
rect 14323 19737 14335 19771
rect 14277 19731 14335 19737
rect 13630 19660 13636 19712
rect 13688 19700 13694 19712
rect 14752 19700 14780 19799
rect 15654 19796 15660 19808
rect 15712 19796 15718 19848
rect 16114 19845 16120 19848
rect 15841 19839 15899 19845
rect 15841 19805 15853 19839
rect 15887 19805 15899 19839
rect 16108 19836 16120 19845
rect 16075 19808 16120 19836
rect 15841 19799 15899 19805
rect 16108 19799 16120 19808
rect 13688 19672 14780 19700
rect 15856 19700 15884 19799
rect 16114 19796 16120 19799
rect 16172 19796 16178 19848
rect 19696 19839 19754 19845
rect 19696 19805 19708 19839
rect 19742 19836 19754 19839
rect 20898 19836 20904 19848
rect 19742 19808 20904 19836
rect 19742 19805 19754 19808
rect 19696 19799 19754 19805
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 21266 19836 21272 19848
rect 21227 19808 21272 19836
rect 21266 19796 21272 19808
rect 21324 19796 21330 19848
rect 21358 19796 21364 19848
rect 21416 19836 21422 19848
rect 21634 19836 21640 19848
rect 21416 19808 21461 19836
rect 21595 19808 21640 19836
rect 21416 19796 21422 19808
rect 21634 19796 21640 19808
rect 21692 19796 21698 19848
rect 21775 19839 21833 19845
rect 21775 19805 21787 19839
rect 21821 19836 21833 19839
rect 22066 19836 22094 19876
rect 22462 19864 22468 19916
rect 22520 19904 22526 19916
rect 22520 19876 24808 19904
rect 22520 19864 22526 19876
rect 23658 19836 23664 19848
rect 21821 19808 22094 19836
rect 23619 19808 23664 19836
rect 21821 19805 21833 19808
rect 21775 19799 21833 19805
rect 23658 19796 23664 19808
rect 23716 19796 23722 19848
rect 24780 19845 24808 19876
rect 25056 19845 25084 19944
rect 24765 19839 24823 19845
rect 24765 19805 24777 19839
rect 24811 19805 24823 19839
rect 24765 19799 24823 19805
rect 24858 19839 24916 19845
rect 24858 19805 24870 19839
rect 24904 19805 24916 19839
rect 24858 19799 24916 19805
rect 25041 19839 25099 19845
rect 25041 19805 25053 19839
rect 25087 19805 25099 19839
rect 25148 19836 25176 20012
rect 27525 20009 27537 20043
rect 27571 20040 27583 20043
rect 28166 20040 28172 20052
rect 27571 20012 28172 20040
rect 27571 20009 27583 20012
rect 27525 20003 27583 20009
rect 28166 20000 28172 20012
rect 28224 20000 28230 20052
rect 28350 20040 28356 20052
rect 28311 20012 28356 20040
rect 28350 20000 28356 20012
rect 28408 20000 28414 20052
rect 28626 20040 28632 20052
rect 28587 20012 28632 20040
rect 28626 20000 28632 20012
rect 28684 20000 28690 20052
rect 30742 20000 30748 20052
rect 30800 20040 30806 20052
rect 31113 20043 31171 20049
rect 31113 20040 31125 20043
rect 30800 20012 31125 20040
rect 30800 20000 30806 20012
rect 31113 20009 31125 20012
rect 31159 20040 31171 20043
rect 33318 20040 33324 20052
rect 31159 20012 33324 20040
rect 31159 20009 31171 20012
rect 31113 20003 31171 20009
rect 33318 20000 33324 20012
rect 33376 20000 33382 20052
rect 34790 20000 34796 20052
rect 34848 20040 34854 20052
rect 34977 20043 35035 20049
rect 34977 20040 34989 20043
rect 34848 20012 34989 20040
rect 34848 20000 34854 20012
rect 34977 20009 34989 20012
rect 35023 20009 35035 20043
rect 34977 20003 35035 20009
rect 36262 20000 36268 20052
rect 36320 20040 36326 20052
rect 36725 20043 36783 20049
rect 36725 20040 36737 20043
rect 36320 20012 36737 20040
rect 36320 20000 36326 20012
rect 36725 20009 36737 20012
rect 36771 20009 36783 20043
rect 36725 20003 36783 20009
rect 30006 19904 30012 19916
rect 29967 19876 30012 19904
rect 30006 19864 30012 19876
rect 30064 19864 30070 19916
rect 33318 19864 33324 19916
rect 33376 19904 33382 19916
rect 36081 19907 36139 19913
rect 33376 19876 35112 19904
rect 33376 19864 33382 19876
rect 25230 19839 25288 19845
rect 25230 19836 25242 19839
rect 25148 19808 25242 19836
rect 25041 19799 25099 19805
rect 25230 19805 25242 19808
rect 25276 19805 25288 19839
rect 26050 19836 26056 19848
rect 26011 19808 26056 19836
rect 25230 19799 25288 19805
rect 17034 19728 17040 19780
rect 17092 19768 17098 19780
rect 21174 19768 21180 19780
rect 17092 19740 21180 19768
rect 17092 19728 17098 19740
rect 21174 19728 21180 19740
rect 21232 19728 21238 19780
rect 21450 19728 21456 19780
rect 21508 19768 21514 19780
rect 21545 19771 21603 19777
rect 21545 19768 21557 19771
rect 21508 19740 21557 19768
rect 21508 19728 21514 19740
rect 21545 19737 21557 19740
rect 21591 19737 21603 19771
rect 21545 19731 21603 19737
rect 23842 19728 23848 19780
rect 23900 19768 23906 19780
rect 24872 19768 24900 19799
rect 26050 19796 26056 19808
rect 26108 19796 26114 19848
rect 28258 19836 28264 19848
rect 28219 19808 28264 19836
rect 28258 19796 28264 19808
rect 28316 19796 28322 19848
rect 28445 19839 28503 19845
rect 28445 19805 28457 19839
rect 28491 19836 28503 19839
rect 28994 19836 29000 19848
rect 28491 19808 29000 19836
rect 28491 19805 28503 19808
rect 28445 19799 28503 19805
rect 28994 19796 29000 19808
rect 29052 19796 29058 19848
rect 29638 19796 29644 19848
rect 29696 19836 29702 19848
rect 29733 19839 29791 19845
rect 29733 19836 29745 19839
rect 29696 19808 29745 19836
rect 29696 19796 29702 19808
rect 29733 19805 29745 19808
rect 29779 19805 29791 19839
rect 29733 19799 29791 19805
rect 32033 19839 32091 19845
rect 32033 19805 32045 19839
rect 32079 19805 32091 19839
rect 32306 19836 32312 19848
rect 32267 19808 32312 19836
rect 32033 19799 32091 19805
rect 23900 19740 24900 19768
rect 25133 19771 25191 19777
rect 23900 19728 23906 19740
rect 25133 19737 25145 19771
rect 25179 19768 25191 19771
rect 26878 19768 26884 19780
rect 25179 19740 26884 19768
rect 25179 19737 25191 19740
rect 25133 19731 25191 19737
rect 26878 19728 26884 19740
rect 26936 19728 26942 19780
rect 32048 19768 32076 19799
rect 32306 19796 32312 19808
rect 32364 19796 32370 19848
rect 35084 19845 35112 19876
rect 36081 19873 36093 19907
rect 36127 19904 36139 19907
rect 36170 19904 36176 19916
rect 36127 19876 36176 19904
rect 36127 19873 36139 19876
rect 36081 19867 36139 19873
rect 36170 19864 36176 19876
rect 36228 19864 36234 19916
rect 34977 19839 35035 19845
rect 34977 19805 34989 19839
rect 35023 19805 35035 19839
rect 34977 19799 35035 19805
rect 35069 19839 35127 19845
rect 35069 19805 35081 19839
rect 35115 19805 35127 19839
rect 35069 19799 35127 19805
rect 32490 19768 32496 19780
rect 32048 19740 32496 19768
rect 32490 19728 32496 19740
rect 32548 19728 32554 19780
rect 34992 19768 35020 19799
rect 35342 19796 35348 19848
rect 35400 19836 35406 19848
rect 35713 19839 35771 19845
rect 35713 19836 35725 19839
rect 35400 19808 35725 19836
rect 35400 19796 35406 19808
rect 35713 19805 35725 19808
rect 35759 19805 35771 19839
rect 35986 19836 35992 19848
rect 35947 19808 35992 19836
rect 35713 19799 35771 19805
rect 35986 19796 35992 19808
rect 36044 19796 36050 19848
rect 36538 19836 36544 19848
rect 36499 19808 36544 19836
rect 36538 19796 36544 19808
rect 36596 19796 36602 19848
rect 36695 19839 36753 19845
rect 36695 19805 36707 19839
rect 36741 19836 36753 19839
rect 36906 19836 36912 19848
rect 36741 19808 36912 19836
rect 36741 19805 36753 19808
rect 36695 19799 36753 19805
rect 36906 19796 36912 19808
rect 36964 19796 36970 19848
rect 36446 19768 36452 19780
rect 34992 19740 36452 19768
rect 36446 19728 36452 19740
rect 36504 19728 36510 19780
rect 16298 19700 16304 19712
rect 15856 19672 16304 19700
rect 13688 19660 13694 19672
rect 16298 19660 16304 19672
rect 16356 19660 16362 19712
rect 22922 19660 22928 19712
rect 22980 19700 22986 19712
rect 23382 19700 23388 19712
rect 22980 19672 23388 19700
rect 22980 19660 22986 19672
rect 23382 19660 23388 19672
rect 23440 19700 23446 19712
rect 23753 19703 23811 19709
rect 23753 19700 23765 19703
rect 23440 19672 23765 19700
rect 23440 19660 23446 19672
rect 23753 19669 23765 19672
rect 23799 19669 23811 19703
rect 23753 19663 23811 19669
rect 25409 19703 25467 19709
rect 25409 19669 25421 19703
rect 25455 19700 25467 19703
rect 27522 19700 27528 19712
rect 25455 19672 27528 19700
rect 25455 19669 25467 19672
rect 25409 19663 25467 19669
rect 27522 19660 27528 19672
rect 27580 19660 27586 19712
rect 31202 19660 31208 19712
rect 31260 19700 31266 19712
rect 31849 19703 31907 19709
rect 31849 19700 31861 19703
rect 31260 19672 31861 19700
rect 31260 19660 31266 19672
rect 31849 19669 31861 19672
rect 31895 19669 31907 19703
rect 32214 19700 32220 19712
rect 32175 19672 32220 19700
rect 31849 19663 31907 19669
rect 32214 19660 32220 19672
rect 32272 19660 32278 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 7098 19456 7104 19508
rect 7156 19496 7162 19508
rect 7653 19499 7711 19505
rect 7653 19496 7665 19499
rect 7156 19468 7665 19496
rect 7156 19456 7162 19468
rect 7653 19465 7665 19468
rect 7699 19465 7711 19499
rect 13998 19496 14004 19508
rect 13959 19468 14004 19496
rect 7653 19459 7711 19465
rect 13998 19456 14004 19468
rect 14056 19456 14062 19508
rect 18325 19499 18383 19505
rect 18325 19465 18337 19499
rect 18371 19496 18383 19499
rect 22094 19496 22100 19508
rect 18371 19468 22100 19496
rect 18371 19465 18383 19468
rect 18325 19459 18383 19465
rect 22094 19456 22100 19468
rect 22152 19456 22158 19508
rect 23842 19496 23848 19508
rect 23803 19468 23848 19496
rect 23842 19456 23848 19468
rect 23900 19456 23906 19508
rect 26602 19496 26608 19508
rect 26563 19468 26608 19496
rect 26602 19456 26608 19468
rect 26660 19456 26666 19508
rect 35894 19456 35900 19508
rect 35952 19496 35958 19508
rect 36633 19499 36691 19505
rect 36633 19496 36645 19499
rect 35952 19468 36645 19496
rect 35952 19456 35958 19468
rect 36633 19465 36645 19468
rect 36679 19465 36691 19499
rect 36633 19459 36691 19465
rect 7469 19431 7527 19437
rect 7469 19397 7481 19431
rect 7515 19397 7527 19431
rect 7469 19391 7527 19397
rect 25492 19431 25550 19437
rect 25492 19397 25504 19431
rect 25538 19428 25550 19431
rect 25866 19428 25872 19440
rect 25538 19400 25872 19428
rect 25538 19397 25550 19400
rect 25492 19391 25550 19397
rect 4798 19360 4804 19372
rect 4759 19332 4804 19360
rect 4798 19320 4804 19332
rect 4856 19320 4862 19372
rect 5074 19360 5080 19372
rect 5035 19332 5080 19360
rect 5074 19320 5080 19332
rect 5132 19320 5138 19372
rect 6730 19360 6736 19372
rect 6643 19332 6736 19360
rect 6730 19320 6736 19332
rect 6788 19360 6794 19372
rect 6914 19360 6920 19372
rect 6788 19332 6920 19360
rect 6788 19320 6794 19332
rect 6914 19320 6920 19332
rect 6972 19360 6978 19372
rect 7484 19360 7512 19391
rect 25866 19388 25872 19400
rect 25924 19388 25930 19440
rect 26878 19388 26884 19440
rect 26936 19428 26942 19440
rect 27525 19431 27583 19437
rect 27525 19428 27537 19431
rect 26936 19400 27537 19428
rect 26936 19388 26942 19400
rect 27525 19397 27537 19400
rect 27571 19397 27583 19431
rect 27525 19391 27583 19397
rect 31297 19431 31355 19437
rect 31297 19397 31309 19431
rect 31343 19428 31355 19431
rect 32214 19428 32220 19440
rect 31343 19400 32220 19428
rect 31343 19397 31355 19400
rect 31297 19391 31355 19397
rect 32214 19388 32220 19400
rect 32272 19388 32278 19440
rect 35544 19400 36216 19428
rect 6972 19332 7512 19360
rect 7929 19363 7987 19369
rect 6972 19320 6978 19332
rect 7929 19329 7941 19363
rect 7975 19360 7987 19363
rect 8938 19360 8944 19372
rect 7975 19332 8944 19360
rect 7975 19329 7987 19332
rect 7929 19323 7987 19329
rect 8938 19320 8944 19332
rect 8996 19320 9002 19372
rect 12713 19363 12771 19369
rect 12713 19329 12725 19363
rect 12759 19360 12771 19363
rect 13446 19360 13452 19372
rect 12759 19332 13452 19360
rect 12759 19329 12771 19332
rect 12713 19323 12771 19329
rect 13446 19320 13452 19332
rect 13504 19320 13510 19372
rect 14550 19320 14556 19372
rect 14608 19360 14614 19372
rect 15378 19360 15384 19372
rect 14608 19332 15384 19360
rect 14608 19320 14614 19332
rect 15378 19320 15384 19332
rect 15436 19320 15442 19372
rect 17957 19363 18015 19369
rect 17957 19329 17969 19363
rect 18003 19360 18015 19363
rect 18782 19360 18788 19372
rect 18003 19332 18788 19360
rect 18003 19329 18015 19332
rect 17957 19323 18015 19329
rect 18782 19320 18788 19332
rect 18840 19320 18846 19372
rect 22002 19320 22008 19372
rect 22060 19360 22066 19372
rect 22465 19363 22523 19369
rect 22465 19360 22477 19363
rect 22060 19332 22477 19360
rect 22060 19320 22066 19332
rect 22465 19329 22477 19332
rect 22511 19329 22523 19363
rect 22465 19323 22523 19329
rect 22732 19363 22790 19369
rect 22732 19329 22744 19363
rect 22778 19360 22790 19363
rect 23198 19360 23204 19372
rect 22778 19332 23204 19360
rect 22778 19329 22790 19332
rect 22732 19323 22790 19329
rect 23198 19320 23204 19332
rect 23256 19320 23262 19372
rect 27341 19363 27399 19369
rect 27341 19360 27353 19363
rect 26252 19332 27353 19360
rect 7006 19292 7012 19304
rect 6967 19264 7012 19292
rect 7006 19252 7012 19264
rect 7064 19252 7070 19304
rect 15194 19252 15200 19304
rect 15252 19292 15258 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 15252 19264 18061 19292
rect 15252 19252 15258 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 25222 19292 25228 19304
rect 25183 19264 25228 19292
rect 18049 19255 18107 19261
rect 25222 19252 25228 19264
rect 25280 19252 25286 19304
rect 4890 19156 4896 19168
rect 4851 19128 4896 19156
rect 4890 19116 4896 19128
rect 4948 19116 4954 19168
rect 6086 19116 6092 19168
rect 6144 19156 6150 19168
rect 6549 19159 6607 19165
rect 6549 19156 6561 19159
rect 6144 19128 6561 19156
rect 6144 19116 6150 19128
rect 6549 19125 6561 19128
rect 6595 19125 6607 19159
rect 6549 19119 6607 19125
rect 6917 19159 6975 19165
rect 6917 19125 6929 19159
rect 6963 19156 6975 19159
rect 7653 19159 7711 19165
rect 7653 19156 7665 19159
rect 6963 19128 7665 19156
rect 6963 19125 6975 19128
rect 6917 19119 6975 19125
rect 7653 19125 7665 19128
rect 7699 19156 7711 19159
rect 7742 19156 7748 19168
rect 7699 19128 7748 19156
rect 7699 19125 7711 19128
rect 7653 19119 7711 19125
rect 7742 19116 7748 19128
rect 7800 19116 7806 19168
rect 18138 19156 18144 19168
rect 18099 19128 18144 19156
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 25866 19116 25872 19168
rect 25924 19156 25930 19168
rect 26252 19156 26280 19332
rect 27341 19329 27353 19332
rect 27387 19329 27399 19363
rect 27614 19360 27620 19372
rect 27575 19332 27620 19360
rect 27341 19323 27399 19329
rect 27614 19320 27620 19332
rect 27672 19320 27678 19372
rect 35544 19369 35572 19400
rect 36188 19372 36216 19400
rect 35529 19363 35587 19369
rect 35529 19329 35541 19363
rect 35575 19329 35587 19363
rect 35529 19323 35587 19329
rect 35713 19363 35771 19369
rect 35713 19329 35725 19363
rect 35759 19360 35771 19363
rect 35759 19332 36124 19360
rect 35759 19329 35771 19332
rect 35713 19323 35771 19329
rect 36096 19304 36124 19332
rect 36170 19320 36176 19372
rect 36228 19360 36234 19372
rect 36449 19363 36507 19369
rect 36228 19332 36273 19360
rect 36228 19320 36234 19332
rect 36449 19329 36461 19363
rect 36495 19360 36507 19363
rect 36906 19360 36912 19372
rect 36495 19332 36912 19360
rect 36495 19329 36507 19332
rect 36449 19323 36507 19329
rect 36906 19320 36912 19332
rect 36964 19320 36970 19372
rect 29638 19292 29644 19304
rect 29599 19264 29644 19292
rect 29638 19252 29644 19264
rect 29696 19252 29702 19304
rect 29917 19295 29975 19301
rect 29917 19261 29929 19295
rect 29963 19292 29975 19295
rect 31202 19292 31208 19304
rect 29963 19264 31208 19292
rect 29963 19261 29975 19264
rect 29917 19255 29975 19261
rect 31202 19252 31208 19264
rect 31260 19252 31266 19304
rect 36078 19292 36084 19304
rect 35991 19264 36084 19292
rect 36078 19252 36084 19264
rect 36136 19292 36142 19304
rect 36265 19295 36323 19301
rect 36265 19292 36277 19295
rect 36136 19264 36277 19292
rect 36136 19252 36142 19264
rect 36265 19261 36277 19264
rect 36311 19261 36323 19295
rect 36265 19255 36323 19261
rect 35529 19227 35587 19233
rect 35529 19193 35541 19227
rect 35575 19224 35587 19227
rect 36538 19224 36544 19236
rect 35575 19196 36544 19224
rect 35575 19193 35587 19196
rect 35529 19187 35587 19193
rect 36538 19184 36544 19196
rect 36596 19184 36602 19236
rect 27154 19156 27160 19168
rect 25924 19128 26280 19156
rect 27115 19128 27160 19156
rect 25924 19116 25930 19128
rect 27154 19116 27160 19128
rect 27212 19116 27218 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 4706 18952 4712 18964
rect 2700 18924 4712 18952
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18717 2191 18751
rect 2133 18711 2191 18717
rect 2317 18751 2375 18757
rect 2317 18717 2329 18751
rect 2363 18748 2375 18751
rect 2700 18748 2728 18924
rect 4706 18912 4712 18924
rect 4764 18912 4770 18964
rect 6917 18955 6975 18961
rect 6917 18921 6929 18955
rect 6963 18952 6975 18955
rect 7006 18952 7012 18964
rect 6963 18924 7012 18952
rect 6963 18921 6975 18924
rect 6917 18915 6975 18921
rect 7006 18912 7012 18924
rect 7064 18912 7070 18964
rect 12986 18912 12992 18964
rect 13044 18952 13050 18964
rect 13265 18955 13323 18961
rect 13265 18952 13277 18955
rect 13044 18924 13277 18952
rect 13044 18912 13050 18924
rect 13265 18921 13277 18924
rect 13311 18921 13323 18955
rect 13446 18952 13452 18964
rect 13407 18924 13452 18952
rect 13265 18915 13323 18921
rect 13446 18912 13452 18924
rect 13504 18912 13510 18964
rect 22189 18955 22247 18961
rect 22189 18921 22201 18955
rect 22235 18921 22247 18955
rect 23198 18952 23204 18964
rect 23159 18924 23204 18952
rect 22189 18915 22247 18921
rect 14734 18844 14740 18896
rect 14792 18884 14798 18896
rect 16761 18887 16819 18893
rect 16761 18884 16773 18887
rect 14792 18856 16773 18884
rect 14792 18844 14798 18856
rect 16761 18853 16773 18856
rect 16807 18853 16819 18887
rect 18506 18884 18512 18896
rect 16761 18847 16819 18853
rect 17144 18856 18512 18884
rect 4249 18819 4307 18825
rect 4249 18785 4261 18819
rect 4295 18816 4307 18819
rect 4614 18816 4620 18828
rect 4295 18788 4620 18816
rect 4295 18785 4307 18788
rect 4249 18779 4307 18785
rect 4614 18776 4620 18788
rect 4672 18776 4678 18828
rect 17144 18816 17172 18856
rect 18506 18844 18512 18856
rect 18564 18844 18570 18896
rect 22204 18884 22232 18915
rect 23198 18912 23204 18924
rect 23256 18912 23262 18964
rect 26234 18952 26240 18964
rect 25516 18924 26240 18952
rect 25516 18884 25544 18924
rect 26234 18912 26240 18924
rect 26292 18912 26298 18964
rect 26878 18952 26884 18964
rect 26839 18924 26884 18952
rect 26878 18912 26884 18924
rect 26936 18912 26942 18964
rect 28258 18912 28264 18964
rect 28316 18952 28322 18964
rect 28445 18955 28503 18961
rect 28445 18952 28457 18955
rect 28316 18924 28457 18952
rect 28316 18912 28322 18924
rect 28445 18921 28457 18924
rect 28491 18921 28503 18955
rect 28445 18915 28503 18921
rect 22204 18856 25544 18884
rect 27522 18844 27528 18896
rect 27580 18884 27586 18896
rect 36078 18884 36084 18896
rect 27580 18856 28948 18884
rect 36039 18856 36084 18884
rect 27580 18844 27586 18856
rect 18877 18819 18935 18825
rect 16776 18788 17172 18816
rect 17236 18788 18552 18816
rect 2363 18720 2728 18748
rect 2777 18751 2835 18757
rect 2363 18717 2375 18720
rect 2317 18711 2375 18717
rect 2777 18717 2789 18751
rect 2823 18748 2835 18751
rect 2866 18748 2872 18760
rect 2823 18720 2872 18748
rect 2823 18717 2835 18720
rect 2777 18711 2835 18717
rect 2148 18680 2176 18711
rect 2866 18708 2872 18720
rect 2924 18708 2930 18760
rect 2958 18708 2964 18760
rect 3016 18748 3022 18760
rect 3970 18748 3976 18760
rect 3016 18720 3061 18748
rect 3931 18720 3976 18748
rect 3016 18708 3022 18720
rect 3970 18708 3976 18720
rect 4028 18708 4034 18760
rect 7098 18708 7104 18760
rect 7156 18708 7162 18760
rect 10045 18751 10103 18757
rect 10045 18717 10057 18751
rect 10091 18748 10103 18751
rect 10594 18748 10600 18760
rect 10091 18720 10600 18748
rect 10091 18717 10103 18720
rect 10045 18711 10103 18717
rect 10594 18708 10600 18720
rect 10652 18708 10658 18760
rect 16776 18757 16804 18788
rect 16577 18751 16635 18757
rect 16577 18717 16589 18751
rect 16623 18717 16635 18751
rect 16577 18711 16635 18717
rect 16761 18751 16819 18757
rect 16761 18717 16773 18751
rect 16807 18717 16819 18751
rect 16761 18711 16819 18717
rect 2148 18652 2774 18680
rect 2130 18572 2136 18624
rect 2188 18612 2194 18624
rect 2225 18615 2283 18621
rect 2225 18612 2237 18615
rect 2188 18584 2237 18612
rect 2188 18572 2194 18584
rect 2225 18581 2237 18584
rect 2271 18581 2283 18615
rect 2746 18612 2774 18652
rect 4890 18640 4896 18692
rect 4948 18640 4954 18692
rect 6730 18680 6736 18692
rect 6691 18652 6736 18680
rect 6730 18640 6736 18652
rect 6788 18640 6794 18692
rect 6917 18683 6975 18689
rect 6917 18649 6929 18683
rect 6963 18680 6975 18683
rect 7116 18680 7144 18708
rect 6963 18652 7144 18680
rect 6963 18649 6975 18652
rect 6917 18643 6975 18649
rect 10686 18640 10692 18692
rect 10744 18680 10750 18692
rect 13081 18683 13139 18689
rect 13081 18680 13093 18683
rect 10744 18652 13093 18680
rect 10744 18640 10750 18652
rect 13081 18649 13093 18652
rect 13127 18649 13139 18683
rect 16592 18680 16620 18711
rect 17236 18692 17264 18788
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 17589 18751 17647 18757
rect 17589 18717 17601 18751
rect 17635 18748 17647 18751
rect 17862 18748 17868 18760
rect 17635 18720 17868 18748
rect 17635 18717 17647 18720
rect 17589 18711 17647 18717
rect 17218 18680 17224 18692
rect 16592 18652 17224 18680
rect 13081 18643 13139 18649
rect 17218 18640 17224 18652
rect 17276 18640 17282 18692
rect 17420 18680 17448 18711
rect 17862 18708 17868 18720
rect 17920 18708 17926 18760
rect 18524 18757 18552 18788
rect 18877 18785 18889 18819
rect 18923 18816 18935 18819
rect 20254 18816 20260 18828
rect 18923 18788 20260 18816
rect 18923 18785 18935 18788
rect 18877 18779 18935 18785
rect 20254 18776 20260 18788
rect 20312 18776 20318 18828
rect 28920 18825 28948 18856
rect 36078 18844 36084 18856
rect 36136 18844 36142 18896
rect 28621 18819 28679 18825
rect 28621 18816 28633 18819
rect 28368 18788 28633 18816
rect 18509 18751 18567 18757
rect 18509 18717 18521 18751
rect 18555 18717 18567 18751
rect 18509 18711 18567 18717
rect 22370 18708 22376 18760
rect 22428 18748 22434 18760
rect 23385 18751 23443 18757
rect 23385 18748 23397 18751
rect 22428 18720 23397 18748
rect 22428 18708 22434 18720
rect 23385 18717 23397 18720
rect 23431 18717 23443 18751
rect 23658 18748 23664 18760
rect 23619 18720 23664 18748
rect 23385 18711 23443 18717
rect 18325 18683 18383 18689
rect 17420 18652 17632 18680
rect 17604 18624 17632 18652
rect 18325 18649 18337 18683
rect 18371 18680 18383 18683
rect 18690 18680 18696 18692
rect 18371 18652 18696 18680
rect 18371 18649 18383 18652
rect 18325 18643 18383 18649
rect 18690 18640 18696 18652
rect 18748 18640 18754 18692
rect 21910 18640 21916 18692
rect 21968 18680 21974 18692
rect 22005 18683 22063 18689
rect 22005 18680 22017 18683
rect 21968 18652 22017 18680
rect 21968 18640 21974 18652
rect 22005 18649 22017 18652
rect 22051 18649 22063 18683
rect 22186 18680 22192 18692
rect 22147 18652 22192 18680
rect 22005 18643 22063 18649
rect 22186 18640 22192 18652
rect 22244 18640 22250 18692
rect 2961 18615 3019 18621
rect 2961 18612 2973 18615
rect 2746 18584 2973 18612
rect 2225 18575 2283 18581
rect 2961 18581 2973 18584
rect 3007 18612 3019 18615
rect 4430 18612 4436 18624
rect 3007 18584 4436 18612
rect 3007 18581 3019 18584
rect 2961 18575 3019 18581
rect 4430 18572 4436 18584
rect 4488 18572 4494 18624
rect 5718 18612 5724 18624
rect 5679 18584 5724 18612
rect 5718 18572 5724 18584
rect 5776 18572 5782 18624
rect 7101 18615 7159 18621
rect 7101 18581 7113 18615
rect 7147 18612 7159 18615
rect 9122 18612 9128 18624
rect 7147 18584 9128 18612
rect 7147 18581 7159 18584
rect 7101 18575 7159 18581
rect 9122 18572 9128 18584
rect 9180 18572 9186 18624
rect 10134 18612 10140 18624
rect 10095 18584 10140 18612
rect 10134 18572 10140 18584
rect 10192 18572 10198 18624
rect 13265 18615 13323 18621
rect 13265 18581 13277 18615
rect 13311 18612 13323 18615
rect 14826 18612 14832 18624
rect 13311 18584 14832 18612
rect 13311 18581 13323 18584
rect 13265 18575 13323 18581
rect 14826 18572 14832 18584
rect 14884 18572 14890 18624
rect 16850 18572 16856 18624
rect 16908 18612 16914 18624
rect 17310 18612 17316 18624
rect 16908 18584 17316 18612
rect 16908 18572 16914 18584
rect 17310 18572 17316 18584
rect 17368 18612 17374 18624
rect 17405 18615 17463 18621
rect 17405 18612 17417 18615
rect 17368 18584 17417 18612
rect 17368 18572 17374 18584
rect 17405 18581 17417 18584
rect 17451 18581 17463 18615
rect 17405 18575 17463 18581
rect 17586 18572 17592 18624
rect 17644 18572 17650 18624
rect 22373 18615 22431 18621
rect 22373 18581 22385 18615
rect 22419 18612 22431 18615
rect 22554 18612 22560 18624
rect 22419 18584 22560 18612
rect 22419 18581 22431 18584
rect 22373 18575 22431 18581
rect 22554 18572 22560 18584
rect 22612 18572 22618 18624
rect 23400 18612 23428 18711
rect 23658 18708 23664 18720
rect 23716 18708 23722 18760
rect 25222 18708 25228 18760
rect 25280 18748 25286 18760
rect 25501 18751 25559 18757
rect 25501 18748 25513 18751
rect 25280 18720 25513 18748
rect 25280 18708 25286 18720
rect 25501 18717 25513 18720
rect 25547 18748 25559 18751
rect 26050 18748 26056 18760
rect 25547 18720 26056 18748
rect 25547 18717 25559 18720
rect 25501 18711 25559 18717
rect 26050 18708 26056 18720
rect 26108 18708 26114 18760
rect 23569 18683 23627 18689
rect 23569 18649 23581 18683
rect 23615 18680 23627 18683
rect 23842 18680 23848 18692
rect 23615 18652 23848 18680
rect 23615 18649 23627 18652
rect 23569 18643 23627 18649
rect 23842 18640 23848 18652
rect 23900 18640 23906 18692
rect 25768 18683 25826 18689
rect 25768 18649 25780 18683
rect 25814 18680 25826 18683
rect 27154 18680 27160 18692
rect 25814 18652 27160 18680
rect 25814 18649 25826 18652
rect 25768 18643 25826 18649
rect 27154 18640 27160 18652
rect 27212 18640 27218 18692
rect 25866 18612 25872 18624
rect 23400 18584 25872 18612
rect 25866 18572 25872 18584
rect 25924 18572 25930 18624
rect 28368 18612 28396 18788
rect 28621 18785 28633 18788
rect 28667 18785 28679 18819
rect 28621 18779 28679 18785
rect 28905 18819 28963 18825
rect 28905 18785 28917 18819
rect 28951 18785 28963 18819
rect 30374 18816 30380 18828
rect 30335 18788 30380 18816
rect 28905 18779 28963 18785
rect 30374 18776 30380 18788
rect 30432 18816 30438 18828
rect 30926 18816 30932 18828
rect 30432 18788 30932 18816
rect 30432 18776 30438 18788
rect 30926 18776 30932 18788
rect 30984 18776 30990 18828
rect 32953 18819 33011 18825
rect 32953 18785 32965 18819
rect 32999 18816 33011 18819
rect 33134 18816 33140 18828
rect 32999 18788 33140 18816
rect 32999 18785 33011 18788
rect 32953 18779 33011 18785
rect 33134 18776 33140 18788
rect 33192 18776 33198 18828
rect 28442 18708 28448 18760
rect 28500 18748 28506 18760
rect 28699 18751 28757 18757
rect 28699 18748 28711 18751
rect 28500 18720 28711 18748
rect 28500 18708 28506 18720
rect 28699 18717 28711 18720
rect 28745 18717 28757 18751
rect 28699 18711 28757 18717
rect 28814 18751 28872 18757
rect 28814 18717 28826 18751
rect 28860 18748 28872 18751
rect 30101 18751 30159 18757
rect 28860 18720 29960 18748
rect 28860 18717 28872 18720
rect 28814 18711 28872 18717
rect 29932 18689 29960 18720
rect 30101 18717 30113 18751
rect 30147 18748 30159 18751
rect 31018 18748 31024 18760
rect 30147 18720 31024 18748
rect 30147 18717 30159 18720
rect 30101 18711 30159 18717
rect 31018 18708 31024 18720
rect 31076 18708 31082 18760
rect 33778 18748 33784 18760
rect 33442 18720 33784 18748
rect 33778 18708 33784 18720
rect 33836 18708 33842 18760
rect 35710 18748 35716 18760
rect 35671 18720 35716 18748
rect 35710 18708 35716 18720
rect 35768 18708 35774 18760
rect 35897 18751 35955 18757
rect 35897 18717 35909 18751
rect 35943 18717 35955 18751
rect 35897 18711 35955 18717
rect 29917 18683 29975 18689
rect 29917 18649 29929 18683
rect 29963 18680 29975 18683
rect 30834 18680 30840 18692
rect 29963 18652 30840 18680
rect 29963 18649 29975 18652
rect 29917 18643 29975 18649
rect 30834 18640 30840 18652
rect 30892 18640 30898 18692
rect 33505 18683 33563 18689
rect 33505 18649 33517 18683
rect 33551 18649 33563 18683
rect 33505 18643 33563 18649
rect 30190 18612 30196 18624
rect 28368 18584 30196 18612
rect 30190 18572 30196 18584
rect 30248 18572 30254 18624
rect 31018 18572 31024 18624
rect 31076 18612 31082 18624
rect 33520 18612 33548 18643
rect 35342 18640 35348 18692
rect 35400 18680 35406 18692
rect 35912 18680 35940 18711
rect 35986 18708 35992 18760
rect 36044 18748 36050 18760
rect 36173 18751 36231 18757
rect 36173 18748 36185 18751
rect 36044 18720 36185 18748
rect 36044 18708 36050 18720
rect 36173 18717 36185 18720
rect 36219 18717 36231 18751
rect 36446 18748 36452 18760
rect 36407 18720 36452 18748
rect 36173 18711 36231 18717
rect 36446 18708 36452 18720
rect 36504 18708 36510 18760
rect 35400 18652 35940 18680
rect 35400 18640 35406 18652
rect 31076 18584 33548 18612
rect 31076 18572 31082 18584
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 3605 18411 3663 18417
rect 3605 18377 3617 18411
rect 3651 18377 3663 18411
rect 3605 18371 3663 18377
rect 2130 18340 2136 18352
rect 2091 18312 2136 18340
rect 2130 18300 2136 18312
rect 2188 18300 2194 18352
rect 2774 18300 2780 18352
rect 2832 18300 2838 18352
rect 3620 18272 3648 18371
rect 3970 18368 3976 18420
rect 4028 18408 4034 18420
rect 4065 18411 4123 18417
rect 4065 18408 4077 18411
rect 4028 18380 4077 18408
rect 4028 18368 4034 18380
rect 4065 18377 4077 18380
rect 4111 18377 4123 18411
rect 13354 18408 13360 18420
rect 4065 18371 4123 18377
rect 12406 18380 13360 18408
rect 12406 18340 12434 18380
rect 13354 18368 13360 18380
rect 13412 18368 13418 18420
rect 14277 18411 14335 18417
rect 14277 18377 14289 18411
rect 14323 18408 14335 18411
rect 15562 18408 15568 18420
rect 14323 18380 15568 18408
rect 14323 18377 14335 18380
rect 14277 18371 14335 18377
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 15930 18368 15936 18420
rect 15988 18408 15994 18420
rect 17221 18411 17279 18417
rect 17221 18408 17233 18411
rect 15988 18380 17233 18408
rect 15988 18368 15994 18380
rect 17221 18377 17233 18380
rect 17267 18377 17279 18411
rect 26050 18408 26056 18420
rect 26011 18380 26056 18408
rect 17221 18371 17279 18377
rect 26050 18368 26056 18380
rect 26108 18368 26114 18420
rect 29638 18368 29644 18420
rect 29696 18408 29702 18420
rect 29917 18411 29975 18417
rect 29917 18408 29929 18411
rect 29696 18380 29929 18408
rect 29696 18368 29702 18380
rect 29917 18377 29929 18380
rect 29963 18377 29975 18411
rect 29917 18371 29975 18377
rect 32214 18368 32220 18420
rect 32272 18408 32278 18420
rect 35805 18411 35863 18417
rect 35805 18408 35817 18411
rect 32272 18380 35817 18408
rect 32272 18368 32278 18380
rect 10428 18312 12434 18340
rect 13164 18343 13222 18349
rect 4249 18275 4307 18281
rect 4249 18272 4261 18275
rect 3620 18244 4261 18272
rect 4249 18241 4261 18244
rect 4295 18241 4307 18275
rect 4798 18272 4804 18284
rect 4249 18235 4307 18241
rect 4448 18244 4804 18272
rect 1857 18207 1915 18213
rect 1857 18173 1869 18207
rect 1903 18204 1915 18207
rect 2682 18204 2688 18216
rect 1903 18176 2688 18204
rect 1903 18173 1915 18176
rect 1857 18167 1915 18173
rect 2682 18164 2688 18176
rect 2740 18204 2746 18216
rect 4448 18204 4476 18244
rect 4798 18232 4804 18244
rect 4856 18272 4862 18284
rect 5442 18272 5448 18284
rect 4856 18244 5448 18272
rect 4856 18232 4862 18244
rect 5442 18232 5448 18244
rect 5500 18232 5506 18284
rect 7837 18275 7895 18281
rect 7837 18241 7849 18275
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 2740 18176 4476 18204
rect 4525 18207 4583 18213
rect 2740 18164 2746 18176
rect 4525 18173 4537 18207
rect 4571 18204 4583 18207
rect 4706 18204 4712 18216
rect 4571 18176 4712 18204
rect 4571 18173 4583 18176
rect 4525 18167 4583 18173
rect 4706 18164 4712 18176
rect 4764 18164 4770 18216
rect 4430 18136 4436 18148
rect 4391 18108 4436 18136
rect 4430 18096 4436 18108
rect 4488 18096 4494 18148
rect 7852 18136 7880 18235
rect 9214 18232 9220 18284
rect 9272 18272 9278 18284
rect 10428 18281 10456 18312
rect 13164 18309 13176 18343
rect 13210 18340 13222 18343
rect 13814 18340 13820 18352
rect 13210 18312 13820 18340
rect 13210 18309 13222 18312
rect 13164 18303 13222 18309
rect 13814 18300 13820 18312
rect 13872 18300 13878 18352
rect 17862 18300 17868 18352
rect 17920 18340 17926 18352
rect 18325 18343 18383 18349
rect 18325 18340 18337 18343
rect 17920 18312 18337 18340
rect 17920 18300 17926 18312
rect 18325 18309 18337 18312
rect 18371 18309 18383 18343
rect 18874 18340 18880 18352
rect 18835 18312 18880 18340
rect 18325 18303 18383 18309
rect 18874 18300 18880 18312
rect 18932 18300 18938 18352
rect 22554 18340 22560 18352
rect 22515 18312 22560 18340
rect 22554 18300 22560 18312
rect 22612 18300 22618 18352
rect 10312 18275 10370 18281
rect 10312 18272 10324 18275
rect 9272 18244 10324 18272
rect 9272 18232 9278 18244
rect 10312 18241 10324 18244
rect 10358 18241 10370 18275
rect 10312 18235 10370 18241
rect 10413 18275 10471 18281
rect 10413 18241 10425 18275
rect 10459 18241 10471 18275
rect 10594 18272 10600 18284
rect 10555 18244 10600 18272
rect 10413 18235 10471 18241
rect 10594 18232 10600 18244
rect 10652 18232 10658 18284
rect 12894 18272 12900 18284
rect 12855 18244 12900 18272
rect 12894 18232 12900 18244
rect 12952 18232 12958 18284
rect 17218 18272 17224 18284
rect 17179 18244 17224 18272
rect 17218 18232 17224 18244
rect 17276 18232 17282 18284
rect 17586 18272 17592 18284
rect 17547 18244 17592 18272
rect 17586 18232 17592 18244
rect 17644 18232 17650 18284
rect 18506 18272 18512 18284
rect 18467 18244 18512 18272
rect 18506 18232 18512 18244
rect 18564 18232 18570 18284
rect 18598 18232 18604 18284
rect 18656 18272 18662 18284
rect 19337 18275 19395 18281
rect 19337 18272 19349 18275
rect 18656 18244 19349 18272
rect 18656 18232 18662 18244
rect 19337 18241 19349 18244
rect 19383 18241 19395 18275
rect 19337 18235 19395 18241
rect 19521 18275 19579 18281
rect 19521 18241 19533 18275
rect 19567 18241 19579 18275
rect 19521 18235 19579 18241
rect 24765 18275 24823 18281
rect 24765 18241 24777 18275
rect 24811 18272 24823 18275
rect 26234 18272 26240 18284
rect 24811 18244 26240 18272
rect 24811 18241 24823 18244
rect 24765 18235 24823 18241
rect 9398 18164 9404 18216
rect 9456 18204 9462 18216
rect 11057 18207 11115 18213
rect 11057 18204 11069 18207
rect 9456 18176 11069 18204
rect 9456 18164 9462 18176
rect 11057 18173 11069 18176
rect 11103 18173 11115 18207
rect 17236 18204 17264 18232
rect 19536 18204 19564 18235
rect 26234 18232 26240 18244
rect 26292 18232 26298 18284
rect 28626 18272 28632 18284
rect 28587 18244 28632 18272
rect 28626 18232 28632 18244
rect 28684 18232 28690 18284
rect 30834 18272 30840 18284
rect 30795 18244 30840 18272
rect 30834 18232 30840 18244
rect 30892 18232 30898 18284
rect 31018 18272 31024 18284
rect 30979 18244 31024 18272
rect 31018 18232 31024 18244
rect 31076 18232 31082 18284
rect 32766 18272 32772 18284
rect 32727 18244 32772 18272
rect 32766 18232 32772 18244
rect 32824 18232 32830 18284
rect 33152 18281 33180 18380
rect 35805 18377 35817 18380
rect 35851 18408 35863 18411
rect 35986 18408 35992 18420
rect 35851 18380 35992 18408
rect 35851 18377 35863 18380
rect 35805 18371 35863 18377
rect 35986 18368 35992 18380
rect 36044 18368 36050 18420
rect 36170 18408 36176 18420
rect 36131 18380 36176 18408
rect 36170 18368 36176 18380
rect 36228 18368 36234 18420
rect 35621 18343 35679 18349
rect 35621 18340 35633 18343
rect 33336 18312 35633 18340
rect 33336 18284 33364 18312
rect 33137 18275 33195 18281
rect 33137 18241 33149 18275
rect 33183 18241 33195 18275
rect 33318 18272 33324 18284
rect 33279 18244 33324 18272
rect 33137 18235 33195 18241
rect 33318 18232 33324 18244
rect 33376 18232 33382 18284
rect 34992 18281 35020 18312
rect 35621 18309 35633 18312
rect 35667 18340 35679 18343
rect 35710 18340 35716 18352
rect 35667 18312 35716 18340
rect 35667 18309 35679 18312
rect 35621 18303 35679 18309
rect 35710 18300 35716 18312
rect 35768 18300 35774 18352
rect 35897 18343 35955 18349
rect 35897 18309 35909 18343
rect 35943 18340 35955 18343
rect 36446 18340 36452 18352
rect 35943 18312 36452 18340
rect 35943 18309 35955 18312
rect 35897 18303 35955 18309
rect 36446 18300 36452 18312
rect 36504 18300 36510 18352
rect 33689 18275 33747 18281
rect 33689 18241 33701 18275
rect 33735 18241 33747 18275
rect 34517 18275 34575 18281
rect 34517 18272 34529 18275
rect 33689 18235 33747 18241
rect 33796 18244 34529 18272
rect 17236 18176 19564 18204
rect 19889 18207 19947 18213
rect 11057 18167 11115 18173
rect 19889 18173 19901 18207
rect 19935 18204 19947 18207
rect 27430 18204 27436 18216
rect 19935 18176 27436 18204
rect 19935 18173 19947 18176
rect 19889 18167 19947 18173
rect 27430 18164 27436 18176
rect 27488 18164 27494 18216
rect 30852 18204 30880 18232
rect 32858 18204 32864 18216
rect 30852 18176 32864 18204
rect 32858 18164 32864 18176
rect 32916 18164 32922 18216
rect 32953 18207 33011 18213
rect 32953 18173 32965 18207
rect 32999 18204 33011 18207
rect 33594 18204 33600 18216
rect 32999 18176 33600 18204
rect 32999 18173 33011 18176
rect 32953 18167 33011 18173
rect 33594 18164 33600 18176
rect 33652 18164 33658 18216
rect 16482 18136 16488 18148
rect 7852 18108 12434 18136
rect 5442 18028 5448 18080
rect 5500 18068 5506 18080
rect 9125 18071 9183 18077
rect 9125 18068 9137 18071
rect 5500 18040 9137 18068
rect 5500 18028 5506 18040
rect 9125 18037 9137 18040
rect 9171 18068 9183 18071
rect 10686 18068 10692 18080
rect 9171 18040 10692 18068
rect 9171 18037 9183 18040
rect 9125 18031 9183 18037
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 12406 18068 12434 18108
rect 14200 18108 16488 18136
rect 14200 18068 14228 18108
rect 16482 18096 16488 18108
rect 16540 18096 16546 18148
rect 32582 18096 32588 18148
rect 32640 18136 32646 18148
rect 33704 18136 33732 18235
rect 32640 18108 33732 18136
rect 32640 18096 32646 18108
rect 12406 18040 14228 18068
rect 20806 18028 20812 18080
rect 20864 18068 20870 18080
rect 23845 18071 23903 18077
rect 23845 18068 23857 18071
rect 20864 18040 23857 18068
rect 20864 18028 20870 18040
rect 23845 18037 23857 18040
rect 23891 18037 23903 18071
rect 23845 18031 23903 18037
rect 28994 18028 29000 18080
rect 29052 18068 29058 18080
rect 30929 18071 30987 18077
rect 30929 18068 30941 18071
rect 29052 18040 30941 18068
rect 29052 18028 29058 18040
rect 30929 18037 30941 18040
rect 30975 18037 30987 18071
rect 30929 18031 30987 18037
rect 32766 18028 32772 18080
rect 32824 18068 32830 18080
rect 33796 18068 33824 18244
rect 34517 18241 34529 18244
rect 34563 18241 34575 18275
rect 34517 18235 34575 18241
rect 34977 18275 35035 18281
rect 34977 18241 34989 18275
rect 35023 18241 35035 18275
rect 34977 18235 35035 18241
rect 35989 18275 36047 18281
rect 35989 18241 36001 18275
rect 36035 18241 36047 18275
rect 35989 18235 36047 18241
rect 34790 18204 34796 18216
rect 34703 18176 34796 18204
rect 34790 18164 34796 18176
rect 34848 18204 34854 18216
rect 35710 18204 35716 18216
rect 34848 18176 35716 18204
rect 34848 18164 34854 18176
rect 35710 18164 35716 18176
rect 35768 18164 35774 18216
rect 36004 18204 36032 18235
rect 35912 18176 36032 18204
rect 35342 18096 35348 18148
rect 35400 18136 35406 18148
rect 35912 18136 35940 18176
rect 35400 18108 35940 18136
rect 35400 18096 35406 18108
rect 32824 18040 33824 18068
rect 32824 18028 32830 18040
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 10594 17864 10600 17876
rect 2832 17836 2877 17864
rect 8588 17836 10600 17864
rect 2832 17824 2838 17836
rect 1394 17688 1400 17740
rect 1452 17728 1458 17740
rect 1452 17700 8432 17728
rect 1452 17688 1458 17700
rect 2774 17620 2780 17672
rect 2832 17660 2838 17672
rect 2961 17663 3019 17669
rect 2832 17632 2877 17660
rect 2832 17620 2838 17632
rect 2961 17629 2973 17663
rect 3007 17660 3019 17663
rect 5074 17660 5080 17672
rect 3007 17632 5080 17660
rect 3007 17629 3019 17632
rect 2961 17623 3019 17629
rect 5074 17620 5080 17632
rect 5132 17620 5138 17672
rect 8205 17595 8263 17601
rect 8205 17561 8217 17595
rect 8251 17592 8263 17595
rect 8294 17592 8300 17604
rect 8251 17564 8300 17592
rect 8251 17561 8263 17564
rect 8205 17555 8263 17561
rect 8294 17552 8300 17564
rect 8352 17552 8358 17604
rect 8404 17592 8432 17700
rect 8478 17620 8484 17672
rect 8536 17660 8542 17672
rect 8588 17660 8616 17836
rect 10594 17824 10600 17836
rect 10652 17824 10658 17876
rect 22002 17824 22008 17876
rect 22060 17864 22066 17876
rect 22097 17867 22155 17873
rect 22097 17864 22109 17867
rect 22060 17836 22109 17864
rect 22060 17824 22066 17836
rect 22097 17833 22109 17836
rect 22143 17833 22155 17867
rect 22097 17827 22155 17833
rect 24857 17867 24915 17873
rect 24857 17833 24869 17867
rect 24903 17864 24915 17867
rect 25038 17864 25044 17876
rect 24903 17836 25044 17864
rect 24903 17833 24915 17836
rect 24857 17827 24915 17833
rect 25038 17824 25044 17836
rect 25096 17864 25102 17876
rect 25406 17864 25412 17876
rect 25096 17836 25412 17864
rect 25096 17824 25102 17836
rect 25406 17824 25412 17836
rect 25464 17824 25470 17876
rect 27798 17824 27804 17876
rect 27856 17864 27862 17876
rect 28261 17867 28319 17873
rect 28261 17864 28273 17867
rect 27856 17836 28273 17864
rect 27856 17824 27862 17836
rect 28261 17833 28273 17836
rect 28307 17833 28319 17867
rect 33410 17864 33416 17876
rect 33371 17836 33416 17864
rect 28261 17827 28319 17833
rect 33410 17824 33416 17836
rect 33468 17824 33474 17876
rect 21542 17756 21548 17808
rect 21600 17796 21606 17808
rect 23474 17796 23480 17808
rect 21600 17768 23480 17796
rect 21600 17756 21606 17768
rect 23474 17756 23480 17768
rect 23532 17756 23538 17808
rect 28994 17796 29000 17808
rect 28552 17768 29000 17796
rect 28442 17728 28448 17740
rect 8680 17700 12480 17728
rect 8536 17632 8629 17660
rect 8536 17620 8542 17632
rect 8680 17592 8708 17700
rect 9122 17660 9128 17672
rect 9083 17632 9128 17660
rect 9122 17620 9128 17632
rect 9180 17620 9186 17672
rect 12158 17620 12164 17672
rect 12216 17660 12222 17672
rect 12345 17663 12403 17669
rect 12345 17660 12357 17663
rect 12216 17632 12357 17660
rect 12216 17620 12222 17632
rect 12345 17629 12357 17632
rect 12391 17629 12403 17663
rect 12452 17660 12480 17700
rect 20548 17700 28448 17728
rect 15381 17663 15439 17669
rect 15381 17660 15393 17663
rect 12452 17632 15393 17660
rect 12345 17623 12403 17629
rect 15381 17629 15393 17632
rect 15427 17629 15439 17663
rect 15381 17623 15439 17629
rect 17402 17620 17408 17672
rect 17460 17660 17466 17672
rect 17862 17660 17868 17672
rect 17460 17632 17868 17660
rect 17460 17620 17466 17632
rect 17862 17620 17868 17632
rect 17920 17660 17926 17672
rect 18141 17663 18199 17669
rect 18141 17660 18153 17663
rect 17920 17632 18153 17660
rect 17920 17620 17926 17632
rect 18141 17629 18153 17632
rect 18187 17629 18199 17663
rect 18690 17660 18696 17672
rect 18603 17632 18696 17660
rect 18141 17623 18199 17629
rect 18690 17620 18696 17632
rect 18748 17660 18754 17672
rect 19242 17660 19248 17672
rect 18748 17632 19248 17660
rect 18748 17620 18754 17632
rect 19242 17620 19248 17632
rect 19300 17620 19306 17672
rect 9398 17592 9404 17604
rect 8404 17564 8708 17592
rect 9359 17564 9404 17592
rect 9398 17552 9404 17564
rect 9456 17552 9462 17604
rect 10778 17592 10784 17604
rect 10626 17564 10784 17592
rect 10778 17552 10784 17564
rect 10836 17552 10842 17604
rect 12612 17595 12670 17601
rect 12612 17561 12624 17595
rect 12658 17592 12670 17595
rect 13354 17592 13360 17604
rect 12658 17564 13360 17592
rect 12658 17561 12670 17564
rect 12612 17555 12670 17561
rect 13354 17552 13360 17564
rect 13412 17552 13418 17604
rect 18877 17595 18935 17601
rect 18877 17561 18889 17595
rect 18923 17561 18935 17595
rect 20548 17592 20576 17700
rect 28442 17688 28448 17700
rect 28500 17688 28506 17740
rect 28552 17737 28580 17768
rect 28994 17756 29000 17768
rect 29052 17756 29058 17808
rect 28537 17731 28595 17737
rect 28537 17697 28549 17731
rect 28583 17697 28595 17731
rect 30374 17728 30380 17740
rect 28537 17691 28595 17697
rect 28644 17700 30380 17728
rect 20622 17620 20628 17672
rect 20680 17660 20686 17672
rect 23201 17663 23259 17669
rect 23201 17660 23213 17663
rect 20680 17632 23213 17660
rect 20680 17620 20686 17632
rect 23201 17629 23213 17632
rect 23247 17629 23259 17663
rect 23474 17660 23480 17672
rect 23435 17632 23480 17660
rect 23201 17623 23259 17629
rect 23474 17620 23480 17632
rect 23532 17620 23538 17672
rect 28644 17669 28672 17700
rect 30374 17688 30380 17700
rect 30432 17688 30438 17740
rect 33594 17728 33600 17740
rect 33555 17700 33600 17728
rect 33594 17688 33600 17700
rect 33652 17688 33658 17740
rect 25133 17663 25191 17669
rect 25133 17629 25145 17663
rect 25179 17660 25191 17663
rect 25593 17663 25651 17669
rect 25593 17660 25605 17663
rect 25179 17632 25605 17660
rect 25179 17629 25191 17632
rect 25133 17623 25191 17629
rect 25593 17629 25605 17632
rect 25639 17629 25651 17663
rect 25593 17623 25651 17629
rect 28629 17663 28687 17669
rect 28629 17629 28641 17663
rect 28675 17629 28687 17663
rect 28629 17623 28687 17629
rect 28721 17663 28779 17669
rect 28721 17629 28733 17663
rect 28767 17629 28779 17663
rect 29730 17660 29736 17672
rect 29691 17632 29736 17660
rect 28721 17623 28779 17629
rect 20806 17592 20812 17604
rect 18877 17555 18935 17561
rect 19306 17564 20576 17592
rect 20767 17564 20812 17592
rect 6822 17484 6828 17536
rect 6880 17524 6886 17536
rect 7911 17527 7969 17533
rect 7911 17524 7923 17527
rect 6880 17496 7923 17524
rect 6880 17484 6886 17496
rect 7911 17493 7923 17496
rect 7957 17493 7969 17527
rect 7911 17487 7969 17493
rect 8389 17527 8447 17533
rect 8389 17493 8401 17527
rect 8435 17524 8447 17527
rect 10134 17524 10140 17536
rect 8435 17496 10140 17524
rect 8435 17493 8447 17496
rect 8389 17487 8447 17493
rect 10134 17484 10140 17496
rect 10192 17484 10198 17536
rect 10873 17527 10931 17533
rect 10873 17493 10885 17527
rect 10919 17524 10931 17527
rect 10962 17524 10968 17536
rect 10919 17496 10968 17524
rect 10919 17493 10931 17496
rect 10873 17487 10931 17493
rect 10962 17484 10968 17496
rect 11020 17484 11026 17536
rect 13722 17524 13728 17536
rect 13683 17496 13728 17524
rect 13722 17484 13728 17496
rect 13780 17484 13786 17536
rect 16482 17484 16488 17536
rect 16540 17524 16546 17536
rect 16669 17527 16727 17533
rect 16669 17524 16681 17527
rect 16540 17496 16681 17524
rect 16540 17484 16546 17496
rect 16669 17493 16681 17496
rect 16715 17493 16727 17527
rect 16669 17487 16727 17493
rect 17310 17484 17316 17536
rect 17368 17524 17374 17536
rect 18414 17524 18420 17536
rect 17368 17496 18420 17524
rect 17368 17484 17374 17496
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 18892 17524 18920 17555
rect 19306 17524 19334 17564
rect 20806 17552 20812 17564
rect 20864 17552 20870 17604
rect 21910 17552 21916 17604
rect 21968 17592 21974 17604
rect 24673 17595 24731 17601
rect 24673 17592 24685 17595
rect 21968 17564 24685 17592
rect 21968 17552 21974 17564
rect 24673 17561 24685 17564
rect 24719 17561 24731 17595
rect 24854 17592 24860 17604
rect 24815 17564 24860 17592
rect 24673 17555 24731 17561
rect 24854 17552 24860 17564
rect 24912 17552 24918 17604
rect 27246 17552 27252 17604
rect 27304 17592 27310 17604
rect 28736 17592 28764 17623
rect 29730 17620 29736 17632
rect 29788 17620 29794 17672
rect 32214 17620 32220 17672
rect 32272 17660 32278 17672
rect 32309 17663 32367 17669
rect 32309 17660 32321 17663
rect 32272 17632 32321 17660
rect 32272 17620 32278 17632
rect 32309 17629 32321 17632
rect 32355 17629 32367 17663
rect 32582 17660 32588 17672
rect 32543 17632 32588 17660
rect 32309 17623 32367 17629
rect 32582 17620 32588 17632
rect 32640 17660 32646 17672
rect 33042 17660 33048 17672
rect 32640 17632 33048 17660
rect 32640 17620 32646 17632
rect 33042 17620 33048 17632
rect 33100 17620 33106 17672
rect 33778 17660 33784 17672
rect 33739 17632 33784 17660
rect 33778 17620 33784 17632
rect 33836 17620 33842 17672
rect 34149 17663 34207 17669
rect 34149 17629 34161 17663
rect 34195 17629 34207 17663
rect 34149 17623 34207 17629
rect 34333 17663 34391 17669
rect 34333 17629 34345 17663
rect 34379 17660 34391 17663
rect 34790 17660 34796 17672
rect 34379 17632 34796 17660
rect 34379 17629 34391 17632
rect 34333 17623 34391 17629
rect 32674 17592 32680 17604
rect 27304 17564 28764 17592
rect 32635 17564 32680 17592
rect 27304 17552 27310 17564
rect 32674 17552 32680 17564
rect 32732 17592 32738 17604
rect 34164 17592 34192 17623
rect 34790 17620 34796 17632
rect 34848 17620 34854 17672
rect 32732 17564 34192 17592
rect 32732 17552 32738 17564
rect 23014 17524 23020 17536
rect 18892 17496 19334 17524
rect 22975 17496 23020 17524
rect 23014 17484 23020 17496
rect 23072 17484 23078 17536
rect 23382 17524 23388 17536
rect 23343 17496 23388 17524
rect 23382 17484 23388 17496
rect 23440 17484 23446 17536
rect 24872 17524 24900 17552
rect 25130 17524 25136 17536
rect 24872 17496 25136 17524
rect 25130 17484 25136 17496
rect 25188 17484 25194 17536
rect 26234 17484 26240 17536
rect 26292 17524 26298 17536
rect 26881 17527 26939 17533
rect 26881 17524 26893 17527
rect 26292 17496 26893 17524
rect 26292 17484 26298 17496
rect 26881 17493 26893 17496
rect 26927 17493 26939 17527
rect 26881 17487 26939 17493
rect 28626 17484 28632 17536
rect 28684 17524 28690 17536
rect 31021 17527 31079 17533
rect 31021 17524 31033 17527
rect 28684 17496 31033 17524
rect 28684 17484 28690 17496
rect 31021 17493 31033 17496
rect 31067 17493 31079 17527
rect 31021 17487 31079 17493
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 5718 17320 5724 17332
rect 5552 17292 5724 17320
rect 5350 17184 5356 17196
rect 5311 17156 5356 17184
rect 5350 17144 5356 17156
rect 5408 17144 5414 17196
rect 5552 17193 5580 17292
rect 5718 17280 5724 17292
rect 5776 17320 5782 17332
rect 8478 17320 8484 17332
rect 5776 17292 8484 17320
rect 5776 17280 5782 17292
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 10045 17323 10103 17329
rect 10045 17289 10057 17323
rect 10091 17320 10103 17323
rect 10318 17320 10324 17332
rect 10091 17292 10324 17320
rect 10091 17289 10103 17292
rect 10045 17283 10103 17289
rect 10318 17280 10324 17292
rect 10376 17280 10382 17332
rect 18138 17280 18144 17332
rect 18196 17320 18202 17332
rect 18877 17323 18935 17329
rect 18877 17320 18889 17323
rect 18196 17292 18889 17320
rect 18196 17280 18202 17292
rect 18877 17289 18889 17292
rect 18923 17289 18935 17323
rect 18877 17283 18935 17289
rect 21361 17323 21419 17329
rect 21361 17289 21373 17323
rect 21407 17320 21419 17323
rect 22370 17320 22376 17332
rect 21407 17292 22376 17320
rect 21407 17289 21419 17292
rect 21361 17283 21419 17289
rect 22370 17280 22376 17292
rect 22428 17280 22434 17332
rect 30190 17280 30196 17332
rect 30248 17320 30254 17332
rect 32493 17323 32551 17329
rect 32493 17320 32505 17323
rect 30248 17292 32505 17320
rect 30248 17280 30254 17292
rect 32493 17289 32505 17292
rect 32539 17289 32551 17323
rect 33134 17320 33140 17332
rect 33095 17292 33140 17320
rect 32493 17283 32551 17289
rect 33134 17280 33140 17292
rect 33192 17280 33198 17332
rect 5902 17212 5908 17264
rect 5960 17252 5966 17264
rect 7377 17255 7435 17261
rect 7377 17252 7389 17255
rect 5960 17224 7389 17252
rect 5960 17212 5966 17224
rect 7377 17221 7389 17224
rect 7423 17252 7435 17255
rect 7423 17224 10916 17252
rect 7423 17221 7435 17224
rect 7377 17215 7435 17221
rect 5537 17187 5595 17193
rect 5537 17153 5549 17187
rect 5583 17153 5595 17187
rect 5537 17147 5595 17153
rect 6733 17187 6791 17193
rect 6733 17153 6745 17187
rect 6779 17184 6791 17187
rect 7650 17184 7656 17196
rect 6779 17156 7656 17184
rect 6779 17153 6791 17156
rect 6733 17147 6791 17153
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 10686 17184 10692 17196
rect 10647 17156 10692 17184
rect 10686 17144 10692 17156
rect 10744 17144 10750 17196
rect 10888 17193 10916 17224
rect 10962 17212 10968 17264
rect 11020 17252 11026 17264
rect 11020 17224 16896 17252
rect 11020 17212 11026 17224
rect 10873 17187 10931 17193
rect 10873 17153 10885 17187
rect 10919 17153 10931 17187
rect 10873 17147 10931 17153
rect 12980 17187 13038 17193
rect 12980 17153 12992 17187
rect 13026 17184 13038 17187
rect 13262 17184 13268 17196
rect 13026 17156 13268 17184
rect 13026 17153 13038 17156
rect 12980 17147 13038 17153
rect 13262 17144 13268 17156
rect 13320 17144 13326 17196
rect 14642 17184 14648 17196
rect 14603 17156 14648 17184
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 16868 17193 16896 17224
rect 18046 17212 18052 17264
rect 18104 17252 18110 17264
rect 18601 17255 18659 17261
rect 18601 17252 18613 17255
rect 18104 17224 18613 17252
rect 18104 17212 18110 17224
rect 18601 17221 18613 17224
rect 18647 17221 18659 17255
rect 18601 17215 18659 17221
rect 21910 17212 21916 17264
rect 21968 17252 21974 17264
rect 32585 17255 32643 17261
rect 21968 17224 23888 17252
rect 21968 17212 21974 17224
rect 16853 17187 16911 17193
rect 16853 17153 16865 17187
rect 16899 17184 16911 17187
rect 17310 17184 17316 17196
rect 16899 17156 17316 17184
rect 16899 17153 16911 17156
rect 16853 17147 16911 17153
rect 17310 17144 17316 17156
rect 17368 17144 17374 17196
rect 17497 17187 17555 17193
rect 17497 17153 17509 17187
rect 17543 17153 17555 17187
rect 18233 17187 18291 17193
rect 18233 17184 18245 17187
rect 17497 17147 17555 17153
rect 18156 17156 18245 17184
rect 5258 17116 5264 17128
rect 5171 17088 5264 17116
rect 5258 17076 5264 17088
rect 5316 17076 5322 17128
rect 5997 17119 6055 17125
rect 5997 17085 6009 17119
rect 6043 17085 6055 17119
rect 5997 17079 6055 17085
rect 10045 17119 10103 17125
rect 10045 17085 10057 17119
rect 10091 17085 10103 17119
rect 10045 17079 10103 17085
rect 10137 17119 10195 17125
rect 10137 17085 10149 17119
rect 10183 17116 10195 17119
rect 10594 17116 10600 17128
rect 10183 17088 10600 17116
rect 10183 17085 10195 17088
rect 10137 17079 10195 17085
rect 5276 16980 5304 17076
rect 5350 17008 5356 17060
rect 5408 17048 5414 17060
rect 6012 17048 6040 17079
rect 5408 17020 6040 17048
rect 10060 17048 10088 17079
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 12158 17076 12164 17128
rect 12216 17116 12222 17128
rect 12713 17119 12771 17125
rect 12713 17116 12725 17119
rect 12216 17088 12725 17116
rect 12216 17076 12222 17088
rect 12713 17085 12725 17088
rect 12759 17085 12771 17119
rect 15010 17116 15016 17128
rect 14971 17088 15016 17116
rect 12713 17079 12771 17085
rect 15010 17076 15016 17088
rect 15068 17076 15074 17128
rect 17512 17116 17540 17147
rect 16868 17088 17540 17116
rect 16868 17060 16896 17088
rect 10226 17048 10232 17060
rect 10060 17020 10232 17048
rect 5408 17008 5414 17020
rect 10226 17008 10232 17020
rect 10284 17008 10290 17060
rect 10778 17048 10784 17060
rect 10739 17020 10784 17048
rect 10778 17008 10784 17020
rect 10836 17008 10842 17060
rect 16850 17008 16856 17060
rect 16908 17008 16914 17060
rect 18156 17048 18184 17156
rect 18233 17153 18245 17156
rect 18279 17153 18291 17187
rect 18233 17147 18291 17153
rect 18322 17144 18328 17196
rect 18380 17184 18386 17196
rect 18509 17187 18567 17193
rect 18380 17156 18425 17184
rect 18380 17144 18386 17156
rect 18509 17153 18521 17187
rect 18555 17153 18567 17187
rect 18690 17184 18696 17196
rect 18748 17193 18754 17196
rect 18656 17156 18696 17184
rect 18509 17147 18567 17153
rect 18414 17076 18420 17128
rect 18472 17116 18478 17128
rect 18524 17116 18552 17147
rect 18690 17144 18696 17156
rect 18748 17147 18756 17193
rect 21174 17184 21180 17196
rect 21087 17156 21180 17184
rect 18748 17144 18754 17147
rect 21174 17144 21180 17156
rect 21232 17144 21238 17196
rect 21453 17187 21511 17193
rect 21453 17153 21465 17187
rect 21499 17184 21511 17187
rect 21542 17184 21548 17196
rect 21499 17156 21548 17184
rect 21499 17153 21511 17156
rect 21453 17147 21511 17153
rect 21542 17144 21548 17156
rect 21600 17144 21606 17196
rect 22002 17184 22008 17196
rect 21963 17156 22008 17184
rect 22002 17144 22008 17156
rect 22060 17144 22066 17196
rect 22272 17187 22330 17193
rect 22272 17153 22284 17187
rect 22318 17184 22330 17187
rect 23014 17184 23020 17196
rect 22318 17156 23020 17184
rect 22318 17153 22330 17156
rect 22272 17147 22330 17153
rect 23014 17144 23020 17156
rect 23072 17144 23078 17196
rect 23860 17193 23888 17224
rect 32585 17221 32597 17255
rect 32631 17252 32643 17255
rect 33410 17252 33416 17264
rect 32631 17224 33416 17252
rect 32631 17221 32643 17224
rect 32585 17215 32643 17221
rect 33410 17212 33416 17224
rect 33468 17212 33474 17264
rect 23845 17187 23903 17193
rect 23845 17153 23857 17187
rect 23891 17153 23903 17187
rect 23845 17147 23903 17153
rect 23934 17144 23940 17196
rect 23992 17184 23998 17196
rect 24101 17187 24159 17193
rect 24101 17184 24113 17187
rect 23992 17156 24113 17184
rect 23992 17144 23998 17156
rect 24101 17153 24113 17156
rect 24147 17153 24159 17187
rect 24101 17147 24159 17153
rect 32401 17187 32459 17193
rect 32401 17153 32413 17187
rect 32447 17153 32459 17187
rect 32401 17147 32459 17153
rect 18472 17088 18552 17116
rect 21192 17116 21220 17144
rect 21818 17116 21824 17128
rect 21192 17088 21824 17116
rect 18472 17076 18478 17088
rect 21818 17076 21824 17088
rect 21876 17076 21882 17128
rect 22002 17048 22008 17060
rect 18156 17020 22008 17048
rect 22002 17008 22008 17020
rect 22060 17008 22066 17060
rect 32416 17048 32444 17147
rect 32674 17144 32680 17196
rect 32732 17184 32738 17196
rect 33321 17187 33379 17193
rect 32732 17156 32777 17184
rect 32732 17144 32738 17156
rect 33321 17153 33333 17187
rect 33367 17184 33379 17187
rect 33502 17184 33508 17196
rect 33367 17156 33508 17184
rect 33367 17153 33379 17156
rect 33321 17147 33379 17153
rect 33502 17144 33508 17156
rect 33560 17144 33566 17196
rect 33597 17187 33655 17193
rect 33597 17153 33609 17187
rect 33643 17153 33655 17187
rect 33597 17147 33655 17153
rect 33781 17187 33839 17193
rect 33781 17153 33793 17187
rect 33827 17184 33839 17187
rect 34790 17184 34796 17196
rect 33827 17156 34796 17184
rect 33827 17153 33839 17156
rect 33781 17147 33839 17153
rect 32692 17116 32720 17144
rect 33226 17116 33232 17128
rect 32692 17088 33232 17116
rect 33226 17076 33232 17088
rect 33284 17116 33290 17128
rect 33612 17116 33640 17147
rect 34790 17144 34796 17156
rect 34848 17144 34854 17196
rect 33284 17088 33640 17116
rect 33284 17076 33290 17088
rect 33502 17048 33508 17060
rect 32416 17020 33508 17048
rect 33502 17008 33508 17020
rect 33560 17008 33566 17060
rect 6546 16980 6552 16992
rect 5276 16952 6552 16980
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 9490 16940 9496 16992
rect 9548 16980 9554 16992
rect 9585 16983 9643 16989
rect 9585 16980 9597 16983
rect 9548 16952 9597 16980
rect 9548 16940 9554 16952
rect 9585 16949 9597 16952
rect 9631 16949 9643 16983
rect 14090 16980 14096 16992
rect 14051 16952 14096 16980
rect 9585 16943 9643 16949
rect 14090 16940 14096 16952
rect 14148 16940 14154 16992
rect 17313 16983 17371 16989
rect 17313 16949 17325 16983
rect 17359 16980 17371 16983
rect 17402 16980 17408 16992
rect 17359 16952 17408 16980
rect 17359 16949 17371 16952
rect 17313 16943 17371 16949
rect 17402 16940 17408 16952
rect 17460 16940 17466 16992
rect 20993 16983 21051 16989
rect 20993 16949 21005 16983
rect 21039 16980 21051 16983
rect 21082 16980 21088 16992
rect 21039 16952 21088 16980
rect 21039 16949 21051 16952
rect 20993 16943 21051 16949
rect 21082 16940 21088 16952
rect 21140 16940 21146 16992
rect 23382 16980 23388 16992
rect 23343 16952 23388 16980
rect 23382 16940 23388 16952
rect 23440 16940 23446 16992
rect 25222 16980 25228 16992
rect 25183 16952 25228 16980
rect 25222 16940 25228 16952
rect 25280 16940 25286 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 3237 16779 3295 16785
rect 3237 16776 3249 16779
rect 2924 16748 3249 16776
rect 2924 16736 2930 16748
rect 3237 16745 3249 16748
rect 3283 16745 3295 16779
rect 3237 16739 3295 16745
rect 5074 16736 5080 16788
rect 5132 16776 5138 16788
rect 13262 16776 13268 16788
rect 5132 16748 6592 16776
rect 13223 16748 13268 16776
rect 5132 16736 5138 16748
rect 3421 16711 3479 16717
rect 3421 16677 3433 16711
rect 3467 16708 3479 16711
rect 4614 16708 4620 16720
rect 3467 16680 4620 16708
rect 3467 16677 3479 16680
rect 3421 16671 3479 16677
rect 4614 16668 4620 16680
rect 4672 16668 4678 16720
rect 5074 16640 5080 16652
rect 5035 16612 5080 16640
rect 5074 16600 5080 16612
rect 5132 16600 5138 16652
rect 5350 16640 5356 16652
rect 5311 16612 5356 16640
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 6564 16572 6592 16748
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 21910 16776 21916 16788
rect 21008 16748 21916 16776
rect 21008 16649 21036 16748
rect 21910 16736 21916 16748
rect 21968 16736 21974 16788
rect 22002 16736 22008 16788
rect 22060 16776 22066 16788
rect 23385 16779 23443 16785
rect 22060 16736 22094 16776
rect 23385 16745 23397 16779
rect 23431 16776 23443 16779
rect 23934 16776 23940 16788
rect 23431 16748 23940 16776
rect 23431 16745 23443 16748
rect 23385 16739 23443 16745
rect 23934 16736 23940 16748
rect 23992 16736 23998 16788
rect 32858 16736 32864 16788
rect 32916 16776 32922 16788
rect 33045 16779 33103 16785
rect 33045 16776 33057 16779
rect 32916 16748 33057 16776
rect 32916 16736 32922 16748
rect 33045 16745 33057 16748
rect 33091 16745 33103 16779
rect 33045 16739 33103 16745
rect 33778 16736 33784 16788
rect 33836 16776 33842 16788
rect 36173 16779 36231 16785
rect 36173 16776 36185 16779
rect 33836 16748 36185 16776
rect 33836 16736 33842 16748
rect 36173 16745 36185 16748
rect 36219 16745 36231 16779
rect 36722 16776 36728 16788
rect 36683 16748 36728 16776
rect 36173 16739 36231 16745
rect 36722 16736 36728 16748
rect 36780 16736 36786 16788
rect 22066 16708 22094 16736
rect 28166 16708 28172 16720
rect 22066 16680 28172 16708
rect 28166 16668 28172 16680
rect 28224 16668 28230 16720
rect 20993 16643 21051 16649
rect 20993 16609 21005 16643
rect 21039 16609 21051 16643
rect 20993 16603 21051 16609
rect 22002 16600 22008 16652
rect 22060 16640 22066 16652
rect 26326 16640 26332 16652
rect 22060 16612 26332 16640
rect 22060 16600 22066 16612
rect 26326 16600 26332 16612
rect 26384 16600 26390 16652
rect 7377 16575 7435 16581
rect 7377 16572 7389 16575
rect 6564 16544 7389 16572
rect 7377 16541 7389 16544
rect 7423 16541 7435 16575
rect 13446 16572 13452 16584
rect 13407 16544 13452 16572
rect 7377 16535 7435 16541
rect 13446 16532 13452 16544
rect 13504 16532 13510 16584
rect 13630 16532 13636 16584
rect 13688 16572 13694 16584
rect 13725 16575 13783 16581
rect 13725 16572 13737 16575
rect 13688 16544 13737 16572
rect 13688 16532 13694 16544
rect 13725 16541 13737 16544
rect 13771 16541 13783 16575
rect 13725 16535 13783 16541
rect 17221 16575 17279 16581
rect 17221 16541 17233 16575
rect 17267 16541 17279 16575
rect 17402 16572 17408 16584
rect 17363 16544 17408 16572
rect 17221 16535 17279 16541
rect 2958 16464 2964 16516
rect 3016 16504 3022 16516
rect 3053 16507 3111 16513
rect 3053 16504 3065 16507
rect 3016 16476 3065 16504
rect 3016 16464 3022 16476
rect 3053 16473 3065 16476
rect 3099 16473 3111 16507
rect 3053 16467 3111 16473
rect 3269 16507 3327 16513
rect 3269 16473 3281 16507
rect 3315 16504 3327 16507
rect 4706 16504 4712 16516
rect 3315 16476 4712 16504
rect 3315 16473 3327 16476
rect 3269 16467 3327 16473
rect 4706 16464 4712 16476
rect 4764 16464 4770 16516
rect 5994 16464 6000 16516
rect 6052 16464 6058 16516
rect 7650 16504 7656 16516
rect 7611 16476 7656 16504
rect 7650 16464 7656 16476
rect 7708 16464 7714 16516
rect 16850 16504 16856 16516
rect 12406 16476 16856 16504
rect 6178 16396 6184 16448
rect 6236 16436 6242 16448
rect 6825 16439 6883 16445
rect 6825 16436 6837 16439
rect 6236 16408 6837 16436
rect 6236 16396 6242 16408
rect 6825 16405 6837 16408
rect 6871 16436 6883 16439
rect 12406 16436 12434 16476
rect 16850 16464 16856 16476
rect 16908 16464 16914 16516
rect 17236 16504 17264 16535
rect 17402 16532 17408 16544
rect 17460 16532 17466 16584
rect 17678 16572 17684 16584
rect 17591 16544 17684 16572
rect 17678 16532 17684 16544
rect 17736 16572 17742 16584
rect 20714 16572 20720 16584
rect 17736 16544 20720 16572
rect 17736 16532 17742 16544
rect 20714 16532 20720 16544
rect 20772 16572 20778 16584
rect 20898 16572 20904 16584
rect 20772 16544 20904 16572
rect 20772 16532 20778 16544
rect 20898 16532 20904 16544
rect 20956 16532 20962 16584
rect 21082 16532 21088 16584
rect 21140 16572 21146 16584
rect 21249 16575 21307 16581
rect 21249 16572 21261 16575
rect 21140 16544 21261 16572
rect 21140 16532 21146 16544
rect 21249 16541 21261 16544
rect 21295 16541 21307 16575
rect 21249 16535 21307 16541
rect 21818 16532 21824 16584
rect 21876 16572 21882 16584
rect 22020 16572 22048 16600
rect 23566 16572 23572 16584
rect 21876 16544 22048 16572
rect 23527 16544 23572 16572
rect 21876 16532 21882 16544
rect 23566 16532 23572 16544
rect 23624 16532 23630 16584
rect 23658 16532 23664 16584
rect 23716 16572 23722 16584
rect 23845 16575 23903 16581
rect 23845 16572 23857 16575
rect 23716 16544 23857 16572
rect 23716 16532 23722 16544
rect 23845 16541 23857 16544
rect 23891 16541 23903 16575
rect 23845 16535 23903 16541
rect 25961 16575 26019 16581
rect 25961 16541 25973 16575
rect 26007 16572 26019 16575
rect 26142 16572 26148 16584
rect 26007 16544 26148 16572
rect 26007 16541 26019 16544
rect 25961 16535 26019 16541
rect 26142 16532 26148 16544
rect 26200 16532 26206 16584
rect 26237 16575 26295 16581
rect 26237 16541 26249 16575
rect 26283 16541 26295 16575
rect 26237 16535 26295 16541
rect 17954 16504 17960 16516
rect 17236 16476 17960 16504
rect 17954 16464 17960 16476
rect 18012 16504 18018 16516
rect 18598 16504 18604 16516
rect 18012 16476 18604 16504
rect 18012 16464 18018 16476
rect 18598 16464 18604 16476
rect 18656 16464 18662 16516
rect 23753 16507 23811 16513
rect 23753 16473 23765 16507
rect 23799 16504 23811 16507
rect 24854 16504 24860 16516
rect 23799 16476 24860 16504
rect 23799 16473 23811 16476
rect 23753 16467 23811 16473
rect 24854 16464 24860 16476
rect 24912 16504 24918 16516
rect 25222 16504 25228 16516
rect 24912 16476 25228 16504
rect 24912 16464 24918 16476
rect 25222 16464 25228 16476
rect 25280 16464 25286 16516
rect 26050 16464 26056 16516
rect 26108 16504 26114 16516
rect 26252 16504 26280 16535
rect 29454 16532 29460 16584
rect 29512 16572 29518 16584
rect 29733 16575 29791 16581
rect 29733 16572 29745 16575
rect 29512 16544 29745 16572
rect 29512 16532 29518 16544
rect 29733 16541 29745 16544
rect 29779 16541 29791 16575
rect 33226 16572 33232 16584
rect 33187 16544 33232 16572
rect 29733 16535 29791 16541
rect 33226 16532 33232 16544
rect 33284 16532 33290 16584
rect 33502 16572 33508 16584
rect 33415 16544 33508 16572
rect 33502 16532 33508 16544
rect 33560 16572 33566 16584
rect 34330 16572 34336 16584
rect 33560 16544 34336 16572
rect 33560 16532 33566 16544
rect 34330 16532 34336 16544
rect 34388 16532 34394 16584
rect 36081 16575 36139 16581
rect 36081 16541 36093 16575
rect 36127 16572 36139 16575
rect 36127 16544 36860 16572
rect 36127 16541 36139 16544
rect 36081 16535 36139 16541
rect 26108 16476 26280 16504
rect 26108 16464 26114 16476
rect 28534 16464 28540 16516
rect 28592 16504 28598 16516
rect 29978 16507 30036 16513
rect 29978 16504 29990 16507
rect 28592 16476 29990 16504
rect 28592 16464 28598 16476
rect 29978 16473 29990 16476
rect 30024 16473 30036 16507
rect 35894 16504 35900 16516
rect 35855 16476 35900 16504
rect 29978 16467 30036 16473
rect 35894 16464 35900 16476
rect 35952 16464 35958 16516
rect 36832 16504 36860 16544
rect 36906 16532 36912 16584
rect 36964 16572 36970 16584
rect 37093 16575 37151 16581
rect 36964 16544 37009 16572
rect 36964 16532 36970 16544
rect 37093 16541 37105 16575
rect 37139 16541 37151 16575
rect 37093 16535 37151 16541
rect 37108 16504 37136 16535
rect 37182 16532 37188 16584
rect 37240 16572 37246 16584
rect 37240 16544 37285 16572
rect 37240 16532 37246 16544
rect 37826 16504 37832 16516
rect 36832 16476 37832 16504
rect 37826 16464 37832 16476
rect 37884 16464 37890 16516
rect 6871 16408 12434 16436
rect 13633 16439 13691 16445
rect 6871 16405 6883 16408
rect 6825 16399 6883 16405
rect 13633 16405 13645 16439
rect 13679 16436 13691 16439
rect 14090 16436 14096 16448
rect 13679 16408 14096 16436
rect 13679 16405 13691 16408
rect 13633 16399 13691 16405
rect 14090 16396 14096 16408
rect 14148 16436 14154 16448
rect 14642 16436 14648 16448
rect 14148 16408 14648 16436
rect 14148 16396 14154 16408
rect 14642 16396 14648 16408
rect 14700 16396 14706 16448
rect 22370 16436 22376 16448
rect 22331 16408 22376 16436
rect 22370 16396 22376 16408
rect 22428 16396 22434 16448
rect 25774 16436 25780 16448
rect 25735 16408 25780 16436
rect 25774 16396 25780 16408
rect 25832 16396 25838 16448
rect 26142 16436 26148 16448
rect 26103 16408 26148 16436
rect 26142 16396 26148 16408
rect 26200 16396 26206 16448
rect 30926 16396 30932 16448
rect 30984 16436 30990 16448
rect 31113 16439 31171 16445
rect 31113 16436 31125 16439
rect 30984 16408 31125 16436
rect 30984 16396 30990 16408
rect 31113 16405 31125 16408
rect 31159 16405 31171 16439
rect 33410 16436 33416 16448
rect 33371 16408 33416 16436
rect 31113 16399 31171 16405
rect 33410 16396 33416 16408
rect 33468 16396 33474 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 5074 16192 5080 16244
rect 5132 16232 5138 16244
rect 9122 16232 9128 16244
rect 5132 16204 9128 16232
rect 5132 16192 5138 16204
rect 3234 16124 3240 16176
rect 3292 16164 3298 16176
rect 5994 16164 6000 16176
rect 3292 16136 5764 16164
rect 5955 16136 6000 16164
rect 3292 16124 3298 16136
rect 5534 16056 5540 16108
rect 5592 16096 5598 16108
rect 5629 16099 5687 16105
rect 5629 16096 5641 16099
rect 5592 16068 5641 16096
rect 5592 16056 5598 16068
rect 5629 16065 5641 16068
rect 5675 16065 5687 16099
rect 5736 16096 5764 16136
rect 5994 16124 6000 16136
rect 6052 16124 6058 16176
rect 6656 16164 6684 16204
rect 9122 16192 9128 16204
rect 9180 16192 9186 16244
rect 13354 16232 13360 16244
rect 13315 16204 13360 16232
rect 13354 16192 13360 16204
rect 13412 16192 13418 16244
rect 15010 16232 15016 16244
rect 13556 16204 15016 16232
rect 6822 16164 6828 16176
rect 6564 16136 6684 16164
rect 6783 16136 6828 16164
rect 5902 16096 5908 16108
rect 5736 16068 5908 16096
rect 5629 16059 5687 16065
rect 5902 16056 5908 16068
rect 5960 16056 5966 16108
rect 6564 16105 6592 16136
rect 6822 16124 6828 16136
rect 6880 16124 6886 16176
rect 7282 16124 7288 16176
rect 7340 16124 7346 16176
rect 9950 16124 9956 16176
rect 10008 16124 10014 16176
rect 6549 16099 6607 16105
rect 6549 16065 6561 16099
rect 6595 16065 6607 16099
rect 6549 16059 6607 16065
rect 9122 16056 9128 16108
rect 9180 16096 9186 16108
rect 13556 16105 13584 16204
rect 15010 16192 15016 16204
rect 15068 16192 15074 16244
rect 15194 16232 15200 16244
rect 15155 16204 15200 16232
rect 15194 16192 15200 16204
rect 15252 16192 15258 16244
rect 20809 16235 20867 16241
rect 20809 16201 20821 16235
rect 20855 16232 20867 16235
rect 21266 16232 21272 16244
rect 20855 16204 21272 16232
rect 20855 16201 20867 16204
rect 20809 16195 20867 16201
rect 21266 16192 21272 16204
rect 21324 16192 21330 16244
rect 28534 16232 28540 16244
rect 28495 16204 28540 16232
rect 28534 16192 28540 16204
rect 28592 16192 28598 16244
rect 35894 16232 35900 16244
rect 35855 16204 35900 16232
rect 35894 16192 35900 16204
rect 35952 16192 35958 16244
rect 36817 16235 36875 16241
rect 36817 16201 36829 16235
rect 36863 16232 36875 16235
rect 37182 16232 37188 16244
rect 36863 16204 37188 16232
rect 36863 16201 36875 16204
rect 36817 16195 36875 16201
rect 37182 16192 37188 16204
rect 37240 16192 37246 16244
rect 37826 16232 37832 16244
rect 37787 16204 37832 16232
rect 37826 16192 37832 16204
rect 37884 16192 37890 16244
rect 13630 16124 13636 16176
rect 13688 16164 13694 16176
rect 14826 16164 14832 16176
rect 13688 16136 13860 16164
rect 14739 16136 14832 16164
rect 13688 16124 13694 16136
rect 9217 16099 9275 16105
rect 9217 16096 9229 16099
rect 9180 16068 9229 16096
rect 9180 16056 9186 16068
rect 9217 16065 9229 16068
rect 9263 16065 9275 16099
rect 9217 16059 9275 16065
rect 13541 16099 13599 16105
rect 13541 16065 13553 16099
rect 13587 16065 13599 16099
rect 13722 16096 13728 16108
rect 13683 16068 13728 16096
rect 13541 16059 13599 16065
rect 13722 16056 13728 16068
rect 13780 16056 13786 16108
rect 13832 16105 13860 16136
rect 14826 16124 14832 16136
rect 14884 16164 14890 16176
rect 16666 16164 16672 16176
rect 14884 16136 16672 16164
rect 14884 16124 14890 16136
rect 16666 16124 16672 16136
rect 16724 16164 16730 16176
rect 17678 16164 17684 16176
rect 16724 16136 17684 16164
rect 16724 16124 16730 16136
rect 17678 16124 17684 16136
rect 17736 16124 17742 16176
rect 23382 16164 23388 16176
rect 21100 16136 23388 16164
rect 13817 16099 13875 16105
rect 13817 16065 13829 16099
rect 13863 16065 13875 16099
rect 13817 16059 13875 16065
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 5442 15988 5448 16040
rect 5500 16028 5506 16040
rect 6822 16028 6828 16040
rect 5500 16000 6828 16028
rect 5500 15988 5506 16000
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 9490 16028 9496 16040
rect 9451 16000 9496 16028
rect 9490 15988 9496 16000
rect 9548 15988 9554 16040
rect 14568 16028 14596 16059
rect 14642 16056 14648 16108
rect 14700 16096 14706 16108
rect 14700 16068 14745 16096
rect 14700 16056 14706 16068
rect 14918 16056 14924 16108
rect 14976 16096 14982 16108
rect 15059 16099 15117 16105
rect 14976 16068 15021 16096
rect 14976 16056 14982 16068
rect 15059 16065 15071 16099
rect 15105 16096 15117 16099
rect 16022 16096 16028 16108
rect 15105 16068 16028 16096
rect 15105 16065 15117 16068
rect 15059 16059 15117 16065
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 16850 16096 16856 16108
rect 16811 16068 16856 16096
rect 16850 16056 16856 16068
rect 16908 16056 16914 16108
rect 17218 16096 17224 16108
rect 17179 16068 17224 16096
rect 17218 16056 17224 16068
rect 17276 16056 17282 16108
rect 17310 16056 17316 16108
rect 17368 16096 17374 16108
rect 17405 16099 17463 16105
rect 17405 16096 17417 16099
rect 17368 16068 17417 16096
rect 17368 16056 17374 16068
rect 17405 16065 17417 16068
rect 17451 16065 17463 16099
rect 17405 16059 17463 16065
rect 17862 16056 17868 16108
rect 17920 16096 17926 16108
rect 18049 16099 18107 16105
rect 18049 16096 18061 16099
rect 17920 16068 18061 16096
rect 17920 16056 17926 16068
rect 18049 16065 18061 16068
rect 18095 16065 18107 16099
rect 18049 16059 18107 16065
rect 18417 16099 18475 16105
rect 18417 16065 18429 16099
rect 18463 16096 18475 16099
rect 18506 16096 18512 16108
rect 18463 16068 18512 16096
rect 18463 16065 18475 16068
rect 18417 16059 18475 16065
rect 18506 16056 18512 16068
rect 18564 16056 18570 16108
rect 21100 16105 21128 16136
rect 23382 16124 23388 16136
rect 23440 16124 23446 16176
rect 25492 16167 25550 16173
rect 25492 16133 25504 16167
rect 25538 16164 25550 16167
rect 25774 16164 25780 16176
rect 25538 16136 25780 16164
rect 25538 16133 25550 16136
rect 25492 16127 25550 16133
rect 25774 16124 25780 16136
rect 25832 16124 25838 16176
rect 28905 16167 28963 16173
rect 28905 16133 28917 16167
rect 28951 16164 28963 16167
rect 30926 16164 30932 16176
rect 28951 16136 30932 16164
rect 28951 16133 28963 16136
rect 28905 16127 28963 16133
rect 30926 16124 30932 16136
rect 30984 16124 30990 16176
rect 37366 16164 37372 16176
rect 35820 16136 37372 16164
rect 18601 16099 18659 16105
rect 18601 16065 18613 16099
rect 18647 16065 18659 16099
rect 18601 16059 18659 16065
rect 20993 16099 21051 16105
rect 20993 16065 21005 16099
rect 21039 16065 21051 16099
rect 20993 16059 21051 16065
rect 21085 16099 21143 16105
rect 21085 16065 21097 16099
rect 21131 16065 21143 16099
rect 21266 16096 21272 16108
rect 21227 16068 21272 16096
rect 21085 16059 21143 16065
rect 16390 16028 16396 16040
rect 14568 16000 16396 16028
rect 16390 15988 16396 16000
rect 16448 15988 16454 16040
rect 18616 16028 18644 16059
rect 16868 16000 18644 16028
rect 21008 16028 21036 16059
rect 21266 16056 21272 16068
rect 21324 16056 21330 16108
rect 21358 16056 21364 16108
rect 21416 16096 21422 16108
rect 28721 16099 28779 16105
rect 21416 16068 21461 16096
rect 21416 16056 21422 16068
rect 28721 16065 28733 16099
rect 28767 16065 28779 16099
rect 28721 16059 28779 16065
rect 22186 16028 22192 16040
rect 21008 16000 22192 16028
rect 16868 15972 16896 16000
rect 22186 15988 22192 16000
rect 22244 15988 22250 16040
rect 24670 15988 24676 16040
rect 24728 16028 24734 16040
rect 25225 16031 25283 16037
rect 25225 16028 25237 16031
rect 24728 16000 25237 16028
rect 24728 15988 24734 16000
rect 25225 15997 25237 16000
rect 25271 15997 25283 16031
rect 28736 16028 28764 16059
rect 28994 16056 29000 16108
rect 29052 16096 29058 16108
rect 29724 16099 29782 16105
rect 29052 16068 29097 16096
rect 29052 16056 29058 16068
rect 29724 16065 29736 16099
rect 29770 16096 29782 16099
rect 30650 16096 30656 16108
rect 29770 16068 30656 16096
rect 29770 16065 29782 16068
rect 29724 16059 29782 16065
rect 30650 16056 30656 16068
rect 30708 16056 30714 16108
rect 35820 16105 35848 16136
rect 37366 16124 37372 16136
rect 37424 16164 37430 16176
rect 37424 16136 37688 16164
rect 37424 16124 37430 16136
rect 35805 16099 35863 16105
rect 35805 16065 35817 16099
rect 35851 16065 35863 16099
rect 35805 16059 35863 16065
rect 35989 16099 36047 16105
rect 35989 16065 36001 16099
rect 36035 16096 36047 16099
rect 36354 16096 36360 16108
rect 36035 16068 36360 16096
rect 36035 16065 36047 16068
rect 35989 16059 36047 16065
rect 36354 16056 36360 16068
rect 36412 16096 36418 16108
rect 36412 16068 36584 16096
rect 36412 16056 36418 16068
rect 29086 16028 29092 16040
rect 28736 16000 29092 16028
rect 25225 15991 25283 15997
rect 29086 15988 29092 16000
rect 29144 15988 29150 16040
rect 29454 16028 29460 16040
rect 29415 16000 29460 16028
rect 29454 15988 29460 16000
rect 29512 15988 29518 16040
rect 36446 16028 36452 16040
rect 36407 16000 36452 16028
rect 36446 15988 36452 16000
rect 36504 15988 36510 16040
rect 36556 16028 36584 16068
rect 36630 16056 36636 16108
rect 36688 16096 36694 16108
rect 37660 16105 37688 16136
rect 37645 16099 37703 16105
rect 36688 16068 36733 16096
rect 36688 16056 36694 16068
rect 37645 16065 37657 16099
rect 37691 16065 37703 16099
rect 37645 16059 37703 16065
rect 37461 16031 37519 16037
rect 37461 16028 37473 16031
rect 36556 16000 37473 16028
rect 37461 15997 37473 16000
rect 37507 15997 37519 16031
rect 37461 15991 37519 15997
rect 16850 15920 16856 15972
rect 16908 15920 16914 15972
rect 35894 15920 35900 15972
rect 35952 15960 35958 15972
rect 36630 15960 36636 15972
rect 35952 15932 36636 15960
rect 35952 15920 35958 15932
rect 36630 15920 36636 15932
rect 36688 15920 36694 15972
rect 8202 15852 8208 15904
rect 8260 15892 8266 15904
rect 8297 15895 8355 15901
rect 8297 15892 8309 15895
rect 8260 15864 8309 15892
rect 8260 15852 8266 15864
rect 8297 15861 8309 15864
rect 8343 15861 8355 15895
rect 8297 15855 8355 15861
rect 10502 15852 10508 15904
rect 10560 15892 10566 15904
rect 10965 15895 11023 15901
rect 10965 15892 10977 15895
rect 10560 15864 10977 15892
rect 10560 15852 10566 15864
rect 10965 15861 10977 15864
rect 11011 15861 11023 15895
rect 10965 15855 11023 15861
rect 25038 15852 25044 15904
rect 25096 15892 25102 15904
rect 26142 15892 26148 15904
rect 25096 15864 26148 15892
rect 25096 15852 25102 15864
rect 26142 15852 26148 15864
rect 26200 15892 26206 15904
rect 26605 15895 26663 15901
rect 26605 15892 26617 15895
rect 26200 15864 26617 15892
rect 26200 15852 26206 15864
rect 26605 15861 26617 15864
rect 26651 15861 26663 15895
rect 26605 15855 26663 15861
rect 30837 15895 30895 15901
rect 30837 15861 30849 15895
rect 30883 15892 30895 15895
rect 31202 15892 31208 15904
rect 30883 15864 31208 15892
rect 30883 15861 30895 15864
rect 30837 15855 30895 15861
rect 31202 15852 31208 15864
rect 31260 15852 31266 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 30650 15688 30656 15700
rect 30611 15660 30656 15688
rect 30650 15648 30656 15660
rect 30708 15648 30714 15700
rect 33410 15648 33416 15700
rect 33468 15688 33474 15700
rect 34241 15691 34299 15697
rect 34241 15688 34253 15691
rect 33468 15660 34253 15688
rect 33468 15648 33474 15660
rect 34241 15657 34253 15660
rect 34287 15657 34299 15691
rect 34241 15651 34299 15657
rect 34330 15648 34336 15700
rect 34388 15688 34394 15700
rect 35253 15691 35311 15697
rect 35253 15688 35265 15691
rect 34388 15660 35265 15688
rect 34388 15648 34394 15660
rect 35253 15657 35265 15660
rect 35299 15657 35311 15691
rect 37366 15688 37372 15700
rect 37327 15660 37372 15688
rect 35253 15651 35311 15657
rect 37366 15648 37372 15660
rect 37424 15648 37430 15700
rect 8202 15580 8208 15632
rect 8260 15620 8266 15632
rect 36817 15623 36875 15629
rect 8260 15592 16574 15620
rect 8260 15580 8266 15592
rect 7193 15555 7251 15561
rect 7193 15521 7205 15555
rect 7239 15552 7251 15555
rect 7282 15552 7288 15564
rect 7239 15524 7288 15552
rect 7239 15521 7251 15524
rect 7193 15515 7251 15521
rect 7282 15512 7288 15524
rect 7340 15512 7346 15564
rect 9950 15552 9956 15564
rect 8128 15524 9812 15552
rect 9911 15524 9956 15552
rect 5534 15444 5540 15496
rect 5592 15484 5598 15496
rect 6825 15487 6883 15493
rect 6825 15484 6837 15487
rect 5592 15456 6837 15484
rect 5592 15444 5598 15456
rect 6825 15453 6837 15456
rect 6871 15453 6883 15487
rect 6825 15447 6883 15453
rect 7101 15487 7159 15493
rect 7101 15453 7113 15487
rect 7147 15484 7159 15487
rect 7650 15484 7656 15496
rect 7147 15456 7656 15484
rect 7147 15453 7159 15456
rect 7101 15447 7159 15453
rect 6840 15416 6868 15447
rect 7650 15444 7656 15456
rect 7708 15484 7714 15496
rect 8128 15484 8156 15524
rect 9784 15496 9812 15524
rect 9950 15512 9956 15524
rect 10008 15512 10014 15564
rect 12158 15552 12164 15564
rect 12119 15524 12164 15552
rect 12158 15512 12164 15524
rect 12216 15512 12222 15564
rect 7708 15456 8156 15484
rect 9677 15487 9735 15493
rect 7708 15444 7714 15456
rect 9677 15453 9689 15487
rect 9723 15453 9735 15487
rect 9677 15447 9735 15453
rect 9692 15416 9720 15447
rect 9766 15444 9772 15496
rect 9824 15484 9830 15496
rect 10413 15487 10471 15493
rect 9824 15456 9869 15484
rect 9824 15444 9830 15456
rect 10413 15453 10425 15487
rect 10459 15484 10471 15487
rect 13998 15484 14004 15496
rect 10459 15456 14004 15484
rect 10459 15453 10471 15456
rect 10413 15447 10471 15453
rect 13998 15444 14004 15456
rect 14056 15444 14062 15496
rect 16393 15487 16451 15493
rect 16393 15453 16405 15487
rect 16439 15453 16451 15487
rect 16546 15484 16574 15592
rect 36817 15589 36829 15623
rect 36863 15620 36875 15623
rect 36906 15620 36912 15632
rect 36863 15592 36912 15620
rect 36863 15589 36875 15592
rect 36817 15583 36875 15589
rect 36906 15580 36912 15592
rect 36964 15580 36970 15632
rect 16666 15552 16672 15564
rect 16627 15524 16672 15552
rect 16666 15512 16672 15524
rect 16724 15552 16730 15564
rect 17586 15552 17592 15564
rect 16724 15524 17592 15552
rect 16724 15512 16730 15524
rect 17586 15512 17592 15524
rect 17644 15552 17650 15564
rect 18141 15555 18199 15561
rect 17644 15524 17816 15552
rect 17644 15512 17650 15524
rect 16850 15484 16856 15496
rect 16546 15456 16856 15484
rect 16393 15447 16451 15453
rect 6840 15388 9720 15416
rect 10502 15376 10508 15428
rect 10560 15416 10566 15428
rect 16408 15416 16436 15447
rect 16850 15444 16856 15456
rect 16908 15484 16914 15496
rect 17788 15493 17816 15524
rect 18141 15521 18153 15555
rect 18187 15552 18199 15555
rect 18690 15552 18696 15564
rect 18187 15524 18696 15552
rect 18187 15521 18199 15524
rect 18141 15515 18199 15521
rect 18690 15512 18696 15524
rect 18748 15512 18754 15564
rect 24670 15512 24676 15564
rect 24728 15552 24734 15564
rect 25777 15555 25835 15561
rect 25777 15552 25789 15555
rect 24728 15524 25789 15552
rect 24728 15512 24734 15524
rect 25777 15521 25789 15524
rect 25823 15521 25835 15555
rect 25777 15515 25835 15521
rect 28994 15512 29000 15564
rect 29052 15552 29058 15564
rect 29917 15555 29975 15561
rect 29917 15552 29929 15555
rect 29052 15524 29929 15552
rect 29052 15512 29058 15524
rect 29917 15521 29929 15524
rect 29963 15552 29975 15555
rect 30190 15552 30196 15564
rect 29963 15524 30196 15552
rect 29963 15521 29975 15524
rect 29917 15515 29975 15521
rect 30190 15512 30196 15524
rect 30248 15552 30254 15564
rect 34882 15552 34888 15564
rect 30248 15524 31156 15552
rect 30248 15512 30254 15524
rect 17037 15487 17095 15493
rect 17037 15484 17049 15487
rect 16908 15456 17049 15484
rect 16908 15444 16914 15456
rect 17037 15453 17049 15456
rect 17083 15453 17095 15487
rect 17037 15447 17095 15453
rect 17773 15487 17831 15493
rect 17773 15453 17785 15487
rect 17819 15453 17831 15487
rect 17773 15447 17831 15453
rect 18049 15487 18107 15493
rect 18049 15453 18061 15487
rect 18095 15484 18107 15487
rect 19150 15484 19156 15496
rect 18095 15456 19156 15484
rect 18095 15453 18107 15456
rect 18049 15447 18107 15453
rect 19150 15444 19156 15456
rect 19208 15444 19214 15496
rect 19242 15444 19248 15496
rect 19300 15484 19306 15496
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 19300 15456 19441 15484
rect 19300 15444 19306 15456
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 19613 15487 19671 15493
rect 19613 15453 19625 15487
rect 19659 15453 19671 15487
rect 19613 15447 19671 15453
rect 24765 15487 24823 15493
rect 24765 15453 24777 15487
rect 24811 15484 24823 15487
rect 24854 15484 24860 15496
rect 24811 15456 24860 15484
rect 24811 15453 24823 15456
rect 24765 15447 24823 15453
rect 16758 15416 16764 15428
rect 10560 15388 16764 15416
rect 10560 15376 10566 15388
rect 16758 15376 16764 15388
rect 16816 15376 16822 15428
rect 19168 15416 19196 15444
rect 19628 15416 19656 15447
rect 24854 15444 24860 15456
rect 24912 15444 24918 15496
rect 25038 15484 25044 15496
rect 24999 15456 25044 15484
rect 25038 15444 25044 15456
rect 25096 15444 25102 15496
rect 25130 15444 25136 15496
rect 25188 15484 25194 15496
rect 25188 15456 25233 15484
rect 25188 15444 25194 15456
rect 29546 15444 29552 15496
rect 29604 15484 29610 15496
rect 31128 15493 31156 15524
rect 34348 15524 34888 15552
rect 29733 15487 29791 15493
rect 29733 15484 29745 15487
rect 29604 15456 29745 15484
rect 29604 15444 29610 15456
rect 29733 15453 29745 15456
rect 29779 15453 29791 15487
rect 29733 15447 29791 15453
rect 30837 15487 30895 15493
rect 30837 15453 30849 15487
rect 30883 15453 30895 15487
rect 30837 15447 30895 15453
rect 31113 15487 31171 15493
rect 31113 15453 31125 15487
rect 31159 15453 31171 15487
rect 31113 15447 31171 15453
rect 19168 15388 19656 15416
rect 19797 15419 19855 15425
rect 19797 15385 19809 15419
rect 19843 15416 19855 15419
rect 20254 15416 20260 15428
rect 19843 15388 20260 15416
rect 19843 15385 19855 15388
rect 19797 15379 19855 15385
rect 20254 15376 20260 15388
rect 20312 15416 20318 15428
rect 22186 15416 22192 15428
rect 20312 15388 22192 15416
rect 20312 15376 20318 15388
rect 22186 15376 22192 15388
rect 22244 15416 22250 15428
rect 24949 15419 25007 15425
rect 24949 15416 24961 15419
rect 22244 15388 24961 15416
rect 22244 15376 22250 15388
rect 24949 15385 24961 15388
rect 24995 15385 25007 15419
rect 24949 15379 25007 15385
rect 26044 15419 26102 15425
rect 26044 15385 26056 15419
rect 26090 15416 26102 15419
rect 26142 15416 26148 15428
rect 26090 15388 26148 15416
rect 26090 15385 26102 15388
rect 26044 15379 26102 15385
rect 26142 15376 26148 15388
rect 26200 15376 26206 15428
rect 30852 15416 30880 15447
rect 33686 15444 33692 15496
rect 33744 15484 33750 15496
rect 34348 15493 34376 15524
rect 34882 15512 34888 15524
rect 34940 15512 34946 15564
rect 36354 15552 36360 15564
rect 36315 15524 36360 15552
rect 36354 15512 36360 15524
rect 36412 15512 36418 15564
rect 34149 15487 34207 15493
rect 34149 15484 34161 15487
rect 33744 15456 34161 15484
rect 33744 15444 33750 15456
rect 34149 15453 34161 15456
rect 34195 15453 34207 15487
rect 34149 15447 34207 15453
rect 34333 15487 34391 15493
rect 34333 15453 34345 15487
rect 34379 15453 34391 15487
rect 34333 15447 34391 15453
rect 31386 15416 31392 15428
rect 30852 15388 31392 15416
rect 31386 15376 31392 15388
rect 31444 15376 31450 15428
rect 13446 15308 13452 15360
rect 13504 15348 13510 15360
rect 17034 15348 17040 15360
rect 13504 15320 17040 15348
rect 13504 15308 13510 15320
rect 17034 15308 17040 15320
rect 17092 15308 17098 15360
rect 25317 15351 25375 15357
rect 25317 15317 25329 15351
rect 25363 15348 25375 15351
rect 25866 15348 25872 15360
rect 25363 15320 25872 15348
rect 25363 15317 25375 15320
rect 25317 15311 25375 15317
rect 25866 15308 25872 15320
rect 25924 15308 25930 15360
rect 26510 15308 26516 15360
rect 26568 15348 26574 15360
rect 27157 15351 27215 15357
rect 27157 15348 27169 15351
rect 26568 15320 27169 15348
rect 26568 15308 26574 15320
rect 27157 15317 27169 15320
rect 27203 15317 27215 15351
rect 27157 15311 27215 15317
rect 31021 15351 31079 15357
rect 31021 15317 31033 15351
rect 31067 15348 31079 15351
rect 31202 15348 31208 15360
rect 31067 15320 31208 15348
rect 31067 15317 31079 15320
rect 31021 15311 31079 15317
rect 31202 15308 31208 15320
rect 31260 15308 31266 15360
rect 34164 15348 34192 15447
rect 34698 15444 34704 15496
rect 34756 15484 34762 15496
rect 35069 15487 35127 15493
rect 35069 15484 35081 15487
rect 34756 15456 35081 15484
rect 34756 15444 34762 15456
rect 35069 15453 35081 15456
rect 35115 15484 35127 15487
rect 36372 15484 36400 15512
rect 36538 15484 36544 15496
rect 35115 15456 36400 15484
rect 36499 15456 36544 15484
rect 35115 15453 35127 15456
rect 35069 15447 35127 15453
rect 36538 15444 36544 15456
rect 36596 15444 36602 15496
rect 36906 15484 36912 15496
rect 36867 15456 36912 15484
rect 36906 15444 36912 15456
rect 36964 15444 36970 15496
rect 37182 15444 37188 15496
rect 37240 15484 37246 15496
rect 37369 15487 37427 15493
rect 37369 15484 37381 15487
rect 37240 15456 37381 15484
rect 37240 15444 37246 15456
rect 37369 15453 37381 15456
rect 37415 15453 37427 15487
rect 37369 15447 37427 15453
rect 37553 15487 37611 15493
rect 37553 15453 37565 15487
rect 37599 15453 37611 15487
rect 37553 15447 37611 15453
rect 34790 15376 34796 15428
rect 34848 15416 34854 15428
rect 34885 15419 34943 15425
rect 34885 15416 34897 15419
rect 34848 15388 34897 15416
rect 34848 15376 34854 15388
rect 34885 15385 34897 15388
rect 34931 15385 34943 15419
rect 36924 15416 36952 15444
rect 37568 15416 37596 15447
rect 36924 15388 37596 15416
rect 34885 15379 34943 15385
rect 35158 15348 35164 15360
rect 34164 15320 35164 15348
rect 35158 15308 35164 15320
rect 35216 15308 35222 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 2130 15104 2136 15156
rect 2188 15144 2194 15156
rect 2593 15147 2651 15153
rect 2593 15144 2605 15147
rect 2188 15116 2605 15144
rect 2188 15104 2194 15116
rect 2593 15113 2605 15116
rect 2639 15144 2651 15147
rect 2961 15147 3019 15153
rect 2961 15144 2973 15147
rect 2639 15116 2973 15144
rect 2639 15113 2651 15116
rect 2593 15107 2651 15113
rect 2961 15113 2973 15116
rect 3007 15113 3019 15147
rect 2961 15107 3019 15113
rect 3145 15147 3203 15153
rect 3145 15113 3157 15147
rect 3191 15144 3203 15147
rect 7098 15144 7104 15156
rect 3191 15116 7104 15144
rect 3191 15113 3203 15116
rect 3145 15107 3203 15113
rect 3896 15017 3924 15116
rect 7098 15104 7104 15116
rect 7156 15104 7162 15156
rect 21269 15147 21327 15153
rect 21269 15113 21281 15147
rect 21315 15144 21327 15147
rect 21358 15144 21364 15156
rect 21315 15116 21364 15144
rect 21315 15113 21327 15116
rect 21269 15107 21327 15113
rect 21358 15104 21364 15116
rect 21416 15104 21422 15156
rect 26142 15144 26148 15156
rect 26103 15116 26148 15144
rect 26142 15104 26148 15116
rect 26200 15104 26206 15156
rect 26510 15144 26516 15156
rect 26471 15116 26516 15144
rect 26510 15104 26516 15116
rect 26568 15104 26574 15156
rect 28166 15144 28172 15156
rect 28127 15116 28172 15144
rect 28166 15104 28172 15116
rect 28224 15104 28230 15156
rect 32766 15144 32772 15156
rect 31864 15116 32772 15144
rect 31864 15088 31892 15116
rect 32766 15104 32772 15116
rect 32824 15144 32830 15156
rect 33505 15147 33563 15153
rect 33505 15144 33517 15147
rect 32824 15116 33517 15144
rect 32824 15104 32830 15116
rect 33505 15113 33517 15116
rect 33551 15113 33563 15147
rect 34514 15144 34520 15156
rect 33505 15107 33563 15113
rect 33612 15116 34520 15144
rect 13722 15036 13728 15088
rect 13780 15076 13786 15088
rect 20898 15076 20904 15088
rect 13780 15048 20760 15076
rect 20859 15048 20904 15076
rect 13780 15036 13786 15048
rect 3237 15011 3295 15017
rect 3237 14977 3249 15011
rect 3283 15008 3295 15011
rect 3697 15011 3755 15017
rect 3697 15008 3709 15011
rect 3283 14980 3709 15008
rect 3283 14977 3295 14980
rect 3237 14971 3295 14977
rect 3697 14977 3709 14980
rect 3743 14977 3755 15011
rect 3697 14971 3755 14977
rect 3881 15011 3939 15017
rect 3881 14977 3893 15011
rect 3927 14977 3939 15011
rect 13906 15008 13912 15020
rect 13819 14980 13912 15008
rect 3881 14971 3939 14977
rect 2682 14900 2688 14952
rect 2740 14940 2746 14952
rect 2777 14943 2835 14949
rect 2777 14940 2789 14943
rect 2740 14912 2789 14940
rect 2740 14900 2746 14912
rect 2777 14909 2789 14912
rect 2823 14909 2835 14943
rect 2777 14903 2835 14909
rect 2869 14943 2927 14949
rect 2869 14909 2881 14943
rect 2915 14940 2927 14943
rect 3142 14940 3148 14952
rect 2915 14912 3148 14940
rect 2915 14909 2927 14912
rect 2869 14903 2927 14909
rect 3142 14900 3148 14912
rect 3200 14900 3206 14952
rect 3712 14940 3740 14971
rect 13906 14968 13912 14980
rect 13964 14968 13970 15020
rect 16850 15008 16856 15020
rect 16811 14980 16856 15008
rect 16850 14968 16856 14980
rect 16908 14968 16914 15020
rect 17497 15011 17555 15017
rect 17497 14977 17509 15011
rect 17543 15008 17555 15011
rect 17862 15008 17868 15020
rect 17543 14980 17868 15008
rect 17543 14977 17555 14980
rect 17497 14971 17555 14977
rect 4706 14940 4712 14952
rect 3712 14912 4712 14940
rect 4706 14900 4712 14912
rect 4764 14900 4770 14952
rect 3786 14804 3792 14816
rect 3747 14776 3792 14804
rect 3786 14764 3792 14776
rect 3844 14764 3850 14816
rect 13924 14804 13952 14968
rect 14182 14940 14188 14952
rect 14143 14912 14188 14940
rect 14182 14900 14188 14912
rect 14240 14900 14246 14952
rect 16758 14900 16764 14952
rect 16816 14940 16822 14952
rect 17512 14940 17540 14971
rect 17862 14968 17868 14980
rect 17920 14968 17926 15020
rect 18506 14968 18512 15020
rect 18564 15008 18570 15020
rect 18785 15011 18843 15017
rect 18785 15008 18797 15011
rect 18564 14980 18797 15008
rect 18564 14968 18570 14980
rect 18785 14977 18797 14980
rect 18831 14977 18843 15011
rect 18785 14971 18843 14977
rect 19150 14968 19156 15020
rect 19208 15008 19214 15020
rect 20732 15017 20760 15048
rect 20898 15036 20904 15048
rect 20956 15036 20962 15088
rect 20993 15079 21051 15085
rect 20993 15045 21005 15079
rect 21039 15076 21051 15079
rect 22278 15076 22284 15088
rect 21039 15048 22284 15076
rect 21039 15045 21051 15048
rect 20993 15039 21051 15045
rect 22278 15036 22284 15048
rect 22336 15036 22342 15088
rect 25314 15036 25320 15088
rect 25372 15076 25378 15088
rect 26050 15076 26056 15088
rect 25372 15048 26056 15076
rect 25372 15036 25378 15048
rect 26050 15036 26056 15048
rect 26108 15076 26114 15088
rect 30837 15079 30895 15085
rect 26108 15048 26648 15076
rect 26108 15036 26114 15048
rect 21174 15017 21180 15020
rect 19245 15011 19303 15017
rect 19245 15008 19257 15011
rect 19208 14980 19257 15008
rect 19208 14968 19214 14980
rect 19245 14977 19257 14980
rect 19291 14977 19303 15011
rect 19245 14971 19303 14977
rect 20632 15011 20690 15017
rect 20632 14977 20644 15011
rect 20678 14977 20690 15011
rect 20632 14971 20690 14977
rect 20718 15011 20776 15017
rect 20718 14977 20730 15011
rect 20764 14977 20776 15011
rect 21131 15011 21180 15017
rect 21131 15008 21143 15011
rect 21087 14980 21143 15008
rect 20718 14971 20776 14977
rect 21131 14977 21143 14980
rect 21177 14977 21180 15011
rect 21131 14971 21180 14977
rect 16816 14912 17540 14940
rect 17589 14943 17647 14949
rect 16816 14900 16822 14912
rect 17589 14909 17601 14943
rect 17635 14909 17647 14943
rect 17589 14903 17647 14909
rect 19521 14943 19579 14949
rect 19521 14909 19533 14943
rect 19567 14909 19579 14943
rect 19521 14903 19579 14909
rect 17604 14872 17632 14903
rect 19242 14872 19248 14884
rect 17604 14844 19248 14872
rect 19242 14832 19248 14844
rect 19300 14832 19306 14884
rect 19334 14804 19340 14816
rect 13924 14776 19340 14804
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 19536 14804 19564 14903
rect 20640 14872 20668 14971
rect 21174 14968 21180 14971
rect 21232 15008 21238 15020
rect 24118 15008 24124 15020
rect 21232 14980 24124 15008
rect 21232 14968 21238 14980
rect 24118 14968 24124 14980
rect 24176 14968 24182 15020
rect 26326 15008 26332 15020
rect 26287 14980 26332 15008
rect 26326 14968 26332 14980
rect 26384 14968 26390 15020
rect 26620 15017 26648 15048
rect 30837 15045 30849 15079
rect 30883 15076 30895 15079
rect 31846 15076 31852 15088
rect 30883 15048 31852 15076
rect 30883 15045 30895 15048
rect 30837 15039 30895 15045
rect 31846 15036 31852 15048
rect 31904 15036 31910 15088
rect 32692 15048 33548 15076
rect 26605 15011 26663 15017
rect 26605 14977 26617 15011
rect 26651 14977 26663 15011
rect 28442 15008 28448 15020
rect 28403 14980 28448 15008
rect 26605 14971 26663 14977
rect 28442 14968 28448 14980
rect 28500 14968 28506 15020
rect 28629 15011 28687 15017
rect 28629 14977 28641 15011
rect 28675 15008 28687 15011
rect 28718 15008 28724 15020
rect 28675 14980 28724 15008
rect 28675 14977 28687 14980
rect 28629 14971 28687 14977
rect 28718 14968 28724 14980
rect 28776 14968 28782 15020
rect 30558 15008 30564 15020
rect 30519 14980 30564 15008
rect 30558 14968 30564 14980
rect 30616 14968 30622 15020
rect 30745 15011 30803 15017
rect 30745 14977 30757 15011
rect 30791 14977 30803 15011
rect 30926 15008 30932 15020
rect 30887 14980 30932 15008
rect 30745 14971 30803 14977
rect 28353 14943 28411 14949
rect 28353 14909 28365 14943
rect 28399 14909 28411 14943
rect 28353 14903 28411 14909
rect 28537 14943 28595 14949
rect 28537 14909 28549 14943
rect 28583 14909 28595 14943
rect 30760 14940 30788 14971
rect 30926 14968 30932 14980
rect 30984 15008 30990 15020
rect 32692 15017 32720 15048
rect 33520 15020 33548 15048
rect 32677 15011 32735 15017
rect 30984 14980 31754 15008
rect 30984 14968 30990 14980
rect 31202 14940 31208 14952
rect 30760 14912 31208 14940
rect 28537 14903 28595 14909
rect 21082 14872 21088 14884
rect 20640 14844 21088 14872
rect 21082 14832 21088 14844
rect 21140 14832 21146 14884
rect 25130 14804 25136 14816
rect 19536 14776 25136 14804
rect 25130 14764 25136 14776
rect 25188 14804 25194 14816
rect 26418 14804 26424 14816
rect 25188 14776 26424 14804
rect 25188 14764 25194 14776
rect 26418 14764 26424 14776
rect 26476 14764 26482 14816
rect 28368 14804 28396 14903
rect 28552 14872 28580 14903
rect 31202 14900 31208 14912
rect 31260 14900 31266 14952
rect 31726 14940 31754 14980
rect 32677 14977 32689 15011
rect 32723 14977 32735 15011
rect 32677 14971 32735 14977
rect 33042 14968 33048 15020
rect 33100 15008 33106 15020
rect 33321 15011 33379 15017
rect 33321 15008 33333 15011
rect 33100 14980 33333 15008
rect 33100 14968 33106 14980
rect 33321 14977 33333 14980
rect 33367 14977 33379 15011
rect 33321 14971 33379 14977
rect 33502 14968 33508 15020
rect 33560 14968 33566 15020
rect 33612 15017 33640 15116
rect 34514 15104 34520 15116
rect 34572 15144 34578 15156
rect 34885 15147 34943 15153
rect 34885 15144 34897 15147
rect 34572 15116 34897 15144
rect 34572 15104 34578 15116
rect 34885 15113 34897 15116
rect 34931 15113 34943 15147
rect 34885 15107 34943 15113
rect 34977 15147 35035 15153
rect 34977 15113 34989 15147
rect 35023 15113 35035 15147
rect 34977 15107 35035 15113
rect 36817 15147 36875 15153
rect 36817 15113 36829 15147
rect 36863 15144 36875 15147
rect 36906 15144 36912 15156
rect 36863 15116 36912 15144
rect 36863 15113 36875 15116
rect 36817 15107 36875 15113
rect 34606 15036 34612 15088
rect 34664 15076 34670 15088
rect 34992 15076 35020 15107
rect 36906 15104 36912 15116
rect 36964 15104 36970 15156
rect 35158 15076 35164 15088
rect 34664 15048 35020 15076
rect 35119 15048 35164 15076
rect 34664 15036 34670 15048
rect 35158 15036 35164 15048
rect 35216 15036 35222 15088
rect 36449 15079 36507 15085
rect 36449 15076 36461 15079
rect 35268 15048 36461 15076
rect 33597 15011 33655 15017
rect 33597 14977 33609 15011
rect 33643 14977 33655 15011
rect 33597 14971 33655 14977
rect 33689 15011 33747 15017
rect 33689 14977 33701 15011
rect 33735 14977 33747 15011
rect 33689 14971 33747 14977
rect 34793 15011 34851 15017
rect 34793 14977 34805 15011
rect 34839 15008 34851 15011
rect 34882 15008 34888 15020
rect 34839 14980 34888 15008
rect 34839 14977 34851 14980
rect 34793 14971 34851 14977
rect 33612 14940 33640 14971
rect 31726 14912 33640 14940
rect 32769 14875 32827 14881
rect 32769 14872 32781 14875
rect 28552 14844 32781 14872
rect 32769 14841 32781 14844
rect 32815 14841 32827 14875
rect 33704 14872 33732 14971
rect 34882 14968 34888 14980
rect 34940 14968 34946 15020
rect 34609 14943 34667 14949
rect 34609 14909 34621 14943
rect 34655 14940 34667 14943
rect 34698 14940 34704 14952
rect 34655 14912 34704 14940
rect 34655 14909 34667 14912
rect 34609 14903 34667 14909
rect 34698 14900 34704 14912
rect 34756 14900 34762 14952
rect 32769 14835 32827 14841
rect 33612 14844 33732 14872
rect 33612 14816 33640 14844
rect 34514 14832 34520 14884
rect 34572 14872 34578 14884
rect 35268 14872 35296 15048
rect 36449 15045 36461 15048
rect 36495 15045 36507 15079
rect 36649 15079 36707 15085
rect 36649 15076 36661 15079
rect 36449 15039 36507 15045
rect 36556 15048 36661 15076
rect 35805 15011 35863 15017
rect 35805 14977 35817 15011
rect 35851 15008 35863 15011
rect 35894 15008 35900 15020
rect 35851 14980 35900 15008
rect 35851 14977 35863 14980
rect 35805 14971 35863 14977
rect 35894 14968 35900 14980
rect 35952 14968 35958 15020
rect 36556 15008 36584 15048
rect 36649 15045 36661 15048
rect 36695 15045 36707 15079
rect 36649 15039 36707 15045
rect 36004 14980 36584 15008
rect 35342 14900 35348 14952
rect 35400 14940 35406 14952
rect 35621 14943 35679 14949
rect 35621 14940 35633 14943
rect 35400 14912 35633 14940
rect 35400 14900 35406 14912
rect 35621 14909 35633 14912
rect 35667 14909 35679 14943
rect 35621 14903 35679 14909
rect 34572 14844 35296 14872
rect 34572 14832 34578 14844
rect 31113 14807 31171 14813
rect 31113 14804 31125 14807
rect 28368 14776 31125 14804
rect 31113 14773 31125 14776
rect 31159 14773 31171 14807
rect 31113 14767 31171 14773
rect 31202 14764 31208 14816
rect 31260 14804 31266 14816
rect 33594 14804 33600 14816
rect 31260 14776 33600 14804
rect 31260 14764 31266 14776
rect 33594 14764 33600 14776
rect 33652 14764 33658 14816
rect 33686 14764 33692 14816
rect 33744 14804 33750 14816
rect 33873 14807 33931 14813
rect 33873 14804 33885 14807
rect 33744 14776 33885 14804
rect 33744 14764 33750 14776
rect 33873 14773 33885 14776
rect 33919 14773 33931 14807
rect 33873 14767 33931 14773
rect 34882 14764 34888 14816
rect 34940 14804 34946 14816
rect 35802 14804 35808 14816
rect 34940 14776 35808 14804
rect 34940 14764 34946 14776
rect 35802 14764 35808 14776
rect 35860 14804 35866 14816
rect 36004 14813 36032 14980
rect 35989 14807 36047 14813
rect 35989 14804 36001 14807
rect 35860 14776 36001 14804
rect 35860 14764 35866 14776
rect 35989 14773 36001 14776
rect 36035 14773 36047 14807
rect 35989 14767 36047 14773
rect 36170 14764 36176 14816
rect 36228 14804 36234 14816
rect 36538 14804 36544 14816
rect 36228 14776 36544 14804
rect 36228 14764 36234 14776
rect 36538 14764 36544 14776
rect 36596 14804 36602 14816
rect 36633 14807 36691 14813
rect 36633 14804 36645 14807
rect 36596 14776 36645 14804
rect 36596 14764 36602 14776
rect 36633 14773 36645 14776
rect 36679 14773 36691 14807
rect 36633 14767 36691 14773
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 1670 14560 1676 14612
rect 1728 14600 1734 14612
rect 3050 14600 3056 14612
rect 1728 14572 3056 14600
rect 1728 14560 1734 14572
rect 3050 14560 3056 14572
rect 3108 14600 3114 14612
rect 3970 14600 3976 14612
rect 3108 14572 3976 14600
rect 3108 14560 3114 14572
rect 3970 14560 3976 14572
rect 4028 14560 4034 14612
rect 16390 14560 16396 14612
rect 16448 14600 16454 14612
rect 20625 14603 20683 14609
rect 20625 14600 20637 14603
rect 16448 14572 20637 14600
rect 16448 14560 16454 14572
rect 20625 14569 20637 14572
rect 20671 14569 20683 14603
rect 20625 14563 20683 14569
rect 26881 14603 26939 14609
rect 26881 14569 26893 14603
rect 26927 14600 26939 14603
rect 28718 14600 28724 14612
rect 26927 14572 28724 14600
rect 26927 14569 26939 14572
rect 26881 14563 26939 14569
rect 28718 14560 28724 14572
rect 28776 14560 28782 14612
rect 30558 14560 30564 14612
rect 30616 14600 30622 14612
rect 33042 14600 33048 14612
rect 30616 14572 33048 14600
rect 30616 14560 30622 14572
rect 33042 14560 33048 14572
rect 33100 14560 33106 14612
rect 34790 14560 34796 14612
rect 34848 14600 34854 14612
rect 34885 14603 34943 14609
rect 34885 14600 34897 14603
rect 34848 14572 34897 14600
rect 34848 14560 34854 14572
rect 34885 14569 34897 14572
rect 34931 14569 34943 14603
rect 34885 14563 34943 14569
rect 35897 14603 35955 14609
rect 35897 14569 35909 14603
rect 35943 14600 35955 14603
rect 37182 14600 37188 14612
rect 35943 14572 37188 14600
rect 35943 14569 35955 14572
rect 35897 14563 35955 14569
rect 37182 14560 37188 14572
rect 37240 14560 37246 14612
rect 19058 14532 19064 14544
rect 18892 14504 19064 14532
rect 3050 14464 3056 14476
rect 3011 14436 3056 14464
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 3142 14424 3148 14476
rect 3200 14464 3206 14476
rect 16666 14464 16672 14476
rect 3200 14436 3245 14464
rect 16040 14436 16672 14464
rect 3200 14424 3206 14436
rect 2130 14396 2136 14408
rect 2091 14368 2136 14396
rect 2130 14356 2136 14368
rect 2188 14356 2194 14408
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2774 14396 2780 14408
rect 2271 14368 2780 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2774 14356 2780 14368
rect 2832 14356 2838 14408
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14365 3019 14399
rect 2961 14359 3019 14365
rect 2976 14328 3004 14359
rect 3234 14356 3240 14408
rect 3292 14396 3298 14408
rect 13446 14396 13452 14408
rect 3292 14368 3337 14396
rect 13407 14368 13452 14396
rect 3292 14356 3298 14368
rect 13446 14356 13452 14368
rect 13504 14356 13510 14408
rect 13725 14399 13783 14405
rect 13725 14365 13737 14399
rect 13771 14396 13783 14399
rect 14182 14396 14188 14408
rect 13771 14368 14188 14396
rect 13771 14365 13783 14368
rect 13725 14359 13783 14365
rect 14182 14356 14188 14368
rect 14240 14396 14246 14408
rect 15470 14396 15476 14408
rect 14240 14368 15476 14396
rect 14240 14356 14246 14368
rect 15470 14356 15476 14368
rect 15528 14356 15534 14408
rect 16040 14405 16068 14436
rect 16666 14424 16672 14436
rect 16724 14424 16730 14476
rect 17313 14467 17371 14473
rect 17313 14433 17325 14467
rect 17359 14464 17371 14467
rect 17954 14464 17960 14476
rect 17359 14436 17960 14464
rect 17359 14433 17371 14436
rect 17313 14427 17371 14433
rect 17954 14424 17960 14436
rect 18012 14424 18018 14476
rect 18506 14464 18512 14476
rect 18432 14436 18512 14464
rect 16025 14399 16083 14405
rect 16025 14365 16037 14399
rect 16071 14365 16083 14399
rect 16206 14396 16212 14408
rect 16167 14368 16212 14396
rect 16025 14359 16083 14365
rect 16206 14356 16212 14368
rect 16264 14356 16270 14408
rect 16758 14396 16764 14408
rect 16719 14368 16764 14396
rect 16758 14356 16764 14368
rect 16816 14356 16822 14408
rect 16850 14356 16856 14408
rect 16908 14396 16914 14408
rect 18432 14405 18460 14436
rect 18506 14424 18512 14436
rect 18564 14424 18570 14476
rect 18892 14473 18920 14504
rect 19058 14492 19064 14504
rect 19116 14532 19122 14544
rect 21174 14532 21180 14544
rect 19116 14504 21180 14532
rect 19116 14492 19122 14504
rect 21174 14492 21180 14504
rect 21232 14492 21238 14544
rect 24118 14492 24124 14544
rect 24176 14532 24182 14544
rect 24176 14504 26648 14532
rect 24176 14492 24182 14504
rect 18877 14467 18935 14473
rect 18877 14433 18889 14467
rect 18923 14433 18935 14467
rect 22370 14464 22376 14476
rect 18877 14427 18935 14433
rect 20088 14436 22376 14464
rect 16945 14399 17003 14405
rect 16945 14396 16957 14399
rect 16908 14368 16957 14396
rect 16908 14356 16914 14368
rect 16945 14365 16957 14368
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 18417 14399 18475 14405
rect 18417 14365 18429 14399
rect 18463 14365 18475 14399
rect 18598 14396 18604 14408
rect 18559 14368 18604 14396
rect 18417 14359 18475 14365
rect 18598 14356 18604 14368
rect 18656 14356 18662 14408
rect 20088 14405 20116 14436
rect 22370 14424 22376 14436
rect 22428 14424 22434 14476
rect 23198 14464 23204 14476
rect 23111 14436 23204 14464
rect 23198 14424 23204 14436
rect 23256 14464 23262 14476
rect 25314 14464 25320 14476
rect 23256 14436 25320 14464
rect 23256 14424 23262 14436
rect 25314 14424 25320 14436
rect 25372 14424 25378 14476
rect 20073 14399 20131 14405
rect 20073 14365 20085 14399
rect 20119 14365 20131 14399
rect 20254 14396 20260 14408
rect 20215 14368 20260 14396
rect 20073 14359 20131 14365
rect 20254 14356 20260 14368
rect 20312 14356 20318 14408
rect 20438 14396 20444 14408
rect 20399 14368 20444 14396
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 22922 14396 22928 14408
rect 22883 14368 22928 14396
rect 22922 14356 22928 14368
rect 22980 14356 22986 14408
rect 26237 14399 26295 14405
rect 26237 14365 26249 14399
rect 26283 14365 26295 14399
rect 26237 14359 26295 14365
rect 3786 14328 3792 14340
rect 2976 14300 3792 14328
rect 3786 14288 3792 14300
rect 3844 14288 3850 14340
rect 20346 14288 20352 14340
rect 20404 14328 20410 14340
rect 20404 14300 20449 14328
rect 20404 14288 20410 14300
rect 1854 14220 1860 14272
rect 1912 14260 1918 14272
rect 2682 14260 2688 14272
rect 1912 14232 2688 14260
rect 1912 14220 1918 14232
rect 2682 14220 2688 14232
rect 2740 14260 2746 14272
rect 2777 14263 2835 14269
rect 2777 14260 2789 14263
rect 2740 14232 2789 14260
rect 2740 14220 2746 14232
rect 2777 14229 2789 14232
rect 2823 14229 2835 14263
rect 2777 14223 2835 14229
rect 3050 14220 3056 14272
rect 3108 14260 3114 14272
rect 3234 14260 3240 14272
rect 3108 14232 3240 14260
rect 3108 14220 3114 14232
rect 3234 14220 3240 14232
rect 3292 14220 3298 14272
rect 13262 14260 13268 14272
rect 13223 14232 13268 14260
rect 13262 14220 13268 14232
rect 13320 14220 13326 14272
rect 13633 14263 13691 14269
rect 13633 14229 13645 14263
rect 13679 14260 13691 14263
rect 14274 14260 14280 14272
rect 13679 14232 14280 14260
rect 13679 14229 13691 14232
rect 13633 14223 13691 14229
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 16022 14260 16028 14272
rect 15983 14232 16028 14260
rect 16022 14220 16028 14232
rect 16080 14220 16086 14272
rect 26252 14260 26280 14359
rect 26326 14356 26332 14408
rect 26384 14396 26390 14408
rect 26620 14396 26648 14504
rect 30374 14492 30380 14544
rect 30432 14532 30438 14544
rect 30926 14532 30932 14544
rect 30432 14504 30932 14532
rect 30432 14492 30438 14504
rect 30926 14492 30932 14504
rect 30984 14492 30990 14544
rect 26702 14399 26760 14405
rect 26702 14396 26714 14399
rect 26384 14368 26429 14396
rect 26620 14368 26714 14396
rect 26384 14356 26390 14368
rect 26702 14365 26714 14368
rect 26748 14365 26760 14399
rect 26702 14359 26760 14365
rect 34514 14356 34520 14408
rect 34572 14396 34578 14408
rect 35161 14399 35219 14405
rect 35161 14396 35173 14399
rect 34572 14368 35173 14396
rect 34572 14356 34578 14368
rect 35161 14365 35173 14368
rect 35207 14365 35219 14399
rect 35161 14359 35219 14365
rect 26510 14328 26516 14340
rect 26471 14300 26516 14328
rect 26510 14288 26516 14300
rect 26568 14288 26574 14340
rect 26605 14331 26663 14337
rect 26605 14297 26617 14331
rect 26651 14328 26663 14331
rect 26786 14328 26792 14340
rect 26651 14300 26792 14328
rect 26651 14297 26663 14300
rect 26605 14291 26663 14297
rect 26786 14288 26792 14300
rect 26844 14288 26850 14340
rect 31846 14288 31852 14340
rect 31904 14328 31910 14340
rect 34606 14328 34612 14340
rect 31904 14300 34612 14328
rect 31904 14288 31910 14300
rect 34606 14288 34612 14300
rect 34664 14328 34670 14340
rect 34885 14331 34943 14337
rect 34885 14328 34897 14331
rect 34664 14300 34897 14328
rect 34664 14288 34670 14300
rect 34885 14297 34897 14300
rect 34931 14297 34943 14331
rect 34885 14291 34943 14297
rect 35069 14331 35127 14337
rect 35069 14297 35081 14331
rect 35115 14297 35127 14331
rect 35176 14328 35204 14359
rect 35250 14356 35256 14408
rect 35308 14405 35314 14408
rect 35308 14396 35316 14405
rect 35308 14368 35353 14396
rect 35308 14359 35316 14368
rect 35308 14356 35314 14359
rect 35802 14356 35808 14408
rect 35860 14396 35866 14408
rect 35897 14399 35955 14405
rect 35897 14396 35909 14399
rect 35860 14368 35909 14396
rect 35860 14356 35866 14368
rect 35897 14365 35909 14368
rect 35943 14365 35955 14399
rect 36170 14396 36176 14408
rect 36131 14368 36176 14396
rect 35897 14359 35955 14365
rect 36170 14356 36176 14368
rect 36228 14356 36234 14408
rect 36081 14331 36139 14337
rect 36081 14328 36093 14331
rect 35176 14300 36093 14328
rect 35069 14291 35127 14297
rect 36081 14297 36093 14300
rect 36127 14297 36139 14331
rect 36081 14291 36139 14297
rect 26694 14260 26700 14272
rect 26252 14232 26700 14260
rect 26694 14220 26700 14232
rect 26752 14220 26758 14272
rect 33594 14220 33600 14272
rect 33652 14260 33658 14272
rect 35084 14260 35112 14291
rect 35894 14260 35900 14272
rect 33652 14232 35900 14260
rect 33652 14220 33658 14232
rect 35894 14220 35900 14232
rect 35952 14220 35958 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 1670 14056 1676 14068
rect 1631 14028 1676 14056
rect 1670 14016 1676 14028
rect 1728 14016 1734 14068
rect 2593 14059 2651 14065
rect 2593 14025 2605 14059
rect 2639 14056 2651 14059
rect 2866 14056 2872 14068
rect 2639 14028 2872 14056
rect 2639 14025 2651 14028
rect 2593 14019 2651 14025
rect 2866 14016 2872 14028
rect 2924 14016 2930 14068
rect 2961 14059 3019 14065
rect 2961 14025 2973 14059
rect 3007 14056 3019 14059
rect 3418 14056 3424 14068
rect 3007 14028 3424 14056
rect 3007 14025 3019 14028
rect 2961 14019 3019 14025
rect 3418 14016 3424 14028
rect 3476 14056 3482 14068
rect 4801 14059 4859 14065
rect 4801 14056 4813 14059
rect 3476 14028 4813 14056
rect 3476 14016 3482 14028
rect 4801 14025 4813 14028
rect 4847 14025 4859 14059
rect 14274 14056 14280 14068
rect 14187 14028 14280 14056
rect 4801 14019 4859 14025
rect 14274 14016 14280 14028
rect 14332 14056 14338 14068
rect 14918 14056 14924 14068
rect 14332 14028 14924 14056
rect 14332 14016 14338 14028
rect 14918 14016 14924 14028
rect 14976 14016 14982 14068
rect 16206 14016 16212 14068
rect 16264 14056 16270 14068
rect 17497 14059 17555 14065
rect 17497 14056 17509 14059
rect 16264 14028 17509 14056
rect 16264 14016 16270 14028
rect 17497 14025 17509 14028
rect 17543 14056 17555 14059
rect 18598 14056 18604 14068
rect 17543 14028 18604 14056
rect 17543 14025 17555 14028
rect 17497 14019 17555 14025
rect 18598 14016 18604 14028
rect 18656 14016 18662 14068
rect 26418 14056 26424 14068
rect 22066 14028 26424 14056
rect 3789 13991 3847 13997
rect 3789 13988 3801 13991
rect 2148 13960 3801 13988
rect 1854 13920 1860 13932
rect 1815 13892 1860 13920
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 2148 13929 2176 13960
rect 3789 13957 3801 13960
rect 3835 13957 3847 13991
rect 13164 13991 13222 13997
rect 3789 13951 3847 13957
rect 3988 13960 4752 13988
rect 3988 13932 4016 13960
rect 2041 13923 2099 13929
rect 2041 13889 2053 13923
rect 2087 13889 2099 13923
rect 2041 13883 2099 13889
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13889 2191 13923
rect 3970 13920 3976 13932
rect 3931 13892 3976 13920
rect 2133 13883 2191 13889
rect 2056 13852 2084 13883
rect 3970 13880 3976 13892
rect 4028 13880 4034 13932
rect 4724 13929 4752 13960
rect 13164 13957 13176 13991
rect 13210 13988 13222 13991
rect 13262 13988 13268 14000
rect 13210 13960 13268 13988
rect 13210 13957 13222 13960
rect 13164 13951 13222 13957
rect 13262 13948 13268 13960
rect 13320 13948 13326 14000
rect 16942 13948 16948 14000
rect 17000 13988 17006 14000
rect 17221 13991 17279 13997
rect 17221 13988 17233 13991
rect 17000 13960 17233 13988
rect 17000 13948 17006 13960
rect 17221 13957 17233 13960
rect 17267 13957 17279 13991
rect 17221 13951 17279 13957
rect 19429 13991 19487 13997
rect 19429 13957 19441 13991
rect 19475 13988 19487 13991
rect 22066 13988 22094 14028
rect 26418 14016 26424 14028
rect 26476 14016 26482 14068
rect 32674 14016 32680 14068
rect 32732 14056 32738 14068
rect 33689 14059 33747 14065
rect 33689 14056 33701 14059
rect 32732 14028 33701 14056
rect 32732 14016 32738 14028
rect 33689 14025 33701 14028
rect 33735 14056 33747 14059
rect 35250 14056 35256 14068
rect 33735 14028 35256 14056
rect 33735 14025 33747 14028
rect 33689 14019 33747 14025
rect 35250 14016 35256 14028
rect 35308 14016 35314 14068
rect 19475 13960 22094 13988
rect 19475 13957 19487 13960
rect 19429 13951 19487 13957
rect 22278 13948 22284 14000
rect 22336 13988 22342 14000
rect 22373 13991 22431 13997
rect 22373 13988 22385 13991
rect 22336 13960 22385 13988
rect 22336 13948 22342 13960
rect 22373 13957 22385 13960
rect 22419 13988 22431 13991
rect 23290 13988 23296 14000
rect 22419 13960 23296 13988
rect 22419 13957 22431 13960
rect 22373 13951 22431 13957
rect 23290 13948 23296 13960
rect 23348 13948 23354 14000
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13889 4215 13923
rect 4157 13883 4215 13889
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 4709 13923 4767 13929
rect 4709 13889 4721 13923
rect 4755 13889 4767 13923
rect 4709 13883 4767 13889
rect 9024 13923 9082 13929
rect 9024 13889 9036 13923
rect 9070 13920 9082 13923
rect 9490 13920 9496 13932
rect 9070 13892 9496 13920
rect 9070 13889 9082 13892
rect 9024 13883 9082 13889
rect 2774 13852 2780 13864
rect 2056 13824 2780 13852
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 3053 13855 3111 13861
rect 3053 13821 3065 13855
rect 3099 13852 3111 13855
rect 3142 13852 3148 13864
rect 3099 13824 3148 13852
rect 3099 13821 3111 13824
rect 3053 13815 3111 13821
rect 3142 13812 3148 13824
rect 3200 13812 3206 13864
rect 3237 13855 3295 13861
rect 3237 13821 3249 13855
rect 3283 13852 3295 13855
rect 3786 13852 3792 13864
rect 3283 13824 3792 13852
rect 3283 13821 3295 13824
rect 3237 13815 3295 13821
rect 3786 13812 3792 13824
rect 3844 13812 3850 13864
rect 4172 13852 4200 13883
rect 4080 13824 4200 13852
rect 3160 13784 3188 13812
rect 4080 13784 4108 13824
rect 3160 13756 4108 13784
rect 3786 13676 3792 13728
rect 3844 13716 3850 13728
rect 4264 13716 4292 13883
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13889 14979 13923
rect 15102 13920 15108 13932
rect 15063 13892 15108 13920
rect 14921 13883 14979 13889
rect 8754 13852 8760 13864
rect 8715 13824 8760 13852
rect 8754 13812 8760 13824
rect 8812 13812 8818 13864
rect 12894 13852 12900 13864
rect 12855 13824 12900 13852
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 14936 13852 14964 13883
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 15197 13923 15255 13929
rect 15197 13889 15209 13923
rect 15243 13920 15255 13923
rect 15470 13920 15476 13932
rect 15243 13892 15476 13920
rect 15243 13889 15255 13892
rect 15197 13883 15255 13889
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 17310 13880 17316 13932
rect 17368 13920 17374 13932
rect 17405 13923 17463 13929
rect 17405 13920 17417 13923
rect 17368 13892 17417 13920
rect 17368 13880 17374 13892
rect 17405 13889 17417 13892
rect 17451 13889 17463 13923
rect 17405 13883 17463 13889
rect 17954 13880 17960 13932
rect 18012 13920 18018 13932
rect 18506 13920 18512 13932
rect 18012 13892 18512 13920
rect 18012 13880 18018 13892
rect 18506 13880 18512 13892
rect 18564 13920 18570 13932
rect 18693 13923 18751 13929
rect 18693 13920 18705 13923
rect 18564 13892 18705 13920
rect 18564 13880 18570 13892
rect 18693 13889 18705 13892
rect 18739 13889 18751 13923
rect 19150 13920 19156 13932
rect 19111 13892 19156 13920
rect 18693 13883 18751 13889
rect 19150 13880 19156 13892
rect 19208 13880 19214 13932
rect 22189 13923 22247 13929
rect 22189 13920 22201 13923
rect 19260 13892 22201 13920
rect 15010 13852 15016 13864
rect 14923 13824 15016 13852
rect 15010 13812 15016 13824
rect 15068 13852 15074 13864
rect 16298 13852 16304 13864
rect 15068 13824 16304 13852
rect 15068 13812 15074 13824
rect 16298 13812 16304 13824
rect 16356 13852 16362 13864
rect 19260 13852 19288 13892
rect 22189 13889 22201 13892
rect 22235 13920 22247 13923
rect 22465 13923 22523 13929
rect 22235 13892 22416 13920
rect 22235 13889 22247 13892
rect 22189 13883 22247 13889
rect 16356 13824 19288 13852
rect 22005 13855 22063 13861
rect 16356 13812 16362 13824
rect 22005 13821 22017 13855
rect 22051 13852 22063 13855
rect 22278 13852 22284 13864
rect 22051 13824 22284 13852
rect 22051 13821 22063 13824
rect 22005 13815 22063 13821
rect 22278 13812 22284 13824
rect 22336 13812 22342 13864
rect 22388 13852 22416 13892
rect 22465 13889 22477 13923
rect 22511 13920 22523 13923
rect 23198 13920 23204 13932
rect 22511 13892 23204 13920
rect 22511 13889 22523 13892
rect 22465 13883 22523 13889
rect 23198 13880 23204 13892
rect 23256 13880 23262 13932
rect 23385 13923 23443 13929
rect 23385 13889 23397 13923
rect 23431 13920 23443 13923
rect 24854 13920 24860 13932
rect 23431 13892 24860 13920
rect 23431 13889 23443 13892
rect 23385 13883 23443 13889
rect 24854 13880 24860 13892
rect 24912 13880 24918 13932
rect 32398 13880 32404 13932
rect 32456 13920 32462 13932
rect 32565 13923 32623 13929
rect 32565 13920 32577 13923
rect 32456 13892 32577 13920
rect 32456 13880 32462 13892
rect 32565 13889 32577 13892
rect 32611 13889 32623 13923
rect 32565 13883 32623 13889
rect 25958 13852 25964 13864
rect 22388 13824 25964 13852
rect 25958 13812 25964 13824
rect 26016 13852 26022 13864
rect 32306 13852 32312 13864
rect 26016 13824 28948 13852
rect 32267 13824 32312 13852
rect 26016 13812 26022 13824
rect 28920 13784 28948 13824
rect 32306 13812 32312 13824
rect 32364 13812 32370 13864
rect 29086 13784 29092 13796
rect 28920 13756 29092 13784
rect 29086 13744 29092 13756
rect 29144 13744 29150 13796
rect 10134 13716 10140 13728
rect 3844 13688 4292 13716
rect 10095 13688 10140 13716
rect 3844 13676 3850 13688
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 14734 13716 14740 13728
rect 14695 13688 14740 13716
rect 14734 13676 14740 13688
rect 14792 13676 14798 13728
rect 24578 13676 24584 13728
rect 24636 13716 24642 13728
rect 24673 13719 24731 13725
rect 24673 13716 24685 13719
rect 24636 13688 24685 13716
rect 24636 13676 24642 13688
rect 24673 13685 24685 13688
rect 24719 13685 24731 13719
rect 24673 13679 24731 13685
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 2869 13515 2927 13521
rect 2869 13512 2881 13515
rect 2832 13484 2881 13512
rect 2832 13472 2838 13484
rect 2869 13481 2881 13484
rect 2915 13481 2927 13515
rect 2869 13475 2927 13481
rect 3970 13472 3976 13524
rect 4028 13512 4034 13524
rect 4157 13515 4215 13521
rect 4157 13512 4169 13515
rect 4028 13484 4169 13512
rect 4028 13472 4034 13484
rect 4157 13481 4169 13484
rect 4203 13481 4215 13515
rect 4157 13475 4215 13481
rect 15746 13472 15752 13524
rect 15804 13512 15810 13524
rect 15804 13484 20576 13512
rect 15804 13472 15810 13484
rect 18785 13447 18843 13453
rect 18785 13413 18797 13447
rect 18831 13444 18843 13447
rect 19978 13444 19984 13456
rect 18831 13416 19984 13444
rect 18831 13413 18843 13416
rect 18785 13407 18843 13413
rect 19978 13404 19984 13416
rect 20036 13444 20042 13456
rect 20438 13444 20444 13456
rect 20036 13416 20444 13444
rect 20036 13404 20042 13416
rect 20438 13404 20444 13416
rect 20496 13404 20502 13456
rect 3050 13376 3056 13388
rect 2746 13348 3056 13376
rect 2746 13320 2774 13348
rect 3050 13336 3056 13348
rect 3108 13336 3114 13388
rect 9766 13376 9772 13388
rect 8234 13362 9772 13376
rect 8220 13348 9772 13362
rect 2746 13268 2780 13320
rect 2832 13308 2838 13320
rect 3142 13308 3148 13320
rect 2832 13280 2879 13308
rect 3103 13280 3148 13308
rect 2832 13268 2838 13280
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 6638 13268 6644 13320
rect 6696 13308 6702 13320
rect 8220 13308 8248 13348
rect 9766 13336 9772 13348
rect 9824 13336 9830 13388
rect 17865 13379 17923 13385
rect 17865 13345 17877 13379
rect 17911 13376 17923 13379
rect 19150 13376 19156 13388
rect 17911 13348 19156 13376
rect 17911 13345 17923 13348
rect 17865 13339 17923 13345
rect 19150 13336 19156 13348
rect 19208 13336 19214 13388
rect 20548 13376 20576 13484
rect 21910 13472 21916 13524
rect 21968 13512 21974 13524
rect 22097 13515 22155 13521
rect 22097 13512 22109 13515
rect 21968 13484 22109 13512
rect 21968 13472 21974 13484
rect 22097 13481 22109 13484
rect 22143 13481 22155 13515
rect 22097 13475 22155 13481
rect 23382 13472 23388 13524
rect 23440 13512 23446 13524
rect 28350 13512 28356 13524
rect 23440 13484 28356 13512
rect 23440 13472 23446 13484
rect 28350 13472 28356 13484
rect 28408 13472 28414 13524
rect 32306 13472 32312 13524
rect 32364 13512 32370 13524
rect 32493 13515 32551 13521
rect 32493 13512 32505 13515
rect 32364 13484 32505 13512
rect 32364 13472 32370 13484
rect 32493 13481 32505 13484
rect 32539 13481 32551 13515
rect 32493 13475 32551 13481
rect 24578 13376 24584 13388
rect 20548 13348 22094 13376
rect 24539 13348 24584 13376
rect 6696 13280 8248 13308
rect 12161 13311 12219 13317
rect 6696 13268 6702 13280
rect 12161 13277 12173 13311
rect 12207 13308 12219 13311
rect 12894 13308 12900 13320
rect 12207 13280 12900 13308
rect 12207 13277 12219 13280
rect 12161 13271 12219 13277
rect 12894 13268 12900 13280
rect 12952 13268 12958 13320
rect 16942 13268 16948 13320
rect 17000 13308 17006 13320
rect 17129 13311 17187 13317
rect 17129 13308 17141 13311
rect 17000 13280 17141 13308
rect 17000 13268 17006 13280
rect 17129 13277 17141 13280
rect 17175 13277 17187 13311
rect 17129 13271 17187 13277
rect 17310 13268 17316 13320
rect 17368 13308 17374 13320
rect 17773 13311 17831 13317
rect 17773 13308 17785 13311
rect 17368 13280 17785 13308
rect 17368 13268 17374 13280
rect 17773 13277 17785 13280
rect 17819 13277 17831 13311
rect 18506 13308 18512 13320
rect 18467 13280 18512 13308
rect 17773 13271 17831 13277
rect 18506 13268 18512 13280
rect 18564 13268 18570 13320
rect 18598 13268 18604 13320
rect 18656 13308 18662 13320
rect 18693 13311 18751 13317
rect 18693 13308 18705 13311
rect 18656 13280 18705 13308
rect 18656 13268 18662 13280
rect 18693 13277 18705 13280
rect 18739 13277 18751 13311
rect 18693 13271 18751 13277
rect 2501 13243 2559 13249
rect 2501 13209 2513 13243
rect 2547 13240 2559 13243
rect 2746 13240 2774 13268
rect 2866 13240 2872 13252
rect 2924 13249 2930 13252
rect 2547 13212 2774 13240
rect 2836 13212 2872 13240
rect 2547 13209 2559 13212
rect 2501 13203 2559 13209
rect 2866 13200 2872 13212
rect 2924 13203 2936 13249
rect 2924 13200 2930 13203
rect 3234 13200 3240 13252
rect 3292 13240 3298 13252
rect 3973 13243 4031 13249
rect 3973 13240 3985 13243
rect 3292 13212 3985 13240
rect 3292 13200 3298 13212
rect 3973 13209 3985 13212
rect 4019 13209 4031 13243
rect 3973 13203 4031 13209
rect 4154 13200 4160 13252
rect 4212 13240 4218 13252
rect 4614 13240 4620 13252
rect 4212 13212 4620 13240
rect 4212 13200 4218 13212
rect 4614 13200 4620 13212
rect 4672 13200 4678 13252
rect 7466 13240 7472 13252
rect 7427 13212 7472 13240
rect 7466 13200 7472 13212
rect 7524 13200 7530 13252
rect 7558 13200 7564 13252
rect 7616 13240 7622 13252
rect 7929 13243 7987 13249
rect 7616 13212 7661 13240
rect 7616 13200 7622 13212
rect 7929 13209 7941 13243
rect 7975 13240 7987 13243
rect 8202 13240 8208 13252
rect 7975 13212 8208 13240
rect 7975 13209 7987 13212
rect 7929 13203 7987 13209
rect 8202 13200 8208 13212
rect 8260 13200 8266 13252
rect 8294 13200 8300 13252
rect 8352 13240 8358 13252
rect 10413 13243 10471 13249
rect 8352 13212 8397 13240
rect 8352 13200 8358 13212
rect 10413 13209 10425 13243
rect 10459 13240 10471 13243
rect 10459 13212 12434 13240
rect 10459 13209 10471 13212
rect 10413 13203 10471 13209
rect 4338 13172 4344 13184
rect 4299 13144 4344 13172
rect 4338 13132 4344 13144
rect 4396 13132 4402 13184
rect 5994 13132 6000 13184
rect 6052 13172 6058 13184
rect 7193 13175 7251 13181
rect 7193 13172 7205 13175
rect 6052 13144 7205 13172
rect 6052 13132 6058 13144
rect 7193 13141 7205 13144
rect 7239 13141 7251 13175
rect 8478 13172 8484 13184
rect 8439 13144 8484 13172
rect 7193 13135 7251 13141
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 12406 13172 12434 13212
rect 12802 13200 12808 13252
rect 12860 13240 12866 13252
rect 14277 13243 14335 13249
rect 14277 13240 14289 13243
rect 12860 13212 14289 13240
rect 12860 13200 12866 13212
rect 14277 13209 14289 13212
rect 14323 13209 14335 13243
rect 18708 13240 18736 13271
rect 19242 13268 19248 13320
rect 19300 13308 19306 13320
rect 19429 13311 19487 13317
rect 19429 13308 19441 13311
rect 19300 13280 19441 13308
rect 19300 13268 19306 13280
rect 19429 13277 19441 13280
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 19613 13311 19671 13317
rect 19613 13277 19625 13311
rect 19659 13277 19671 13311
rect 20806 13308 20812 13320
rect 20767 13280 20812 13308
rect 19613 13271 19671 13277
rect 19628 13240 19656 13271
rect 20806 13268 20812 13280
rect 20864 13268 20870 13320
rect 22066 13308 22094 13348
rect 24578 13336 24584 13348
rect 24636 13336 24642 13388
rect 26421 13311 26479 13317
rect 26421 13308 26433 13311
rect 22066 13280 26433 13308
rect 26421 13277 26433 13280
rect 26467 13277 26479 13311
rect 26421 13271 26479 13277
rect 29086 13268 29092 13320
rect 29144 13308 29150 13320
rect 29917 13311 29975 13317
rect 29917 13308 29929 13311
rect 29144 13280 29929 13308
rect 29144 13268 29150 13280
rect 29917 13277 29929 13280
rect 29963 13277 29975 13311
rect 30190 13308 30196 13320
rect 30151 13280 30196 13308
rect 29917 13271 29975 13277
rect 18708 13212 19656 13240
rect 19797 13243 19855 13249
rect 14277 13203 14335 13209
rect 19797 13209 19809 13243
rect 19843 13240 19855 13243
rect 20438 13240 20444 13252
rect 19843 13212 20444 13240
rect 19843 13209 19855 13212
rect 19797 13203 19855 13209
rect 20438 13200 20444 13212
rect 20496 13200 20502 13252
rect 24848 13243 24906 13249
rect 24848 13209 24860 13243
rect 24894 13240 24906 13243
rect 27154 13240 27160 13252
rect 24894 13212 27160 13240
rect 24894 13209 24906 13212
rect 24848 13203 24906 13209
rect 27154 13200 27160 13212
rect 27212 13200 27218 13252
rect 29932 13240 29960 13271
rect 30190 13268 30196 13280
rect 30248 13268 30254 13320
rect 30466 13240 30472 13252
rect 29932 13212 30472 13240
rect 30466 13200 30472 13212
rect 30524 13200 30530 13252
rect 31205 13243 31263 13249
rect 31205 13209 31217 13243
rect 31251 13240 31263 13243
rect 32122 13240 32128 13252
rect 31251 13212 32128 13240
rect 31251 13209 31263 13212
rect 31205 13203 31263 13209
rect 32122 13200 32128 13212
rect 32180 13200 32186 13252
rect 12986 13172 12992 13184
rect 12406 13144 12992 13172
rect 12986 13132 12992 13144
rect 13044 13172 13050 13184
rect 15565 13175 15623 13181
rect 15565 13172 15577 13175
rect 13044 13144 15577 13172
rect 13044 13132 13050 13144
rect 15565 13141 15577 13144
rect 15611 13141 15623 13175
rect 15565 13135 15623 13141
rect 19058 13132 19064 13184
rect 19116 13172 19122 13184
rect 19426 13172 19432 13184
rect 19116 13144 19432 13172
rect 19116 13132 19122 13144
rect 19426 13132 19432 13144
rect 19484 13132 19490 13184
rect 25961 13175 26019 13181
rect 25961 13141 25973 13175
rect 26007 13172 26019 13175
rect 26326 13172 26332 13184
rect 26007 13144 26332 13172
rect 26007 13141 26019 13144
rect 25961 13135 26019 13141
rect 26326 13132 26332 13144
rect 26384 13132 26390 13184
rect 26602 13172 26608 13184
rect 26563 13144 26608 13172
rect 26602 13132 26608 13144
rect 26660 13132 26666 13184
rect 29730 13172 29736 13184
rect 29691 13144 29736 13172
rect 29730 13132 29736 13144
rect 29788 13132 29794 13184
rect 30101 13175 30159 13181
rect 30101 13141 30113 13175
rect 30147 13172 30159 13175
rect 30558 13172 30564 13184
rect 30147 13144 30564 13172
rect 30147 13141 30159 13144
rect 30101 13135 30159 13141
rect 30558 13132 30564 13144
rect 30616 13132 30622 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 3421 12971 3479 12977
rect 3421 12937 3433 12971
rect 3467 12968 3479 12971
rect 4154 12968 4160 12980
rect 3467 12940 4160 12968
rect 3467 12937 3479 12940
rect 3421 12931 3479 12937
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 5994 12968 6000 12980
rect 5955 12940 6000 12968
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 9769 12971 9827 12977
rect 9769 12937 9781 12971
rect 9815 12968 9827 12971
rect 10134 12968 10140 12980
rect 9815 12940 10140 12968
rect 9815 12937 9827 12940
rect 9769 12931 9827 12937
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 10226 12928 10232 12980
rect 10284 12968 10290 12980
rect 10873 12971 10931 12977
rect 10873 12968 10885 12971
rect 10284 12940 10885 12968
rect 10284 12928 10290 12940
rect 10873 12937 10885 12940
rect 10919 12937 10931 12971
rect 14737 12971 14795 12977
rect 10873 12931 10931 12937
rect 12452 12940 12756 12968
rect 2685 12903 2743 12909
rect 2685 12869 2697 12903
rect 2731 12900 2743 12903
rect 3234 12900 3240 12912
rect 2731 12872 3240 12900
rect 2731 12869 2743 12872
rect 2685 12863 2743 12869
rect 3234 12860 3240 12872
rect 3292 12860 3298 12912
rect 3970 12860 3976 12912
rect 4028 12900 4034 12912
rect 4338 12900 4344 12912
rect 4028 12872 4344 12900
rect 4028 12860 4034 12872
rect 4338 12860 4344 12872
rect 4396 12900 4402 12912
rect 8754 12900 8760 12912
rect 4396 12872 8760 12900
rect 4396 12860 4402 12872
rect 2593 12835 2651 12841
rect 2593 12801 2605 12835
rect 2639 12832 2651 12835
rect 3142 12832 3148 12844
rect 2639 12804 3148 12832
rect 2639 12801 2651 12804
rect 2593 12795 2651 12801
rect 3142 12792 3148 12804
rect 3200 12832 3206 12844
rect 4062 12832 4068 12844
rect 3200 12804 4068 12832
rect 3200 12792 3206 12804
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 4632 12841 4660 12872
rect 8754 12860 8760 12872
rect 8812 12860 8818 12912
rect 10502 12900 10508 12912
rect 8864 12872 10180 12900
rect 10463 12872 10508 12900
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12801 4675 12835
rect 4617 12795 4675 12801
rect 4884 12835 4942 12841
rect 4884 12801 4896 12835
rect 4930 12832 4942 12835
rect 5442 12832 5448 12844
rect 4930 12804 5448 12832
rect 4930 12801 4942 12804
rect 4884 12795 4942 12801
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 7558 12792 7564 12844
rect 7616 12832 7622 12844
rect 8864 12832 8892 12872
rect 10042 12832 10048 12844
rect 7616 12804 8892 12832
rect 10003 12804 10048 12832
rect 7616 12792 7622 12804
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 10152 12841 10180 12872
rect 10502 12860 10508 12872
rect 10560 12860 10566 12912
rect 12452 12909 12480 12940
rect 12437 12903 12495 12909
rect 12437 12869 12449 12903
rect 12483 12869 12495 12903
rect 12437 12863 12495 12869
rect 12621 12903 12679 12909
rect 12621 12869 12633 12903
rect 12667 12869 12679 12903
rect 12728 12900 12756 12940
rect 14737 12937 14749 12971
rect 14783 12968 14795 12971
rect 15102 12968 15108 12980
rect 14783 12940 15108 12968
rect 14783 12937 14795 12940
rect 14737 12931 14795 12937
rect 15102 12928 15108 12940
rect 15160 12968 15166 12980
rect 16942 12968 16948 12980
rect 15160 12940 16948 12968
rect 15160 12928 15166 12940
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 17126 12928 17132 12980
rect 17184 12968 17190 12980
rect 17497 12971 17555 12977
rect 17184 12940 17356 12968
rect 17184 12928 17190 12940
rect 14182 12900 14188 12912
rect 12728 12872 14188 12900
rect 12621 12863 12679 12869
rect 10137 12835 10195 12841
rect 10137 12801 10149 12835
rect 10183 12832 10195 12835
rect 10410 12832 10416 12844
rect 10183 12804 10416 12832
rect 10183 12801 10195 12804
rect 10137 12795 10195 12801
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 10226 12724 10232 12776
rect 10284 12724 10290 12776
rect 12636 12696 12664 12863
rect 14182 12860 14188 12872
rect 14240 12860 14246 12912
rect 15470 12860 15476 12912
rect 15528 12900 15534 12912
rect 17328 12900 17356 12940
rect 17497 12937 17509 12971
rect 17543 12968 17555 12971
rect 21266 12968 21272 12980
rect 17543 12940 21272 12968
rect 17543 12937 17555 12940
rect 17497 12931 17555 12937
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 24670 12968 24676 12980
rect 24631 12940 24676 12968
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 27154 12968 27160 12980
rect 27115 12940 27160 12968
rect 27154 12928 27160 12940
rect 27212 12928 27218 12980
rect 29454 12928 29460 12980
rect 29512 12968 29518 12980
rect 29917 12971 29975 12977
rect 29917 12968 29929 12971
rect 29512 12940 29929 12968
rect 29512 12928 29518 12940
rect 29917 12937 29929 12940
rect 29963 12937 29975 12971
rect 29917 12931 29975 12937
rect 31389 12971 31447 12977
rect 31389 12937 31401 12971
rect 31435 12968 31447 12971
rect 33689 12971 33747 12977
rect 33689 12968 33701 12971
rect 31435 12940 33701 12968
rect 31435 12937 31447 12940
rect 31389 12931 31447 12937
rect 33689 12937 33701 12940
rect 33735 12968 33747 12971
rect 36170 12968 36176 12980
rect 33735 12940 36176 12968
rect 33735 12937 33747 12940
rect 33689 12931 33747 12937
rect 36170 12928 36176 12940
rect 36228 12928 36234 12980
rect 18874 12900 18880 12912
rect 15528 12872 15700 12900
rect 17328 12872 18880 12900
rect 15528 12860 15534 12872
rect 12894 12792 12900 12844
rect 12952 12832 12958 12844
rect 13357 12835 13415 12841
rect 13357 12832 13369 12835
rect 12952 12804 13369 12832
rect 12952 12792 12958 12804
rect 13357 12801 13369 12804
rect 13403 12801 13415 12835
rect 13357 12795 13415 12801
rect 13624 12835 13682 12841
rect 13624 12801 13636 12835
rect 13670 12832 13682 12835
rect 14734 12832 14740 12844
rect 13670 12804 14740 12832
rect 13670 12801 13682 12804
rect 13624 12795 13682 12801
rect 14734 12792 14740 12804
rect 14792 12792 14798 12844
rect 15378 12832 15384 12844
rect 15339 12804 15384 12832
rect 15378 12792 15384 12804
rect 15436 12792 15442 12844
rect 15562 12832 15568 12844
rect 15523 12804 15568 12832
rect 15562 12792 15568 12804
rect 15620 12792 15626 12844
rect 15672 12841 15700 12872
rect 18874 12860 18880 12872
rect 18932 12900 18938 12912
rect 19245 12903 19303 12909
rect 19245 12900 19257 12903
rect 18932 12872 19257 12900
rect 18932 12860 18938 12872
rect 19245 12869 19257 12872
rect 19291 12869 19303 12903
rect 19245 12863 19303 12869
rect 19337 12903 19395 12909
rect 19337 12869 19349 12903
rect 19383 12900 19395 12903
rect 23385 12903 23443 12909
rect 19383 12872 22094 12900
rect 19383 12869 19395 12872
rect 19337 12863 19395 12869
rect 15657 12835 15715 12841
rect 15657 12801 15669 12835
rect 15703 12801 15715 12835
rect 15657 12795 15715 12801
rect 16853 12835 16911 12841
rect 16853 12801 16865 12835
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 16868 12764 16896 12795
rect 16942 12792 16948 12844
rect 17000 12832 17006 12844
rect 17126 12832 17132 12844
rect 17000 12804 17045 12832
rect 17087 12804 17132 12832
rect 17000 12792 17006 12804
rect 17126 12792 17132 12804
rect 17184 12792 17190 12844
rect 17218 12792 17224 12844
rect 17276 12832 17282 12844
rect 17359 12835 17417 12841
rect 17276 12804 17321 12832
rect 17276 12792 17282 12804
rect 17359 12801 17371 12835
rect 17405 12832 17417 12835
rect 18690 12832 18696 12844
rect 17405 12804 18696 12832
rect 17405 12801 17417 12804
rect 17359 12795 17417 12801
rect 18690 12792 18696 12804
rect 18748 12792 18754 12844
rect 18966 12832 18972 12844
rect 18927 12804 18972 12832
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 19150 12841 19156 12844
rect 19117 12835 19156 12841
rect 19117 12801 19129 12835
rect 19117 12795 19156 12801
rect 19150 12792 19156 12795
rect 19208 12792 19214 12844
rect 19426 12792 19432 12844
rect 19484 12841 19490 12844
rect 19484 12832 19492 12841
rect 22066 12832 22094 12872
rect 23385 12869 23397 12903
rect 23431 12900 23443 12903
rect 26234 12900 26240 12912
rect 23431 12872 26240 12900
rect 23431 12869 23443 12872
rect 23385 12863 23443 12869
rect 26234 12860 26240 12872
rect 26292 12860 26298 12912
rect 26326 12860 26332 12912
rect 26384 12900 26390 12912
rect 26786 12900 26792 12912
rect 26384 12872 26792 12900
rect 26384 12860 26390 12872
rect 26786 12860 26792 12872
rect 26844 12900 26850 12912
rect 27525 12903 27583 12909
rect 27525 12900 27537 12903
rect 26844 12872 27537 12900
rect 26844 12860 26850 12872
rect 27525 12869 27537 12872
rect 27571 12869 27583 12903
rect 28626 12900 28632 12912
rect 28587 12872 28632 12900
rect 27525 12863 27583 12869
rect 28626 12860 28632 12872
rect 28684 12860 28690 12912
rect 30190 12860 30196 12912
rect 30248 12900 30254 12912
rect 30248 12872 31524 12900
rect 30248 12860 30254 12872
rect 25774 12832 25780 12844
rect 19484 12804 19529 12832
rect 22066 12804 23612 12832
rect 25735 12804 25780 12832
rect 19484 12795 19492 12804
rect 19484 12792 19490 12795
rect 23584 12776 23612 12804
rect 25774 12792 25780 12804
rect 25832 12792 25838 12844
rect 25961 12835 26019 12841
rect 25961 12832 25973 12835
rect 25884 12804 25973 12832
rect 16868 12736 19196 12764
rect 19168 12696 19196 12736
rect 19306 12736 23520 12764
rect 19306 12696 19334 12736
rect 12636 12668 13400 12696
rect 3418 12628 3424 12640
rect 3379 12600 3424 12628
rect 3418 12588 3424 12600
rect 3476 12588 3482 12640
rect 3605 12631 3663 12637
rect 3605 12597 3617 12631
rect 3651 12628 3663 12631
rect 4614 12628 4620 12640
rect 3651 12600 4620 12628
rect 3651 12597 3663 12600
rect 3605 12591 3663 12597
rect 4614 12588 4620 12600
rect 4672 12588 4678 12640
rect 11054 12628 11060 12640
rect 11015 12600 11060 12628
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 12618 12628 12624 12640
rect 12579 12600 12624 12628
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 12802 12628 12808 12640
rect 12763 12600 12808 12628
rect 12802 12588 12808 12600
rect 12860 12588 12866 12640
rect 13372 12628 13400 12668
rect 15028 12668 15516 12696
rect 19168 12668 19334 12696
rect 19613 12699 19671 12705
rect 15028 12628 15056 12668
rect 15194 12628 15200 12640
rect 13372 12600 15056 12628
rect 15155 12600 15200 12628
rect 15194 12588 15200 12600
rect 15252 12588 15258 12640
rect 15488 12628 15516 12668
rect 19613 12665 19625 12699
rect 19659 12696 19671 12699
rect 23382 12696 23388 12708
rect 19659 12668 23388 12696
rect 19659 12665 19671 12668
rect 19613 12659 19671 12665
rect 23382 12656 23388 12668
rect 23440 12656 23446 12708
rect 23492 12696 23520 12736
rect 23566 12724 23572 12776
rect 23624 12764 23630 12776
rect 25884 12764 25912 12804
rect 25961 12801 25973 12804
rect 26007 12801 26019 12835
rect 25961 12795 26019 12801
rect 26053 12835 26111 12841
rect 26053 12801 26065 12835
rect 26099 12832 26111 12835
rect 26099 12804 26188 12832
rect 26099 12801 26111 12804
rect 26053 12795 26111 12801
rect 26160 12776 26188 12804
rect 26602 12792 26608 12844
rect 26660 12832 26666 12844
rect 27338 12832 27344 12844
rect 26660 12804 27344 12832
rect 26660 12792 26666 12804
rect 27338 12792 27344 12804
rect 27396 12792 27402 12844
rect 27617 12835 27675 12841
rect 27617 12801 27629 12835
rect 27663 12801 27675 12835
rect 27617 12795 27675 12801
rect 23624 12736 25912 12764
rect 23624 12724 23630 12736
rect 26142 12724 26148 12776
rect 26200 12764 26206 12776
rect 27632 12764 27660 12795
rect 31110 12792 31116 12844
rect 31168 12832 31174 12844
rect 31496 12841 31524 12872
rect 31205 12835 31263 12841
rect 31205 12832 31217 12835
rect 31168 12804 31217 12832
rect 31168 12792 31174 12804
rect 31205 12801 31217 12804
rect 31251 12801 31263 12835
rect 31205 12795 31263 12801
rect 31481 12835 31539 12841
rect 31481 12801 31493 12835
rect 31527 12801 31539 12835
rect 32306 12832 32312 12844
rect 32267 12804 32312 12832
rect 31481 12795 31539 12801
rect 32306 12792 32312 12804
rect 32364 12792 32370 12844
rect 26200 12736 27660 12764
rect 31021 12767 31079 12773
rect 26200 12724 26206 12736
rect 31021 12733 31033 12767
rect 31067 12764 31079 12767
rect 32585 12767 32643 12773
rect 32585 12764 32597 12767
rect 31067 12736 32597 12764
rect 31067 12733 31079 12736
rect 31021 12727 31079 12733
rect 32585 12733 32597 12736
rect 32631 12733 32643 12767
rect 32585 12727 32643 12733
rect 28074 12696 28080 12708
rect 23492 12668 28080 12696
rect 28074 12656 28080 12668
rect 28132 12656 28138 12708
rect 16022 12628 16028 12640
rect 15488 12600 16028 12628
rect 16022 12588 16028 12600
rect 16080 12628 16086 12640
rect 17126 12628 17132 12640
rect 16080 12600 17132 12628
rect 16080 12588 16086 12600
rect 17126 12588 17132 12600
rect 17184 12588 17190 12640
rect 18874 12588 18880 12640
rect 18932 12628 18938 12640
rect 19242 12628 19248 12640
rect 18932 12600 19248 12628
rect 18932 12588 18938 12600
rect 19242 12588 19248 12600
rect 19300 12588 19306 12640
rect 23474 12588 23480 12640
rect 23532 12628 23538 12640
rect 25593 12631 25651 12637
rect 25593 12628 25605 12631
rect 23532 12600 25605 12628
rect 23532 12588 23538 12600
rect 25593 12597 25605 12600
rect 25639 12597 25651 12631
rect 25593 12591 25651 12597
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 6825 12427 6883 12433
rect 6825 12393 6837 12427
rect 6871 12424 6883 12427
rect 7466 12424 7472 12436
rect 6871 12396 7472 12424
rect 6871 12393 6883 12396
rect 6825 12387 6883 12393
rect 7466 12384 7472 12396
rect 7524 12384 7530 12436
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10505 12427 10563 12433
rect 10505 12424 10517 12427
rect 10100 12396 10517 12424
rect 10100 12384 10106 12396
rect 10505 12393 10517 12396
rect 10551 12393 10563 12427
rect 15470 12424 15476 12436
rect 10505 12387 10563 12393
rect 13740 12396 15476 12424
rect 5442 12316 5448 12368
rect 5500 12316 5506 12368
rect 4614 12248 4620 12300
rect 4672 12288 4678 12300
rect 5460 12288 5488 12316
rect 4672 12260 5304 12288
rect 5460 12260 5580 12288
rect 4672 12248 4678 12260
rect 5276 12232 5304 12260
rect 4062 12220 4068 12232
rect 4023 12192 4068 12220
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 4706 12220 4712 12232
rect 4203 12192 4712 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 5258 12180 5264 12232
rect 5316 12220 5322 12232
rect 5445 12223 5503 12229
rect 5445 12220 5457 12223
rect 5316 12192 5457 12220
rect 5316 12180 5322 12192
rect 5445 12189 5457 12192
rect 5491 12189 5503 12223
rect 5552 12220 5580 12260
rect 5701 12223 5759 12229
rect 5701 12220 5713 12223
rect 5552 12192 5713 12220
rect 5445 12183 5503 12189
rect 5701 12189 5713 12192
rect 5747 12189 5759 12223
rect 9122 12220 9128 12232
rect 9083 12192 9128 12220
rect 5701 12183 5759 12189
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 13740 12229 13768 12396
rect 15470 12384 15476 12396
rect 15528 12384 15534 12436
rect 15562 12384 15568 12436
rect 15620 12424 15626 12436
rect 15657 12427 15715 12433
rect 15657 12424 15669 12427
rect 15620 12396 15669 12424
rect 15620 12384 15626 12396
rect 15657 12393 15669 12396
rect 15703 12424 15715 12427
rect 19150 12424 19156 12436
rect 15703 12396 19156 12424
rect 15703 12393 15715 12396
rect 15657 12387 15715 12393
rect 19150 12384 19156 12396
rect 19208 12384 19214 12436
rect 20073 12427 20131 12433
rect 20073 12393 20085 12427
rect 20119 12424 20131 12427
rect 23290 12424 23296 12436
rect 20119 12396 23152 12424
rect 23251 12396 23296 12424
rect 20119 12393 20131 12396
rect 20073 12387 20131 12393
rect 21358 12356 21364 12368
rect 18156 12328 21364 12356
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12189 13507 12223
rect 13449 12183 13507 12189
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12189 13783 12223
rect 14274 12220 14280 12232
rect 14235 12192 14280 12220
rect 13725 12183 13783 12189
rect 9392 12155 9450 12161
rect 9392 12121 9404 12155
rect 9438 12152 9450 12155
rect 9490 12152 9496 12164
rect 9438 12124 9496 12152
rect 9438 12121 9450 12124
rect 9392 12115 9450 12121
rect 9490 12112 9496 12124
rect 9548 12112 9554 12164
rect 13464 12152 13492 12183
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 14826 12220 14832 12232
rect 14476 12192 14832 12220
rect 14476 12152 14504 12192
rect 14826 12180 14832 12192
rect 14884 12220 14890 12232
rect 15286 12220 15292 12232
rect 14884 12192 15292 12220
rect 14884 12180 14890 12192
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 18156 12229 18184 12328
rect 21358 12316 21364 12328
rect 21416 12316 21422 12368
rect 23124 12356 23152 12396
rect 23290 12384 23296 12396
rect 23348 12384 23354 12436
rect 23842 12384 23848 12436
rect 23900 12424 23906 12436
rect 25314 12424 25320 12436
rect 23900 12396 25320 12424
rect 23900 12384 23906 12396
rect 25314 12384 25320 12396
rect 25372 12424 25378 12436
rect 26050 12424 26056 12436
rect 25372 12396 26056 12424
rect 25372 12384 25378 12396
rect 26050 12384 26056 12396
rect 26108 12384 26114 12436
rect 26786 12424 26792 12436
rect 26747 12396 26792 12424
rect 26786 12384 26792 12396
rect 26844 12384 26850 12436
rect 27157 12427 27215 12433
rect 27157 12393 27169 12427
rect 27203 12424 27215 12427
rect 27246 12424 27252 12436
rect 27203 12396 27252 12424
rect 27203 12393 27215 12396
rect 27157 12387 27215 12393
rect 27246 12384 27252 12396
rect 27304 12384 27310 12436
rect 28074 12424 28080 12436
rect 28035 12396 28080 12424
rect 28074 12384 28080 12396
rect 28132 12384 28138 12436
rect 23124 12328 26924 12356
rect 19058 12288 19064 12300
rect 18340 12260 19064 12288
rect 18340 12229 18368 12260
rect 19058 12248 19064 12260
rect 19116 12248 19122 12300
rect 20530 12248 20536 12300
rect 20588 12288 20594 12300
rect 20588 12260 21588 12288
rect 20588 12248 20594 12260
rect 18141 12223 18199 12229
rect 18141 12189 18153 12223
rect 18187 12189 18199 12223
rect 18141 12183 18199 12189
rect 18325 12223 18383 12229
rect 18325 12189 18337 12223
rect 18371 12189 18383 12223
rect 18506 12220 18512 12232
rect 18467 12192 18512 12220
rect 18325 12183 18383 12189
rect 18506 12180 18512 12192
rect 18564 12180 18570 12232
rect 19429 12223 19487 12229
rect 19429 12220 19441 12223
rect 18708 12192 19441 12220
rect 13464 12124 14504 12152
rect 14544 12155 14602 12161
rect 14544 12121 14556 12155
rect 14590 12152 14602 12155
rect 15194 12152 15200 12164
rect 14590 12124 15200 12152
rect 14590 12121 14602 12124
rect 14544 12115 14602 12121
rect 15194 12112 15200 12124
rect 15252 12112 15258 12164
rect 15562 12112 15568 12164
rect 15620 12152 15626 12164
rect 18417 12155 18475 12161
rect 18417 12152 18429 12155
rect 15620 12124 18429 12152
rect 15620 12112 15626 12124
rect 18417 12121 18429 12124
rect 18463 12121 18475 12155
rect 18417 12115 18475 12121
rect 4341 12087 4399 12093
rect 4341 12053 4353 12087
rect 4387 12084 4399 12087
rect 4614 12084 4620 12096
rect 4387 12056 4620 12084
rect 4387 12053 4399 12056
rect 4341 12047 4399 12053
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 13262 12084 13268 12096
rect 13223 12056 13268 12084
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 13630 12084 13636 12096
rect 13591 12056 13636 12084
rect 13630 12044 13636 12056
rect 13688 12044 13694 12096
rect 18708 12093 18736 12192
rect 19429 12189 19441 12192
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 19518 12180 19524 12232
rect 19576 12220 19582 12232
rect 19978 12229 19984 12232
rect 19935 12223 19984 12229
rect 19576 12192 19621 12220
rect 19576 12180 19582 12192
rect 19935 12189 19947 12223
rect 19981 12189 19984 12223
rect 19935 12183 19984 12189
rect 19978 12180 19984 12183
rect 20036 12220 20042 12232
rect 20898 12220 20904 12232
rect 20036 12192 20904 12220
rect 20036 12180 20042 12192
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 21174 12180 21180 12232
rect 21232 12220 21238 12232
rect 21450 12220 21456 12232
rect 21232 12192 21277 12220
rect 21411 12192 21456 12220
rect 21232 12180 21238 12192
rect 21450 12180 21456 12192
rect 21508 12180 21514 12232
rect 19242 12112 19248 12164
rect 19300 12152 19306 12164
rect 19705 12155 19763 12161
rect 19705 12152 19717 12155
rect 19300 12124 19717 12152
rect 19300 12112 19306 12124
rect 19705 12121 19717 12124
rect 19751 12121 19763 12155
rect 19705 12115 19763 12121
rect 19797 12155 19855 12161
rect 19797 12121 19809 12155
rect 19843 12152 19855 12155
rect 20162 12152 20168 12164
rect 19843 12124 20168 12152
rect 19843 12121 19855 12124
rect 19797 12115 19855 12121
rect 20162 12112 20168 12124
rect 20220 12112 20226 12164
rect 21560 12152 21588 12260
rect 24578 12248 24584 12300
rect 24636 12248 24642 12300
rect 26896 12297 26924 12328
rect 26881 12291 26939 12297
rect 26881 12257 26893 12291
rect 26927 12257 26939 12291
rect 28442 12288 28448 12300
rect 26881 12251 26939 12257
rect 28276 12260 28448 12288
rect 21913 12223 21971 12229
rect 21913 12189 21925 12223
rect 21959 12220 21971 12223
rect 24596 12220 24624 12248
rect 28276 12229 28304 12260
rect 28442 12248 28448 12260
rect 28500 12248 28506 12300
rect 30374 12288 30380 12300
rect 28644 12260 30380 12288
rect 21959 12192 24624 12220
rect 26789 12223 26847 12229
rect 21959 12189 21971 12192
rect 21913 12183 21971 12189
rect 26789 12189 26801 12223
rect 26835 12189 26847 12223
rect 26789 12183 26847 12189
rect 28261 12223 28319 12229
rect 28261 12189 28273 12223
rect 28307 12189 28319 12223
rect 28261 12183 28319 12189
rect 28353 12223 28411 12229
rect 28353 12189 28365 12223
rect 28399 12220 28411 12223
rect 28644 12220 28672 12260
rect 30374 12248 30380 12260
rect 30432 12248 30438 12300
rect 28399 12192 28672 12220
rect 28721 12223 28779 12229
rect 28399 12189 28411 12192
rect 28353 12183 28411 12189
rect 28721 12189 28733 12223
rect 28767 12220 28779 12223
rect 30282 12220 30288 12232
rect 28767 12192 30288 12220
rect 28767 12189 28779 12192
rect 28721 12183 28779 12189
rect 22180 12155 22238 12161
rect 21560 12124 22094 12152
rect 18693 12087 18751 12093
rect 18693 12053 18705 12087
rect 18739 12053 18751 12087
rect 20990 12084 20996 12096
rect 20951 12056 20996 12084
rect 18693 12047 18751 12053
rect 20990 12044 20996 12056
rect 21048 12044 21054 12096
rect 21358 12084 21364 12096
rect 21319 12056 21364 12084
rect 21358 12044 21364 12056
rect 21416 12044 21422 12096
rect 22066 12084 22094 12124
rect 22180 12121 22192 12155
rect 22226 12152 22238 12155
rect 22278 12152 22284 12164
rect 22226 12124 22284 12152
rect 22226 12121 22238 12124
rect 22180 12115 22238 12121
rect 22278 12112 22284 12124
rect 22336 12112 22342 12164
rect 24302 12112 24308 12164
rect 24360 12152 24366 12164
rect 24581 12155 24639 12161
rect 24581 12152 24593 12155
rect 24360 12124 24593 12152
rect 24360 12112 24366 12124
rect 24581 12121 24593 12124
rect 24627 12121 24639 12155
rect 26804 12152 26832 12183
rect 30282 12180 30288 12192
rect 30340 12180 30346 12232
rect 24581 12115 24639 12121
rect 24688 12124 26832 12152
rect 28445 12155 28503 12161
rect 24688 12084 24716 12124
rect 28445 12121 28457 12155
rect 28491 12121 28503 12155
rect 28445 12115 28503 12121
rect 22066 12056 24716 12084
rect 24854 12044 24860 12096
rect 24912 12084 24918 12096
rect 25869 12087 25927 12093
rect 25869 12084 25881 12087
rect 24912 12056 25881 12084
rect 24912 12044 24918 12056
rect 25869 12053 25881 12056
rect 25915 12053 25927 12087
rect 28460 12084 28488 12115
rect 28534 12112 28540 12164
rect 28592 12161 28598 12164
rect 28592 12155 28621 12161
rect 28609 12121 28621 12155
rect 30834 12152 30840 12164
rect 30795 12124 30840 12152
rect 28592 12115 28621 12121
rect 28592 12112 28598 12115
rect 30834 12112 30840 12124
rect 30892 12112 30898 12164
rect 30558 12084 30564 12096
rect 28460 12056 30564 12084
rect 25869 12047 25927 12053
rect 30558 12044 30564 12056
rect 30616 12044 30622 12096
rect 32122 12084 32128 12096
rect 32083 12056 32128 12084
rect 32122 12044 32128 12056
rect 32180 12044 32186 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 23477 11883 23535 11889
rect 23477 11849 23489 11883
rect 23523 11880 23535 11883
rect 23566 11880 23572 11892
rect 23523 11852 23572 11880
rect 23523 11849 23535 11852
rect 23477 11843 23535 11849
rect 23566 11840 23572 11852
rect 23624 11840 23630 11892
rect 24118 11880 24124 11892
rect 24079 11852 24124 11880
rect 24118 11840 24124 11852
rect 24176 11840 24182 11892
rect 24302 11880 24308 11892
rect 24263 11852 24308 11880
rect 24302 11840 24308 11852
rect 24360 11840 24366 11892
rect 26513 11883 26571 11889
rect 26513 11849 26525 11883
rect 26559 11880 26571 11883
rect 26786 11880 26792 11892
rect 26559 11852 26792 11880
rect 26559 11849 26571 11852
rect 26513 11843 26571 11849
rect 26786 11840 26792 11852
rect 26844 11840 26850 11892
rect 28442 11880 28448 11892
rect 28403 11852 28448 11880
rect 28442 11840 28448 11852
rect 28500 11840 28506 11892
rect 28629 11883 28687 11889
rect 28629 11849 28641 11883
rect 28675 11880 28687 11883
rect 30834 11880 30840 11892
rect 28675 11852 30840 11880
rect 28675 11849 28687 11852
rect 28629 11843 28687 11849
rect 30834 11840 30840 11852
rect 30892 11840 30898 11892
rect 32309 11883 32367 11889
rect 32309 11849 32321 11883
rect 32355 11880 32367 11883
rect 32398 11880 32404 11892
rect 32355 11852 32404 11880
rect 32355 11849 32367 11852
rect 32309 11843 32367 11849
rect 32398 11840 32404 11852
rect 32456 11840 32462 11892
rect 32674 11880 32680 11892
rect 32635 11852 32680 11880
rect 32674 11840 32680 11852
rect 32732 11840 32738 11892
rect 23842 11812 23848 11824
rect 22066 11784 23848 11812
rect 12989 11747 13047 11753
rect 12989 11713 13001 11747
rect 13035 11744 13047 11747
rect 16482 11744 16488 11756
rect 13035 11716 16488 11744
rect 13035 11713 13047 11716
rect 12989 11707 13047 11713
rect 16482 11704 16488 11716
rect 16540 11704 16546 11756
rect 21450 11704 21456 11756
rect 21508 11744 21514 11756
rect 22066 11744 22094 11784
rect 23842 11772 23848 11784
rect 23900 11772 23906 11824
rect 23937 11815 23995 11821
rect 23937 11781 23949 11815
rect 23983 11812 23995 11815
rect 28258 11812 28264 11824
rect 23983 11784 28264 11812
rect 23983 11781 23995 11784
rect 23937 11775 23995 11781
rect 21508 11716 22094 11744
rect 22364 11747 22422 11753
rect 21508 11704 21514 11716
rect 22364 11713 22376 11747
rect 22410 11744 22422 11747
rect 22410 11716 23152 11744
rect 22410 11713 22422 11716
rect 22364 11707 22422 11713
rect 14182 11636 14188 11688
rect 14240 11676 14246 11688
rect 14737 11679 14795 11685
rect 14737 11676 14749 11679
rect 14240 11648 14749 11676
rect 14240 11636 14246 11648
rect 14737 11645 14749 11648
rect 14783 11676 14795 11679
rect 15102 11676 15108 11688
rect 14783 11648 15108 11676
rect 14783 11645 14795 11648
rect 14737 11639 14795 11645
rect 15102 11636 15108 11648
rect 15160 11636 15166 11688
rect 22002 11636 22008 11688
rect 22060 11676 22066 11688
rect 22097 11679 22155 11685
rect 22097 11676 22109 11679
rect 22060 11648 22109 11676
rect 22060 11636 22066 11648
rect 22097 11645 22109 11648
rect 22143 11645 22155 11679
rect 23124 11676 23152 11716
rect 23474 11676 23480 11688
rect 23124 11648 23480 11676
rect 22097 11639 22155 11645
rect 23474 11636 23480 11648
rect 23532 11636 23538 11688
rect 16482 11568 16488 11620
rect 16540 11608 16546 11620
rect 18230 11608 18236 11620
rect 16540 11580 18236 11608
rect 16540 11568 16546 11580
rect 18230 11568 18236 11580
rect 18288 11568 18294 11620
rect 23382 11568 23388 11620
rect 23440 11608 23446 11620
rect 23952 11608 23980 11775
rect 28258 11772 28264 11784
rect 28316 11772 28322 11824
rect 30190 11772 30196 11824
rect 30248 11812 30254 11824
rect 31665 11815 31723 11821
rect 30248 11784 31616 11812
rect 30248 11772 30254 11784
rect 25866 11744 25872 11756
rect 25827 11716 25872 11744
rect 25866 11704 25872 11716
rect 25924 11704 25930 11756
rect 25962 11747 26020 11753
rect 25962 11713 25974 11747
rect 26008 11713 26020 11747
rect 25962 11707 26020 11713
rect 25222 11636 25228 11688
rect 25280 11676 25286 11688
rect 25976 11676 26004 11707
rect 26050 11704 26056 11756
rect 26108 11744 26114 11756
rect 26418 11753 26424 11756
rect 26145 11747 26203 11753
rect 26145 11744 26157 11747
rect 26108 11716 26157 11744
rect 26108 11704 26114 11716
rect 26145 11713 26157 11716
rect 26191 11713 26203 11747
rect 26145 11707 26203 11713
rect 26237 11747 26295 11753
rect 26237 11713 26249 11747
rect 26283 11713 26295 11747
rect 26237 11707 26295 11713
rect 26375 11747 26424 11753
rect 26375 11713 26387 11747
rect 26421 11713 26424 11747
rect 26375 11707 26424 11713
rect 25280 11648 26004 11676
rect 25280 11636 25286 11648
rect 23440 11580 23980 11608
rect 26252 11608 26280 11707
rect 26418 11704 26424 11707
rect 26476 11744 26482 11756
rect 28534 11744 28540 11756
rect 26476 11716 28540 11744
rect 26476 11704 26482 11716
rect 28534 11704 28540 11716
rect 28592 11704 28598 11756
rect 29457 11747 29515 11753
rect 29457 11713 29469 11747
rect 29503 11744 29515 11747
rect 29730 11744 29736 11756
rect 29503 11716 29736 11744
rect 29503 11713 29515 11716
rect 29457 11707 29515 11713
rect 29730 11704 29736 11716
rect 29788 11704 29794 11756
rect 31386 11704 31392 11756
rect 31444 11744 31450 11756
rect 31481 11747 31539 11753
rect 31481 11744 31493 11747
rect 31444 11716 31493 11744
rect 31444 11704 31450 11716
rect 31481 11713 31493 11716
rect 31527 11713 31539 11747
rect 31588 11744 31616 11784
rect 31665 11781 31677 11815
rect 31711 11812 31723 11815
rect 31846 11812 31852 11824
rect 31711 11784 31852 11812
rect 31711 11781 31723 11784
rect 31665 11775 31723 11781
rect 31846 11772 31852 11784
rect 31904 11812 31910 11824
rect 32582 11812 32588 11824
rect 31904 11784 32588 11812
rect 31904 11772 31910 11784
rect 32582 11772 32588 11784
rect 32640 11772 32646 11824
rect 31757 11747 31815 11753
rect 31757 11744 31769 11747
rect 31588 11716 31769 11744
rect 31481 11707 31539 11713
rect 31757 11713 31769 11716
rect 31803 11713 31815 11747
rect 32490 11744 32496 11756
rect 32451 11716 32496 11744
rect 31757 11707 31815 11713
rect 29178 11676 29184 11688
rect 29139 11648 29184 11676
rect 29178 11636 29184 11648
rect 29236 11636 29242 11688
rect 30558 11676 30564 11688
rect 30519 11648 30564 11676
rect 30558 11636 30564 11648
rect 30616 11636 30622 11688
rect 31772 11676 31800 11707
rect 32490 11704 32496 11716
rect 32548 11704 32554 11756
rect 32769 11747 32827 11753
rect 32769 11713 32781 11747
rect 32815 11713 32827 11747
rect 32769 11707 32827 11713
rect 32784 11676 32812 11707
rect 31772 11648 32812 11676
rect 29086 11608 29092 11620
rect 26252 11580 29092 11608
rect 23440 11568 23446 11580
rect 29086 11568 29092 11580
rect 29144 11568 29150 11620
rect 23566 11500 23572 11552
rect 23624 11540 23630 11552
rect 24121 11543 24179 11549
rect 24121 11540 24133 11543
rect 23624 11512 24133 11540
rect 23624 11500 23630 11512
rect 24121 11509 24133 11512
rect 24167 11540 24179 11543
rect 25406 11540 25412 11552
rect 24167 11512 25412 11540
rect 24167 11509 24179 11512
rect 24121 11503 24179 11509
rect 25406 11500 25412 11512
rect 25464 11540 25470 11552
rect 27982 11540 27988 11552
rect 25464 11512 27988 11540
rect 25464 11500 25470 11512
rect 27982 11500 27988 11512
rect 28040 11540 28046 11552
rect 28445 11543 28503 11549
rect 28445 11540 28457 11543
rect 28040 11512 28457 11540
rect 28040 11500 28046 11512
rect 28445 11509 28457 11512
rect 28491 11509 28503 11543
rect 28445 11503 28503 11509
rect 31297 11543 31355 11549
rect 31297 11509 31309 11543
rect 31343 11540 31355 11543
rect 31478 11540 31484 11552
rect 31343 11512 31484 11540
rect 31343 11509 31355 11512
rect 31297 11503 31355 11509
rect 31478 11500 31484 11512
rect 31536 11500 31542 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 13630 11296 13636 11348
rect 13688 11336 13694 11348
rect 15657 11339 15715 11345
rect 15657 11336 15669 11339
rect 13688 11308 15669 11336
rect 13688 11296 13694 11308
rect 15657 11305 15669 11308
rect 15703 11336 15715 11339
rect 19426 11336 19432 11348
rect 15703 11308 19432 11336
rect 15703 11305 15715 11308
rect 15657 11299 15715 11305
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 21358 11296 21364 11348
rect 21416 11336 21422 11348
rect 23385 11339 23443 11345
rect 23385 11336 23397 11339
rect 21416 11308 23397 11336
rect 21416 11296 21422 11308
rect 23385 11305 23397 11308
rect 23431 11305 23443 11339
rect 32582 11336 32588 11348
rect 32543 11308 32588 11336
rect 23385 11299 23443 11305
rect 32582 11296 32588 11308
rect 32640 11296 32646 11348
rect 16390 11228 16396 11280
rect 16448 11268 16454 11280
rect 17218 11268 17224 11280
rect 16448 11240 17224 11268
rect 16448 11228 16454 11240
rect 17218 11228 17224 11240
rect 17276 11228 17282 11280
rect 6638 11200 6644 11212
rect 6486 11172 6644 11200
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 8754 11160 8760 11212
rect 8812 11200 8818 11212
rect 9125 11203 9183 11209
rect 9125 11200 9137 11203
rect 8812 11172 9137 11200
rect 8812 11160 8818 11172
rect 9125 11169 9137 11172
rect 9171 11169 9183 11203
rect 9125 11163 9183 11169
rect 13262 11160 13268 11212
rect 13320 11200 13326 11212
rect 13320 11172 14412 11200
rect 13320 11160 13326 11172
rect 6178 11132 6184 11144
rect 6139 11104 6184 11132
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 7558 11132 7564 11144
rect 6380 11104 7564 11132
rect 5718 11064 5724 11076
rect 5679 11036 5724 11064
rect 5718 11024 5724 11036
rect 5776 11024 5782 11076
rect 5813 11067 5871 11073
rect 5813 11033 5825 11067
rect 5859 11064 5871 11067
rect 6380 11064 6408 11104
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 9398 11141 9404 11144
rect 9392 11132 9404 11141
rect 9359 11104 9404 11132
rect 9392 11095 9404 11104
rect 9398 11092 9404 11095
rect 9456 11092 9462 11144
rect 14274 11132 14280 11144
rect 14235 11104 14280 11132
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 14384 11132 14412 11172
rect 20990 11160 20996 11212
rect 21048 11200 21054 11212
rect 31478 11200 31484 11212
rect 21048 11172 22140 11200
rect 31439 11172 31484 11200
rect 21048 11160 21054 11172
rect 14533 11135 14591 11141
rect 14533 11132 14545 11135
rect 14384 11104 14545 11132
rect 14533 11101 14545 11104
rect 14579 11101 14591 11135
rect 22002 11132 22008 11144
rect 21963 11104 22008 11132
rect 14533 11095 14591 11101
rect 22002 11092 22008 11104
rect 22060 11092 22066 11144
rect 22112 11132 22140 11172
rect 31478 11160 31484 11172
rect 31536 11160 31542 11212
rect 22261 11135 22319 11141
rect 22261 11132 22273 11135
rect 22112 11104 22273 11132
rect 22261 11101 22273 11104
rect 22307 11101 22319 11135
rect 22261 11095 22319 11101
rect 29914 11092 29920 11144
rect 29972 11132 29978 11144
rect 31205 11135 31263 11141
rect 31205 11132 31217 11135
rect 29972 11104 31217 11132
rect 29972 11092 29978 11104
rect 31205 11101 31217 11104
rect 31251 11101 31263 11135
rect 31205 11095 31263 11101
rect 6546 11064 6552 11076
rect 5859 11036 6408 11064
rect 6507 11036 6552 11064
rect 5859 11033 5871 11036
rect 5813 11027 5871 11033
rect 6546 11024 6552 11036
rect 6604 11024 6610 11076
rect 5442 10996 5448 11008
rect 5403 10968 5448 10996
rect 5442 10956 5448 10968
rect 5500 10956 5506 11008
rect 6454 10956 6460 11008
rect 6512 10996 6518 11008
rect 6733 10999 6791 11005
rect 6733 10996 6745 10999
rect 6512 10968 6745 10996
rect 6512 10956 6518 10968
rect 6733 10965 6745 10968
rect 6779 10965 6791 10999
rect 10502 10996 10508 11008
rect 10463 10968 10508 10996
rect 6733 10959 6791 10965
rect 10502 10956 10508 10968
rect 10560 10956 10566 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 5261 10795 5319 10801
rect 5261 10761 5273 10795
rect 5307 10792 5319 10795
rect 5718 10792 5724 10804
rect 5307 10764 5724 10792
rect 5307 10761 5319 10764
rect 5261 10755 5319 10761
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 9769 10795 9827 10801
rect 9769 10761 9781 10795
rect 9815 10792 9827 10795
rect 10502 10792 10508 10804
rect 9815 10764 10508 10792
rect 9815 10761 9827 10764
rect 9769 10755 9827 10761
rect 10502 10752 10508 10764
rect 10560 10752 10566 10804
rect 14274 10792 14280 10804
rect 14235 10764 14280 10792
rect 14274 10752 14280 10764
rect 14332 10752 14338 10804
rect 29178 10752 29184 10804
rect 29236 10792 29242 10804
rect 29914 10792 29920 10804
rect 29236 10764 29920 10792
rect 29236 10752 29242 10764
rect 29914 10752 29920 10764
rect 29972 10752 29978 10804
rect 3896 10696 5304 10724
rect 3896 10665 3924 10696
rect 5276 10668 5304 10696
rect 9214 10684 9220 10736
rect 9272 10724 9278 10736
rect 10873 10727 10931 10733
rect 10873 10724 10885 10727
rect 9272 10696 10885 10724
rect 9272 10684 9278 10696
rect 10873 10693 10885 10696
rect 10919 10693 10931 10727
rect 12986 10724 12992 10736
rect 12947 10696 12992 10724
rect 10873 10687 10931 10693
rect 12986 10684 12992 10696
rect 13044 10684 13050 10736
rect 18230 10724 18236 10736
rect 18191 10696 18236 10724
rect 18230 10684 18236 10696
rect 18288 10684 18294 10736
rect 28629 10727 28687 10733
rect 28629 10693 28641 10727
rect 28675 10724 28687 10727
rect 32122 10724 32128 10736
rect 28675 10696 32128 10724
rect 28675 10693 28687 10696
rect 28629 10687 28687 10693
rect 32122 10684 32128 10696
rect 32180 10684 32186 10736
rect 3881 10659 3939 10665
rect 3881 10625 3893 10659
rect 3927 10625 3939 10659
rect 3881 10619 3939 10625
rect 4148 10659 4206 10665
rect 4148 10625 4160 10659
rect 4194 10656 4206 10659
rect 4706 10656 4712 10668
rect 4194 10628 4712 10656
rect 4194 10625 4206 10628
rect 4148 10619 4206 10625
rect 4706 10616 4712 10628
rect 4764 10656 4770 10668
rect 5166 10656 5172 10668
rect 4764 10628 5172 10656
rect 4764 10616 4770 10628
rect 5166 10616 5172 10628
rect 5224 10616 5230 10668
rect 5258 10616 5264 10668
rect 5316 10656 5322 10668
rect 9122 10656 9128 10668
rect 5316 10628 9128 10656
rect 5316 10616 5322 10628
rect 9122 10616 9128 10628
rect 9180 10616 9186 10668
rect 10042 10656 10048 10668
rect 10003 10628 10048 10656
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10656 10195 10659
rect 10410 10656 10416 10668
rect 10183 10628 10416 10656
rect 10183 10625 10195 10628
rect 10137 10619 10195 10625
rect 10410 10616 10416 10628
rect 10468 10616 10474 10668
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10656 10563 10659
rect 10962 10656 10968 10668
rect 10551 10628 10968 10656
rect 10551 10625 10563 10628
rect 10505 10619 10563 10625
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 9772 10600 9824 10606
rect 19978 10588 19984 10600
rect 19939 10560 19984 10588
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 9772 10542 9824 10548
rect 11057 10455 11115 10461
rect 11057 10421 11069 10455
rect 11103 10452 11115 10455
rect 11146 10452 11152 10464
rect 11103 10424 11152 10452
rect 11103 10421 11115 10424
rect 11057 10415 11115 10421
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 26418 10412 26424 10464
rect 26476 10452 26482 10464
rect 31110 10452 31116 10464
rect 26476 10424 31116 10452
rect 26476 10412 26482 10424
rect 31110 10412 31116 10424
rect 31168 10412 31174 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 5353 10251 5411 10257
rect 5353 10217 5365 10251
rect 5399 10248 5411 10251
rect 5442 10248 5448 10260
rect 5399 10220 5448 10248
rect 5399 10217 5411 10220
rect 5353 10211 5411 10217
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 10042 10208 10048 10260
rect 10100 10248 10106 10260
rect 10505 10251 10563 10257
rect 10505 10248 10517 10251
rect 10100 10220 10517 10248
rect 10100 10208 10106 10220
rect 10505 10217 10517 10220
rect 10551 10217 10563 10251
rect 10505 10211 10563 10217
rect 22002 10208 22008 10260
rect 22060 10248 22066 10260
rect 22097 10251 22155 10257
rect 22097 10248 22109 10251
rect 22060 10220 22109 10248
rect 22060 10208 22066 10220
rect 22097 10217 22109 10220
rect 22143 10217 22155 10251
rect 26694 10248 26700 10260
rect 22097 10211 22155 10217
rect 25056 10220 26556 10248
rect 26655 10220 26700 10248
rect 3970 10112 3976 10124
rect 3931 10084 3976 10112
rect 3970 10072 3976 10084
rect 4028 10072 4034 10124
rect 9122 10112 9128 10124
rect 9083 10084 9128 10112
rect 9122 10072 9128 10084
rect 9180 10072 9186 10124
rect 19334 10072 19340 10124
rect 19392 10112 19398 10124
rect 19392 10084 19932 10112
rect 19392 10072 19398 10084
rect 19242 10004 19248 10056
rect 19300 10044 19306 10056
rect 19904 10053 19932 10084
rect 21174 10072 21180 10124
rect 21232 10112 21238 10124
rect 25056 10112 25084 10220
rect 21232 10084 25084 10112
rect 26528 10112 26556 10220
rect 26694 10208 26700 10220
rect 26752 10208 26758 10260
rect 27982 10248 27988 10260
rect 27943 10220 27988 10248
rect 27982 10208 27988 10220
rect 28040 10208 28046 10260
rect 26528 10084 29960 10112
rect 21232 10072 21238 10084
rect 19613 10047 19671 10053
rect 19613 10044 19625 10047
rect 19300 10016 19625 10044
rect 19300 10004 19306 10016
rect 19613 10013 19625 10016
rect 19659 10013 19671 10047
rect 19613 10007 19671 10013
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10013 19947 10047
rect 19889 10007 19947 10013
rect 20809 10047 20867 10053
rect 20809 10013 20821 10047
rect 20855 10044 20867 10047
rect 24854 10044 24860 10056
rect 20855 10016 24860 10044
rect 20855 10013 20867 10016
rect 20809 10007 20867 10013
rect 4240 9979 4298 9985
rect 4240 9945 4252 9979
rect 4286 9976 4298 9979
rect 4706 9976 4712 9988
rect 4286 9948 4712 9976
rect 4286 9945 4298 9948
rect 4240 9939 4298 9945
rect 4706 9936 4712 9948
rect 4764 9936 4770 9988
rect 9214 9936 9220 9988
rect 9272 9976 9278 9988
rect 9398 9985 9404 9988
rect 9370 9979 9404 9985
rect 9370 9976 9382 9979
rect 9272 9948 9382 9976
rect 9272 9936 9278 9948
rect 9370 9945 9382 9948
rect 9456 9976 9462 9988
rect 9456 9948 9518 9976
rect 9370 9939 9404 9945
rect 9398 9936 9404 9939
rect 9456 9936 9462 9948
rect 19426 9908 19432 9920
rect 19387 9880 19432 9908
rect 19426 9868 19432 9880
rect 19484 9868 19490 9920
rect 19628 9908 19656 10007
rect 24854 10004 24860 10016
rect 24912 10004 24918 10056
rect 25056 10053 25084 10084
rect 25041 10047 25099 10053
rect 25041 10013 25053 10047
rect 25087 10013 25099 10047
rect 25222 10044 25228 10056
rect 25183 10016 25228 10044
rect 25041 10007 25099 10013
rect 25222 10004 25228 10016
rect 25280 10004 25286 10056
rect 25314 10004 25320 10056
rect 25372 10044 25378 10056
rect 25372 10016 25417 10044
rect 25372 10004 25378 10016
rect 25958 10004 25964 10056
rect 26016 10044 26022 10056
rect 26145 10047 26203 10053
rect 26145 10044 26157 10047
rect 26016 10016 26157 10044
rect 26016 10004 26022 10016
rect 26145 10013 26157 10016
rect 26191 10013 26203 10047
rect 26418 10044 26424 10056
rect 26379 10016 26424 10044
rect 26145 10007 26203 10013
rect 26418 10004 26424 10016
rect 26476 10004 26482 10056
rect 26510 10004 26516 10056
rect 26568 10044 26574 10056
rect 26568 10016 26613 10044
rect 26568 10004 26574 10016
rect 29086 10004 29092 10056
rect 29144 10044 29150 10056
rect 29932 10053 29960 10084
rect 30208 10084 31156 10112
rect 30208 10056 30236 10084
rect 29917 10047 29975 10053
rect 29144 10016 29868 10044
rect 29144 10004 29150 10016
rect 19797 9979 19855 9985
rect 19797 9945 19809 9979
rect 19843 9976 19855 9979
rect 20162 9976 20168 9988
rect 19843 9948 20168 9976
rect 19843 9945 19855 9948
rect 19797 9939 19855 9945
rect 20162 9936 20168 9948
rect 20220 9936 20226 9988
rect 25406 9936 25412 9988
rect 25464 9976 25470 9988
rect 26050 9976 26056 9988
rect 25464 9948 26056 9976
rect 25464 9936 25470 9948
rect 26050 9936 26056 9948
rect 26108 9976 26114 9988
rect 26329 9979 26387 9985
rect 26329 9976 26341 9979
rect 26108 9948 26341 9976
rect 26108 9936 26114 9948
rect 26329 9945 26341 9948
rect 26375 9945 26387 9979
rect 26329 9939 26387 9945
rect 21174 9908 21180 9920
rect 19628 9880 21180 9908
rect 21174 9868 21180 9880
rect 21232 9868 21238 9920
rect 24854 9908 24860 9920
rect 24815 9880 24860 9908
rect 24854 9868 24860 9880
rect 24912 9868 24918 9920
rect 26528 9908 26556 10004
rect 27614 9936 27620 9988
rect 27672 9976 27678 9988
rect 27801 9979 27859 9985
rect 27801 9976 27813 9979
rect 27672 9948 27813 9976
rect 27672 9936 27678 9948
rect 27801 9945 27813 9948
rect 27847 9976 27859 9979
rect 28258 9976 28264 9988
rect 27847 9948 28264 9976
rect 27847 9945 27859 9948
rect 27801 9939 27859 9945
rect 28258 9936 28264 9948
rect 28316 9936 28322 9988
rect 28994 9936 29000 9988
rect 29052 9976 29058 9988
rect 29733 9979 29791 9985
rect 29733 9976 29745 9979
rect 29052 9948 29745 9976
rect 29052 9936 29058 9948
rect 29733 9945 29745 9948
rect 29779 9945 29791 9979
rect 29840 9976 29868 10016
rect 29917 10013 29929 10047
rect 29963 10013 29975 10047
rect 30190 10044 30196 10056
rect 30151 10016 30196 10044
rect 29917 10007 29975 10013
rect 30190 10004 30196 10016
rect 30248 10004 30254 10056
rect 30466 10004 30472 10056
rect 30524 10044 30530 10056
rect 31128 10053 31156 10084
rect 30837 10047 30895 10053
rect 30837 10044 30849 10047
rect 30524 10016 30849 10044
rect 30524 10004 30530 10016
rect 30837 10013 30849 10016
rect 30883 10013 30895 10047
rect 30837 10007 30895 10013
rect 31113 10047 31171 10053
rect 31113 10013 31125 10047
rect 31159 10013 31171 10047
rect 31113 10007 31171 10013
rect 30101 9979 30159 9985
rect 30101 9976 30113 9979
rect 29840 9948 30113 9976
rect 29733 9939 29791 9945
rect 30101 9945 30113 9948
rect 30147 9945 30159 9979
rect 30101 9939 30159 9945
rect 30282 9936 30288 9988
rect 30340 9976 30346 9988
rect 31021 9979 31079 9985
rect 31021 9976 31033 9979
rect 30340 9948 31033 9976
rect 30340 9936 30346 9948
rect 31021 9945 31033 9948
rect 31067 9945 31079 9979
rect 31021 9939 31079 9945
rect 27985 9911 28043 9917
rect 27985 9908 27997 9911
rect 26528 9880 27997 9908
rect 27985 9877 27997 9880
rect 28031 9877 28043 9911
rect 27985 9871 28043 9877
rect 28169 9911 28227 9917
rect 28169 9877 28181 9911
rect 28215 9908 28227 9911
rect 29638 9908 29644 9920
rect 28215 9880 29644 9908
rect 28215 9877 28227 9880
rect 28169 9871 28227 9877
rect 29638 9868 29644 9880
rect 29696 9868 29702 9920
rect 30650 9908 30656 9920
rect 30611 9880 30656 9908
rect 30650 9868 30656 9880
rect 30708 9868 30714 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 11146 9664 11152 9716
rect 11204 9704 11210 9716
rect 17218 9704 17224 9716
rect 11204 9676 17224 9704
rect 11204 9664 11210 9676
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 20073 9707 20131 9713
rect 20073 9673 20085 9707
rect 20119 9704 20131 9707
rect 20162 9704 20168 9716
rect 20119 9676 20168 9704
rect 20119 9673 20131 9676
rect 20073 9667 20131 9673
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 20530 9664 20536 9716
rect 20588 9704 20594 9716
rect 20588 9676 20760 9704
rect 20588 9664 20594 9676
rect 15562 9636 15568 9648
rect 15523 9608 15568 9636
rect 15562 9596 15568 9608
rect 15620 9596 15626 9648
rect 18960 9639 19018 9645
rect 18960 9605 18972 9639
rect 19006 9636 19018 9639
rect 19426 9636 19432 9648
rect 19006 9608 19432 9636
rect 19006 9605 19018 9608
rect 18960 9599 19018 9605
rect 19426 9596 19432 9608
rect 19484 9596 19490 9648
rect 20438 9596 20444 9648
rect 20496 9636 20502 9648
rect 20640 9636 20668 9676
rect 20732 9645 20760 9676
rect 29086 9664 29092 9716
rect 29144 9704 29150 9716
rect 29181 9707 29239 9713
rect 29181 9704 29193 9707
rect 29144 9676 29193 9704
rect 29144 9664 29150 9676
rect 29181 9673 29193 9676
rect 29227 9673 29239 9707
rect 29181 9667 29239 9673
rect 20496 9608 20668 9636
rect 20717 9639 20775 9645
rect 20496 9596 20502 9608
rect 20717 9605 20729 9639
rect 20763 9636 20775 9639
rect 25406 9636 25412 9648
rect 20763 9608 20797 9636
rect 25367 9608 25412 9636
rect 20763 9605 20775 9608
rect 20717 9599 20775 9605
rect 25406 9596 25412 9608
rect 25464 9596 25470 9648
rect 25501 9639 25559 9645
rect 25501 9605 25513 9639
rect 25547 9636 25559 9639
rect 27706 9636 27712 9648
rect 25547 9608 27712 9636
rect 25547 9605 25559 9608
rect 25501 9599 25559 9605
rect 27706 9596 27712 9608
rect 27764 9596 27770 9648
rect 28994 9636 29000 9648
rect 28184 9608 29000 9636
rect 2685 9571 2743 9577
rect 2685 9537 2697 9571
rect 2731 9568 2743 9571
rect 2958 9568 2964 9580
rect 2731 9540 2964 9568
rect 2731 9537 2743 9540
rect 2685 9531 2743 9537
rect 2958 9528 2964 9540
rect 3016 9528 3022 9580
rect 12986 9568 12992 9580
rect 12947 9540 12992 9568
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 15286 9528 15292 9580
rect 15344 9568 15350 9580
rect 15381 9571 15439 9577
rect 15381 9568 15393 9571
rect 15344 9540 15393 9568
rect 15344 9528 15350 9540
rect 15381 9537 15393 9540
rect 15427 9537 15439 9571
rect 15381 9531 15439 9537
rect 15396 9500 15424 9531
rect 15470 9528 15476 9580
rect 15528 9568 15534 9580
rect 15657 9571 15715 9577
rect 15657 9568 15669 9571
rect 15528 9540 15669 9568
rect 15528 9528 15534 9540
rect 15657 9537 15669 9540
rect 15703 9568 15715 9571
rect 16482 9568 16488 9580
rect 15703 9540 16488 9568
rect 15703 9537 15715 9540
rect 15657 9531 15715 9537
rect 16482 9528 16488 9540
rect 16540 9528 16546 9580
rect 19242 9568 19248 9580
rect 18616 9540 19248 9568
rect 18616 9500 18644 9540
rect 19242 9528 19248 9540
rect 19300 9528 19306 9580
rect 20530 9568 20536 9580
rect 20491 9540 20536 9568
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 20805 9571 20863 9577
rect 20805 9537 20817 9571
rect 20851 9537 20863 9571
rect 20805 9531 20863 9537
rect 15396 9472 18644 9500
rect 18693 9503 18751 9509
rect 18693 9469 18705 9503
rect 18739 9469 18751 9503
rect 18693 9463 18751 9469
rect 1854 9324 1860 9376
rect 1912 9364 1918 9376
rect 2777 9367 2835 9373
rect 2777 9364 2789 9367
rect 1912 9336 2789 9364
rect 1912 9324 1918 9336
rect 2777 9333 2789 9336
rect 2823 9333 2835 9367
rect 14274 9364 14280 9376
rect 14235 9336 14280 9364
rect 2777 9327 2835 9333
rect 14274 9324 14280 9336
rect 14332 9324 14338 9376
rect 15194 9364 15200 9376
rect 15155 9336 15200 9364
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 18708 9364 18736 9463
rect 20824 9444 20852 9531
rect 20898 9528 20904 9580
rect 20956 9568 20962 9580
rect 25225 9571 25283 9577
rect 20956 9540 21001 9568
rect 20956 9528 20962 9540
rect 25225 9537 25237 9571
rect 25271 9537 25283 9571
rect 25225 9531 25283 9537
rect 25593 9571 25651 9577
rect 25593 9537 25605 9571
rect 25639 9568 25651 9571
rect 26510 9568 26516 9580
rect 25639 9540 26516 9568
rect 25639 9537 25651 9540
rect 25593 9531 25651 9537
rect 25240 9500 25268 9531
rect 26510 9528 26516 9540
rect 26568 9528 26574 9580
rect 27801 9571 27859 9577
rect 27801 9537 27813 9571
rect 27847 9537 27859 9571
rect 27801 9531 27859 9537
rect 28068 9571 28126 9577
rect 28068 9537 28080 9571
rect 28114 9568 28126 9571
rect 28184 9568 28212 9608
rect 28994 9596 29000 9608
rect 29052 9596 29058 9648
rect 29638 9636 29644 9648
rect 29599 9608 29644 9636
rect 29638 9596 29644 9608
rect 29696 9596 29702 9648
rect 28114 9540 28212 9568
rect 28114 9537 28126 9540
rect 28068 9531 28126 9537
rect 26142 9500 26148 9512
rect 25240 9472 26148 9500
rect 26142 9460 26148 9472
rect 26200 9460 26206 9512
rect 20806 9392 20812 9444
rect 20864 9392 20870 9444
rect 21082 9432 21088 9444
rect 21043 9404 21088 9432
rect 21082 9392 21088 9404
rect 21140 9392 21146 9444
rect 19334 9364 19340 9376
rect 18708 9336 19340 9364
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 20254 9324 20260 9376
rect 20312 9364 20318 9376
rect 25777 9367 25835 9373
rect 25777 9364 25789 9367
rect 20312 9336 25789 9364
rect 20312 9324 20318 9336
rect 25777 9333 25789 9336
rect 25823 9333 25835 9367
rect 27816 9364 27844 9531
rect 28810 9392 28816 9444
rect 28868 9432 28874 9444
rect 30929 9435 30987 9441
rect 30929 9432 30941 9435
rect 28868 9404 30941 9432
rect 28868 9392 28874 9404
rect 30929 9401 30941 9404
rect 30975 9401 30987 9435
rect 30929 9395 30987 9401
rect 29730 9364 29736 9376
rect 27816 9336 29736 9364
rect 25777 9327 25835 9333
rect 29730 9324 29736 9336
rect 29788 9324 29794 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 2958 9120 2964 9172
rect 3016 9160 3022 9172
rect 3329 9163 3387 9169
rect 3329 9160 3341 9163
rect 3016 9132 3341 9160
rect 3016 9120 3022 9132
rect 3329 9129 3341 9132
rect 3375 9160 3387 9163
rect 4062 9160 4068 9172
rect 3375 9132 4068 9160
rect 3375 9129 3387 9132
rect 3329 9123 3387 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 15657 9163 15715 9169
rect 15657 9129 15669 9163
rect 15703 9160 15715 9163
rect 16390 9160 16396 9172
rect 15703 9132 16396 9160
rect 15703 9129 15715 9132
rect 15657 9123 15715 9129
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 18598 9160 18604 9172
rect 16592 9132 18604 9160
rect 16482 9052 16488 9104
rect 16540 9092 16546 9104
rect 16592 9092 16620 9132
rect 18598 9120 18604 9132
rect 18656 9120 18662 9172
rect 18693 9163 18751 9169
rect 18693 9129 18705 9163
rect 18739 9160 18751 9163
rect 18966 9160 18972 9172
rect 18739 9132 18972 9160
rect 18739 9129 18751 9132
rect 18693 9123 18751 9129
rect 18966 9120 18972 9132
rect 19024 9120 19030 9172
rect 20438 9120 20444 9172
rect 20496 9160 20502 9172
rect 23566 9160 23572 9172
rect 20496 9132 20852 9160
rect 23527 9132 23572 9160
rect 20496 9120 20502 9132
rect 16540 9064 16620 9092
rect 20824 9092 20852 9132
rect 23566 9120 23572 9132
rect 23624 9120 23630 9172
rect 25222 9120 25228 9172
rect 25280 9160 25286 9172
rect 25961 9163 26019 9169
rect 25961 9160 25973 9163
rect 25280 9132 25973 9160
rect 25280 9120 25286 9132
rect 25961 9129 25973 9132
rect 26007 9129 26019 9163
rect 25961 9123 26019 9129
rect 27706 9120 27712 9172
rect 27764 9160 27770 9172
rect 29181 9163 29239 9169
rect 29181 9160 29193 9163
rect 27764 9132 29193 9160
rect 27764 9120 27770 9132
rect 29181 9129 29193 9132
rect 29227 9160 29239 9163
rect 30926 9160 30932 9172
rect 29227 9132 30932 9160
rect 29227 9129 29239 9132
rect 29181 9123 29239 9129
rect 30926 9120 30932 9132
rect 30984 9120 30990 9172
rect 31110 9160 31116 9172
rect 31071 9132 31116 9160
rect 31110 9120 31116 9132
rect 31168 9120 31174 9172
rect 20824 9064 23612 9092
rect 16540 9052 16546 9064
rect 1854 9024 1860 9036
rect 1815 8996 1860 9024
rect 1854 8984 1860 8996
rect 1912 8984 1918 9036
rect 14274 9024 14280 9036
rect 14235 8996 14280 9024
rect 14274 8984 14280 8996
rect 14332 8984 14338 9036
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 2958 8916 2964 8968
rect 3016 8916 3022 8968
rect 16298 8956 16304 8968
rect 16259 8928 16304 8956
rect 16298 8916 16304 8928
rect 16356 8916 16362 8968
rect 16390 8916 16396 8968
rect 16448 8956 16454 8968
rect 16592 8965 16620 9064
rect 18874 9024 18880 9036
rect 18156 8996 18880 9024
rect 18156 8965 18184 8996
rect 18874 8984 18880 8996
rect 18932 8984 18938 9036
rect 18984 8996 22140 9024
rect 16485 8959 16543 8965
rect 16485 8956 16497 8959
rect 16448 8928 16497 8956
rect 16448 8916 16454 8928
rect 16485 8925 16497 8928
rect 16531 8925 16543 8959
rect 16485 8919 16543 8925
rect 16577 8959 16635 8965
rect 16577 8925 16589 8959
rect 16623 8925 16635 8959
rect 16577 8919 16635 8925
rect 18141 8959 18199 8965
rect 18141 8925 18153 8959
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 18230 8916 18236 8968
rect 18288 8956 18294 8968
rect 18506 8956 18512 8968
rect 18288 8928 18512 8956
rect 18288 8916 18294 8928
rect 18506 8916 18512 8928
rect 18564 8916 18570 8968
rect 18598 8916 18604 8968
rect 18656 8956 18662 8968
rect 18984 8956 19012 8996
rect 18656 8928 19012 8956
rect 21821 8959 21879 8965
rect 18656 8916 18662 8928
rect 21821 8925 21833 8959
rect 21867 8956 21879 8959
rect 21910 8956 21916 8968
rect 21867 8928 21916 8956
rect 21867 8925 21879 8928
rect 21821 8919 21879 8925
rect 21910 8916 21916 8928
rect 21968 8916 21974 8968
rect 22112 8965 22140 8996
rect 22097 8959 22155 8965
rect 22097 8925 22109 8959
rect 22143 8925 22155 8959
rect 22097 8919 22155 8925
rect 14544 8891 14602 8897
rect 14544 8857 14556 8891
rect 14590 8888 14602 8891
rect 16117 8891 16175 8897
rect 16117 8888 16129 8891
rect 14590 8860 16129 8888
rect 14590 8857 14602 8860
rect 14544 8851 14602 8857
rect 16117 8857 16129 8860
rect 16163 8857 16175 8891
rect 18322 8888 18328 8900
rect 18283 8860 18328 8888
rect 16117 8851 16175 8857
rect 18322 8848 18328 8860
rect 18380 8848 18386 8900
rect 18417 8891 18475 8897
rect 18417 8857 18429 8891
rect 18463 8857 18475 8891
rect 19426 8888 19432 8900
rect 19387 8860 19432 8888
rect 18417 8851 18475 8857
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 5626 8820 5632 8832
rect 2832 8792 5632 8820
rect 2832 8780 2838 8792
rect 5626 8780 5632 8792
rect 5684 8820 5690 8832
rect 6730 8820 6736 8832
rect 5684 8792 6736 8820
rect 5684 8780 5690 8792
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 16666 8780 16672 8832
rect 16724 8820 16730 8832
rect 18432 8820 18460 8851
rect 19426 8848 19432 8860
rect 19484 8848 19490 8900
rect 19978 8848 19984 8900
rect 20036 8888 20042 8900
rect 22186 8888 22192 8900
rect 20036 8860 22192 8888
rect 20036 8848 20042 8860
rect 22186 8848 22192 8860
rect 22244 8888 22250 8900
rect 23382 8888 23388 8900
rect 22244 8860 23388 8888
rect 22244 8848 22250 8860
rect 23382 8848 23388 8860
rect 23440 8848 23446 8900
rect 23584 8897 23612 9064
rect 24578 8956 24584 8968
rect 24539 8928 24584 8956
rect 24578 8916 24584 8928
rect 24636 8916 24642 8968
rect 24854 8965 24860 8968
rect 24848 8956 24860 8965
rect 24815 8928 24860 8956
rect 24848 8919 24860 8928
rect 24854 8916 24860 8919
rect 24912 8916 24918 8968
rect 27801 8959 27859 8965
rect 27801 8925 27813 8959
rect 27847 8956 27859 8959
rect 29086 8956 29092 8968
rect 27847 8928 29092 8956
rect 27847 8925 27859 8928
rect 27801 8919 27859 8925
rect 29086 8916 29092 8928
rect 29144 8916 29150 8968
rect 29730 8956 29736 8968
rect 29691 8928 29736 8956
rect 29730 8916 29736 8928
rect 29788 8916 29794 8968
rect 23569 8891 23627 8897
rect 23569 8857 23581 8891
rect 23615 8888 23627 8891
rect 25406 8888 25412 8900
rect 23615 8860 25412 8888
rect 23615 8857 23627 8860
rect 23569 8851 23627 8857
rect 25406 8848 25412 8860
rect 25464 8848 25470 8900
rect 28068 8891 28126 8897
rect 28068 8857 28080 8891
rect 28114 8888 28126 8891
rect 29638 8888 29644 8900
rect 28114 8860 29644 8888
rect 28114 8857 28126 8860
rect 28068 8851 28126 8857
rect 29638 8848 29644 8860
rect 29696 8848 29702 8900
rect 29822 8848 29828 8900
rect 29880 8888 29886 8900
rect 29978 8891 30036 8897
rect 29978 8888 29990 8891
rect 29880 8860 29990 8888
rect 29880 8848 29886 8860
rect 29978 8857 29990 8860
rect 30024 8857 30036 8891
rect 29978 8851 30036 8857
rect 16724 8792 18460 8820
rect 16724 8780 16730 8792
rect 20070 8780 20076 8832
rect 20128 8820 20134 8832
rect 20717 8823 20775 8829
rect 20717 8820 20729 8823
rect 20128 8792 20729 8820
rect 20128 8780 20134 8792
rect 20717 8789 20729 8792
rect 20763 8789 20775 8823
rect 21634 8820 21640 8832
rect 21595 8792 21640 8820
rect 20717 8783 20775 8789
rect 21634 8780 21640 8792
rect 21692 8780 21698 8832
rect 22002 8820 22008 8832
rect 21963 8792 22008 8820
rect 22002 8780 22008 8792
rect 22060 8780 22066 8832
rect 23753 8823 23811 8829
rect 23753 8789 23765 8823
rect 23799 8820 23811 8823
rect 24670 8820 24676 8832
rect 23799 8792 24676 8820
rect 23799 8789 23811 8792
rect 23753 8783 23811 8789
rect 24670 8780 24676 8792
rect 24728 8780 24734 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1578 8576 1584 8628
rect 1636 8616 1642 8628
rect 5534 8616 5540 8628
rect 1636 8588 5540 8616
rect 1636 8576 1642 8588
rect 2700 8489 2728 8588
rect 5534 8576 5540 8588
rect 5592 8616 5598 8628
rect 13909 8619 13967 8625
rect 5592 8588 6592 8616
rect 5592 8576 5598 8588
rect 2958 8548 2964 8560
rect 2919 8520 2964 8548
rect 2958 8508 2964 8520
rect 3016 8508 3022 8560
rect 4884 8551 4942 8557
rect 4884 8517 4896 8551
rect 4930 8548 4942 8551
rect 5350 8548 5356 8560
rect 4930 8520 5356 8548
rect 4930 8517 4942 8520
rect 4884 8511 4942 8517
rect 5350 8508 5356 8520
rect 5408 8508 5414 8560
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 4614 8480 4620 8492
rect 2832 8452 2877 8480
rect 4575 8452 4620 8480
rect 2832 8440 2838 8452
rect 4614 8440 4620 8452
rect 4672 8480 4678 8492
rect 5442 8480 5448 8492
rect 4672 8452 5448 8480
rect 4672 8440 4678 8452
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 6564 8489 6592 8588
rect 13909 8585 13921 8619
rect 13955 8616 13967 8619
rect 15746 8616 15752 8628
rect 13955 8588 15752 8616
rect 13955 8585 13967 8588
rect 13909 8579 13967 8585
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 17037 8619 17095 8625
rect 17037 8585 17049 8619
rect 17083 8616 17095 8619
rect 18230 8616 18236 8628
rect 17083 8588 18236 8616
rect 17083 8585 17095 8588
rect 17037 8579 17095 8585
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 18693 8619 18751 8625
rect 18693 8585 18705 8619
rect 18739 8616 18751 8619
rect 19426 8616 19432 8628
rect 18739 8588 19432 8616
rect 18739 8585 18751 8588
rect 18693 8579 18751 8585
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 20346 8576 20352 8628
rect 20404 8616 20410 8628
rect 20625 8619 20683 8625
rect 20625 8616 20637 8619
rect 20404 8588 20637 8616
rect 20404 8576 20410 8588
rect 20625 8585 20637 8588
rect 20671 8616 20683 8619
rect 22002 8616 22008 8628
rect 20671 8588 22008 8616
rect 20671 8585 20683 8588
rect 20625 8579 20683 8585
rect 22002 8576 22008 8588
rect 22060 8576 22066 8628
rect 23382 8576 23388 8628
rect 23440 8616 23446 8628
rect 25961 8619 26019 8625
rect 25961 8616 25973 8619
rect 23440 8588 25973 8616
rect 23440 8576 23446 8588
rect 25961 8585 25973 8588
rect 26007 8585 26019 8619
rect 25961 8579 26019 8585
rect 29638 8576 29644 8628
rect 29696 8616 29702 8628
rect 30561 8619 30619 8625
rect 30561 8616 30573 8619
rect 29696 8588 30573 8616
rect 29696 8576 29702 8588
rect 30561 8585 30573 8588
rect 30607 8585 30619 8619
rect 30926 8616 30932 8628
rect 30887 8588 30932 8616
rect 30561 8579 30619 8585
rect 30926 8576 30932 8588
rect 30984 8576 30990 8628
rect 10965 8551 11023 8557
rect 10965 8517 10977 8551
rect 11011 8548 11023 8551
rect 12710 8548 12716 8560
rect 11011 8520 12716 8548
rect 11011 8517 11023 8520
rect 10965 8511 11023 8517
rect 12710 8508 12716 8520
rect 12768 8508 12774 8560
rect 14016 8520 14872 8548
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8449 6607 8483
rect 6730 8480 6736 8492
rect 6691 8452 6736 8480
rect 6549 8443 6607 8449
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 10137 8483 10195 8489
rect 10137 8449 10149 8483
rect 10183 8480 10195 8483
rect 10870 8480 10876 8492
rect 10183 8452 10876 8480
rect 10183 8449 10195 8452
rect 10137 8443 10195 8449
rect 10870 8440 10876 8452
rect 10928 8440 10934 8492
rect 13446 8440 13452 8492
rect 13504 8480 13510 8492
rect 14016 8489 14044 8520
rect 13725 8483 13783 8489
rect 13725 8480 13737 8483
rect 13504 8452 13737 8480
rect 13504 8440 13510 8452
rect 13725 8449 13737 8452
rect 13771 8449 13783 8483
rect 13725 8443 13783 8449
rect 14001 8483 14059 8489
rect 14001 8449 14013 8483
rect 14047 8449 14059 8483
rect 14001 8443 14059 8449
rect 14461 8483 14519 8489
rect 14461 8449 14473 8483
rect 14507 8480 14519 8483
rect 14734 8480 14740 8492
rect 14507 8452 14740 8480
rect 14507 8449 14519 8452
rect 14461 8443 14519 8449
rect 14734 8440 14740 8452
rect 14792 8440 14798 8492
rect 8294 8372 8300 8424
rect 8352 8412 8358 8424
rect 10045 8415 10103 8421
rect 10045 8412 10057 8415
rect 8352 8384 10057 8412
rect 8352 8372 8358 8384
rect 10045 8381 10057 8384
rect 10091 8381 10103 8415
rect 10045 8375 10103 8381
rect 10226 8372 10232 8424
rect 10284 8412 10290 8424
rect 10594 8412 10600 8424
rect 10284 8384 10600 8412
rect 10284 8372 10290 8384
rect 10594 8372 10600 8384
rect 10652 8372 10658 8424
rect 13541 8415 13599 8421
rect 13541 8381 13553 8415
rect 13587 8412 13599 8415
rect 14642 8412 14648 8424
rect 13587 8384 14648 8412
rect 13587 8381 13599 8384
rect 13541 8375 13599 8381
rect 14642 8372 14648 8384
rect 14700 8372 14706 8424
rect 14844 8412 14872 8520
rect 15102 8508 15108 8560
rect 15160 8548 15166 8560
rect 16853 8551 16911 8557
rect 16853 8548 16865 8551
rect 15160 8520 16865 8548
rect 15160 8508 15166 8520
rect 16853 8517 16865 8520
rect 16899 8517 16911 8551
rect 16853 8511 16911 8517
rect 17862 8508 17868 8560
rect 17920 8548 17926 8560
rect 18325 8551 18383 8557
rect 18325 8548 18337 8551
rect 17920 8520 18337 8548
rect 17920 8508 17926 8520
rect 18325 8517 18337 8520
rect 18371 8517 18383 8551
rect 18325 8511 18383 8517
rect 18414 8508 18420 8560
rect 18472 8548 18478 8560
rect 18509 8551 18567 8557
rect 18509 8548 18521 8551
rect 18472 8520 18521 8548
rect 18472 8508 18478 8520
rect 18509 8517 18521 8520
rect 18555 8548 18567 8551
rect 19512 8551 19570 8557
rect 18555 8520 19472 8548
rect 18555 8517 18567 8520
rect 18509 8511 18567 8517
rect 14918 8440 14924 8492
rect 14976 8480 14982 8492
rect 17313 8483 17371 8489
rect 17313 8480 17325 8483
rect 14976 8452 17325 8480
rect 14976 8440 14982 8452
rect 17313 8449 17325 8452
rect 17359 8449 17371 8483
rect 17313 8443 17371 8449
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8480 19303 8483
rect 19334 8480 19340 8492
rect 19291 8452 19340 8480
rect 19291 8449 19303 8452
rect 19245 8443 19303 8449
rect 19334 8440 19340 8452
rect 19392 8440 19398 8492
rect 19444 8480 19472 8520
rect 19512 8517 19524 8551
rect 19558 8548 19570 8551
rect 21634 8548 21640 8560
rect 19558 8520 21640 8548
rect 19558 8517 19570 8520
rect 19512 8511 19570 8517
rect 21634 8508 21640 8520
rect 21692 8508 21698 8560
rect 24486 8548 24492 8560
rect 22848 8520 24492 8548
rect 20898 8480 20904 8492
rect 19444 8452 20904 8480
rect 20898 8440 20904 8452
rect 20956 8440 20962 8492
rect 22848 8489 22876 8520
rect 24486 8508 24492 8520
rect 24544 8508 24550 8560
rect 24670 8548 24676 8560
rect 24631 8520 24676 8548
rect 24670 8508 24676 8520
rect 24728 8508 24734 8560
rect 29086 8548 29092 8560
rect 28736 8520 29092 8548
rect 22833 8483 22891 8489
rect 22833 8449 22845 8483
rect 22879 8449 22891 8483
rect 22833 8443 22891 8449
rect 22922 8440 22928 8492
rect 22980 8480 22986 8492
rect 28736 8489 28764 8520
rect 29086 8508 29092 8520
rect 29144 8548 29150 8560
rect 29914 8548 29920 8560
rect 29144 8520 29920 8548
rect 29144 8508 29150 8520
rect 29914 8508 29920 8520
rect 29972 8508 29978 8560
rect 30190 8508 30196 8560
rect 30248 8548 30254 8560
rect 30248 8520 31064 8548
rect 30248 8508 30254 8520
rect 23089 8483 23147 8489
rect 23089 8480 23101 8483
rect 22980 8452 23101 8480
rect 22980 8440 22986 8452
rect 23089 8449 23101 8452
rect 23135 8449 23147 8483
rect 23089 8443 23147 8449
rect 28721 8483 28779 8489
rect 28721 8449 28733 8483
rect 28767 8449 28779 8483
rect 28721 8443 28779 8449
rect 28988 8483 29046 8489
rect 28988 8449 29000 8483
rect 29034 8480 29046 8483
rect 30650 8480 30656 8492
rect 29034 8452 30656 8480
rect 29034 8449 29046 8452
rect 28988 8443 29046 8449
rect 30650 8440 30656 8452
rect 30708 8440 30714 8492
rect 30742 8440 30748 8492
rect 30800 8480 30806 8492
rect 31036 8489 31064 8520
rect 31021 8483 31079 8489
rect 30800 8452 30845 8480
rect 30800 8440 30806 8452
rect 31021 8449 31033 8483
rect 31067 8449 31079 8483
rect 31021 8443 31079 8449
rect 15286 8412 15292 8424
rect 14844 8384 15292 8412
rect 15286 8372 15292 8384
rect 15344 8412 15350 8424
rect 16482 8412 16488 8424
rect 15344 8384 16488 8412
rect 15344 8372 15350 8384
rect 16482 8372 16488 8384
rect 16540 8372 16546 8424
rect 30760 8412 30788 8440
rect 32490 8412 32496 8424
rect 30760 8384 32496 8412
rect 32490 8372 32496 8384
rect 32548 8372 32554 8424
rect 5997 8347 6055 8353
rect 5997 8313 6009 8347
rect 6043 8344 6055 8347
rect 7006 8344 7012 8356
rect 6043 8316 7012 8344
rect 6043 8313 6055 8316
rect 5997 8307 6055 8313
rect 7006 8304 7012 8316
rect 7064 8304 7070 8356
rect 10134 8304 10140 8356
rect 10192 8344 10198 8356
rect 10505 8347 10563 8353
rect 10505 8344 10517 8347
rect 10192 8316 10517 8344
rect 10192 8304 10198 8316
rect 10505 8313 10517 8316
rect 10551 8313 10563 8347
rect 10505 8307 10563 8313
rect 12986 8304 12992 8356
rect 13044 8344 13050 8356
rect 15749 8347 15807 8353
rect 15749 8344 15761 8347
rect 13044 8316 15761 8344
rect 13044 8304 13050 8316
rect 15749 8313 15761 8316
rect 15795 8313 15807 8347
rect 15749 8307 15807 8313
rect 16298 8304 16304 8356
rect 16356 8344 16362 8356
rect 30101 8347 30159 8353
rect 16356 8316 19288 8344
rect 16356 8304 16362 8316
rect 6546 8236 6552 8288
rect 6604 8276 6610 8288
rect 6641 8279 6699 8285
rect 6641 8276 6653 8279
rect 6604 8248 6653 8276
rect 6604 8236 6610 8248
rect 6641 8245 6653 8248
rect 6687 8245 6699 8279
rect 6641 8239 6699 8245
rect 12618 8236 12624 8288
rect 12676 8276 12682 8288
rect 17037 8279 17095 8285
rect 17037 8276 17049 8279
rect 12676 8248 17049 8276
rect 12676 8236 12682 8248
rect 17037 8245 17049 8248
rect 17083 8276 17095 8279
rect 18506 8276 18512 8288
rect 17083 8248 18512 8276
rect 17083 8245 17095 8248
rect 17037 8239 17095 8245
rect 18506 8236 18512 8248
rect 18564 8236 18570 8288
rect 19260 8276 19288 8316
rect 30101 8313 30113 8347
rect 30147 8344 30159 8347
rect 30282 8344 30288 8356
rect 30147 8316 30288 8344
rect 30147 8313 30159 8316
rect 30101 8307 30159 8313
rect 30282 8304 30288 8316
rect 30340 8304 30346 8356
rect 20622 8276 20628 8288
rect 19260 8248 20628 8276
rect 20622 8236 20628 8248
rect 20680 8236 20686 8288
rect 20714 8236 20720 8288
rect 20772 8276 20778 8288
rect 23106 8276 23112 8288
rect 20772 8248 23112 8276
rect 20772 8236 20778 8248
rect 23106 8236 23112 8248
rect 23164 8236 23170 8288
rect 23198 8236 23204 8288
rect 23256 8276 23262 8288
rect 24213 8279 24271 8285
rect 24213 8276 24225 8279
rect 23256 8248 24225 8276
rect 23256 8236 23262 8248
rect 24213 8245 24225 8248
rect 24259 8245 24271 8279
rect 24213 8239 24271 8245
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 6914 8072 6920 8084
rect 6827 8044 6920 8072
rect 6914 8032 6920 8044
rect 6972 8072 6978 8084
rect 8294 8072 8300 8084
rect 6972 8044 8300 8072
rect 6972 8032 6978 8044
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 10870 8072 10876 8084
rect 10831 8044 10876 8072
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 12710 8072 12716 8084
rect 12406 8044 12716 8072
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7936 5227 7939
rect 8938 7936 8944 7948
rect 5215 7908 8944 7936
rect 5215 7905 5227 7908
rect 5169 7899 5227 7905
rect 8938 7896 8944 7908
rect 8996 7936 9002 7948
rect 9125 7939 9183 7945
rect 9125 7936 9137 7939
rect 8996 7908 9137 7936
rect 8996 7896 9002 7908
rect 9125 7905 9137 7908
rect 9171 7905 9183 7939
rect 9125 7899 9183 7905
rect 9401 7939 9459 7945
rect 9401 7905 9413 7939
rect 9447 7936 9459 7939
rect 9490 7936 9496 7948
rect 9447 7908 9496 7936
rect 9447 7905 9459 7908
rect 9401 7899 9459 7905
rect 9490 7896 9496 7908
rect 9548 7896 9554 7948
rect 12406 7936 12434 8044
rect 12710 8032 12716 8044
rect 12768 8072 12774 8084
rect 15102 8072 15108 8084
rect 12768 8044 15108 8072
rect 12768 8032 12774 8044
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 15562 8032 15568 8084
rect 15620 8072 15626 8084
rect 15841 8075 15899 8081
rect 15841 8072 15853 8075
rect 15620 8044 15853 8072
rect 15620 8032 15626 8044
rect 15841 8041 15853 8044
rect 15887 8041 15899 8075
rect 15841 8035 15899 8041
rect 18506 8032 18512 8084
rect 18564 8072 18570 8084
rect 20806 8072 20812 8084
rect 18564 8044 20668 8072
rect 20767 8044 20812 8072
rect 18564 8032 18570 8044
rect 16482 7964 16488 8016
rect 16540 7964 16546 8016
rect 20640 8004 20668 8044
rect 20806 8032 20812 8044
rect 20864 8032 20870 8084
rect 22833 8075 22891 8081
rect 22833 8041 22845 8075
rect 22879 8072 22891 8075
rect 22922 8072 22928 8084
rect 22879 8044 22928 8072
rect 22879 8041 22891 8044
rect 22833 8035 22891 8041
rect 22922 8032 22928 8044
rect 22980 8032 22986 8084
rect 23106 8032 23112 8084
rect 23164 8072 23170 8084
rect 23566 8072 23572 8084
rect 23164 8044 23572 8072
rect 23164 8032 23170 8044
rect 23566 8032 23572 8044
rect 23624 8032 23630 8084
rect 26142 8032 26148 8084
rect 26200 8072 26206 8084
rect 26237 8075 26295 8081
rect 26237 8072 26249 8075
rect 26200 8044 26249 8072
rect 26200 8032 26206 8044
rect 26237 8041 26249 8044
rect 26283 8041 26295 8075
rect 26237 8035 26295 8041
rect 29733 8075 29791 8081
rect 29733 8041 29745 8075
rect 29779 8072 29791 8075
rect 29822 8072 29828 8084
rect 29779 8044 29828 8072
rect 29779 8041 29791 8044
rect 29733 8035 29791 8041
rect 29822 8032 29828 8044
rect 29880 8032 29886 8084
rect 20714 8004 20720 8016
rect 20640 7976 20720 8004
rect 20714 7964 20720 7976
rect 20772 7964 20778 8016
rect 11440 7908 12434 7936
rect 4062 7868 4068 7880
rect 4023 7840 4068 7868
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 6546 7828 6552 7880
rect 6604 7828 6610 7880
rect 11440 7877 11468 7908
rect 14274 7896 14280 7948
rect 14332 7936 14338 7948
rect 14461 7939 14519 7945
rect 14461 7936 14473 7939
rect 14332 7908 14473 7936
rect 14332 7896 14338 7908
rect 14461 7905 14473 7908
rect 14507 7905 14519 7939
rect 16500 7936 16528 7964
rect 31386 7936 31392 7948
rect 16500 7908 16804 7936
rect 14461 7899 14519 7905
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7868 11667 7871
rect 14728 7871 14786 7877
rect 11655 7840 11836 7868
rect 11655 7837 11667 7840
rect 11609 7831 11667 7837
rect 4249 7803 4307 7809
rect 4249 7769 4261 7803
rect 4295 7800 4307 7803
rect 4614 7800 4620 7812
rect 4295 7772 4620 7800
rect 4295 7769 4307 7772
rect 4249 7763 4307 7769
rect 4614 7760 4620 7772
rect 4672 7760 4678 7812
rect 5350 7760 5356 7812
rect 5408 7800 5414 7812
rect 5445 7803 5503 7809
rect 5445 7800 5457 7803
rect 5408 7772 5457 7800
rect 5408 7760 5414 7772
rect 5445 7769 5457 7772
rect 5491 7769 5503 7803
rect 11701 7803 11759 7809
rect 11701 7800 11713 7803
rect 10626 7772 11713 7800
rect 5445 7763 5503 7769
rect 11701 7769 11713 7772
rect 11747 7769 11759 7803
rect 11701 7763 11759 7769
rect 6730 7692 6736 7744
rect 6788 7732 6794 7744
rect 11808 7732 11836 7840
rect 14728 7837 14740 7871
rect 14774 7868 14786 7871
rect 15194 7868 15200 7880
rect 14774 7840 15200 7868
rect 14774 7837 14786 7840
rect 14728 7831 14786 7837
rect 15194 7828 15200 7840
rect 15252 7828 15258 7880
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 16485 7871 16543 7877
rect 16485 7868 16497 7871
rect 15528 7840 16497 7868
rect 15528 7828 15534 7840
rect 16485 7837 16497 7840
rect 16531 7837 16543 7871
rect 16666 7868 16672 7880
rect 16627 7840 16672 7868
rect 16485 7831 16543 7837
rect 16500 7800 16528 7831
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 16776 7877 16804 7908
rect 29932 7908 31392 7936
rect 16761 7871 16819 7877
rect 16761 7837 16773 7871
rect 16807 7837 16819 7871
rect 16761 7831 16819 7837
rect 18601 7871 18659 7877
rect 18601 7837 18613 7871
rect 18647 7837 18659 7871
rect 18601 7831 18659 7837
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 19242 7868 19248 7880
rect 18923 7840 19248 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 18616 7800 18644 7831
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 19426 7868 19432 7880
rect 19387 7840 19432 7868
rect 19426 7828 19432 7840
rect 19484 7828 19490 7880
rect 20622 7828 20628 7880
rect 20680 7868 20686 7880
rect 23017 7871 23075 7877
rect 23017 7868 23029 7871
rect 20680 7840 23029 7868
rect 20680 7828 20686 7840
rect 23017 7837 23029 7840
rect 23063 7837 23075 7871
rect 23017 7831 23075 7837
rect 23293 7871 23351 7877
rect 23293 7837 23305 7871
rect 23339 7837 23351 7871
rect 23293 7831 23351 7837
rect 16500 7772 18644 7800
rect 16298 7732 16304 7744
rect 6788 7704 11836 7732
rect 16259 7704 16304 7732
rect 6788 7692 6794 7704
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 18414 7732 18420 7744
rect 18375 7704 18420 7732
rect 18414 7692 18420 7704
rect 18472 7692 18478 7744
rect 18785 7735 18843 7741
rect 18785 7701 18797 7735
rect 18831 7732 18843 7735
rect 18874 7732 18880 7744
rect 18831 7704 18880 7732
rect 18831 7701 18843 7704
rect 18785 7695 18843 7701
rect 18874 7692 18880 7704
rect 18932 7692 18938 7744
rect 19260 7732 19288 7828
rect 19696 7803 19754 7809
rect 19696 7769 19708 7803
rect 19742 7800 19754 7803
rect 20438 7800 20444 7812
rect 19742 7772 20444 7800
rect 19742 7769 19754 7772
rect 19696 7763 19754 7769
rect 20438 7760 20444 7772
rect 20496 7760 20502 7812
rect 20530 7760 20536 7812
rect 20588 7800 20594 7812
rect 23198 7800 23204 7812
rect 20588 7772 23204 7800
rect 20588 7760 20594 7772
rect 23198 7760 23204 7772
rect 23256 7760 23262 7812
rect 20898 7732 20904 7744
rect 19260 7704 20904 7732
rect 20898 7692 20904 7704
rect 20956 7692 20962 7744
rect 23308 7732 23336 7831
rect 24670 7828 24676 7880
rect 24728 7868 24734 7880
rect 24857 7871 24915 7877
rect 24857 7868 24869 7871
rect 24728 7840 24869 7868
rect 24728 7828 24734 7840
rect 24857 7837 24869 7840
rect 24903 7837 24915 7871
rect 24857 7831 24915 7837
rect 27430 7828 27436 7880
rect 27488 7868 27494 7880
rect 29932 7877 29960 7908
rect 31386 7896 31392 7908
rect 31444 7896 31450 7948
rect 29917 7871 29975 7877
rect 29917 7868 29929 7871
rect 27488 7840 29929 7868
rect 27488 7828 27494 7840
rect 29917 7837 29929 7840
rect 29963 7837 29975 7871
rect 30190 7868 30196 7880
rect 30151 7840 30196 7868
rect 29917 7831 29975 7837
rect 30190 7828 30196 7840
rect 30248 7828 30254 7880
rect 25124 7803 25182 7809
rect 25124 7769 25136 7803
rect 25170 7800 25182 7803
rect 25590 7800 25596 7812
rect 25170 7772 25596 7800
rect 25170 7769 25182 7772
rect 25124 7763 25182 7769
rect 25590 7760 25596 7772
rect 25648 7760 25654 7812
rect 30101 7803 30159 7809
rect 30101 7769 30113 7803
rect 30147 7800 30159 7803
rect 31110 7800 31116 7812
rect 30147 7772 31116 7800
rect 30147 7769 30159 7772
rect 30101 7763 30159 7769
rect 31110 7760 31116 7772
rect 31168 7760 31174 7812
rect 25314 7732 25320 7744
rect 23308 7704 25320 7732
rect 25314 7692 25320 7704
rect 25372 7692 25378 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 7006 7528 7012 7540
rect 6967 7500 7012 7528
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 10410 7528 10416 7540
rect 9232 7500 10416 7528
rect 6914 7460 6920 7472
rect 6875 7432 6920 7460
rect 6914 7420 6920 7432
rect 6972 7420 6978 7472
rect 7193 7327 7251 7333
rect 7193 7293 7205 7327
rect 7239 7324 7251 7327
rect 9232 7324 9260 7500
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 15286 7528 15292 7540
rect 12176 7500 15292 7528
rect 9582 7401 9588 7404
rect 9565 7395 9588 7401
rect 9565 7361 9577 7395
rect 9565 7355 9588 7361
rect 9582 7352 9588 7355
rect 9640 7352 9646 7404
rect 12176 7401 12204 7500
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 15746 7528 15752 7540
rect 15659 7500 15752 7528
rect 15746 7488 15752 7500
rect 15804 7528 15810 7540
rect 18046 7528 18052 7540
rect 15804 7500 18052 7528
rect 15804 7488 15810 7500
rect 18046 7488 18052 7500
rect 18104 7488 18110 7540
rect 19334 7488 19340 7540
rect 19392 7528 19398 7540
rect 19521 7531 19579 7537
rect 19521 7528 19533 7531
rect 19392 7500 19533 7528
rect 19392 7488 19398 7500
rect 19521 7497 19533 7500
rect 19567 7497 19579 7531
rect 20438 7528 20444 7540
rect 20399 7500 20444 7528
rect 19521 7491 19579 7497
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 20806 7528 20812 7540
rect 20767 7500 20812 7528
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 24578 7488 24584 7540
rect 24636 7528 24642 7540
rect 24673 7531 24731 7537
rect 24673 7528 24685 7531
rect 24636 7500 24685 7528
rect 24636 7488 24642 7500
rect 24673 7497 24685 7500
rect 24719 7497 24731 7531
rect 25590 7528 25596 7540
rect 25551 7500 25596 7528
rect 24673 7491 24731 7497
rect 25590 7488 25596 7500
rect 25648 7488 25654 7540
rect 25961 7531 26019 7537
rect 25961 7497 25973 7531
rect 26007 7528 26019 7531
rect 26142 7528 26148 7540
rect 26007 7500 26148 7528
rect 26007 7497 26019 7500
rect 25961 7491 26019 7497
rect 26142 7488 26148 7500
rect 26200 7488 26206 7540
rect 29730 7488 29736 7540
rect 29788 7528 29794 7540
rect 29917 7531 29975 7537
rect 29917 7528 29929 7531
rect 29788 7500 29929 7528
rect 29788 7488 29794 7500
rect 29917 7497 29929 7500
rect 29963 7497 29975 7531
rect 29917 7491 29975 7497
rect 14642 7469 14648 7472
rect 14636 7460 14648 7469
rect 14603 7432 14648 7460
rect 14636 7423 14648 7432
rect 14642 7420 14648 7423
rect 14700 7420 14706 7472
rect 18233 7463 18291 7469
rect 18233 7429 18245 7463
rect 18279 7460 18291 7463
rect 20070 7460 20076 7472
rect 18279 7432 20076 7460
rect 18279 7429 18291 7432
rect 18233 7423 18291 7429
rect 19352 7404 19380 7432
rect 20070 7420 20076 7432
rect 20128 7420 20134 7472
rect 23382 7460 23388 7472
rect 23343 7432 23388 7460
rect 23382 7420 23388 7432
rect 23440 7420 23446 7472
rect 25314 7420 25320 7472
rect 25372 7460 25378 7472
rect 25682 7460 25688 7472
rect 25372 7432 25688 7460
rect 25372 7420 25378 7432
rect 25682 7420 25688 7432
rect 25740 7460 25746 7472
rect 28629 7463 28687 7469
rect 25740 7432 26096 7460
rect 25740 7420 25746 7432
rect 12161 7395 12219 7401
rect 12161 7361 12173 7395
rect 12207 7361 12219 7395
rect 12161 7355 12219 7361
rect 12345 7395 12403 7401
rect 12345 7361 12357 7395
rect 12391 7392 12403 7395
rect 12618 7392 12624 7404
rect 12391 7364 12624 7392
rect 12391 7361 12403 7364
rect 12345 7355 12403 7361
rect 12618 7352 12624 7364
rect 12676 7352 12682 7404
rect 14369 7395 14427 7401
rect 14369 7361 14381 7395
rect 14415 7392 14427 7395
rect 14458 7392 14464 7404
rect 14415 7364 14464 7392
rect 14415 7361 14427 7364
rect 14369 7355 14427 7361
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 19334 7352 19340 7404
rect 19392 7352 19398 7404
rect 20622 7392 20628 7404
rect 20583 7364 20628 7392
rect 20622 7352 20628 7364
rect 20680 7352 20686 7404
rect 20898 7392 20904 7404
rect 20859 7364 20904 7392
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 26068 7401 26096 7432
rect 28629 7429 28641 7463
rect 28675 7460 28687 7463
rect 28810 7460 28816 7472
rect 28675 7432 28816 7460
rect 28675 7429 28687 7432
rect 28629 7423 28687 7429
rect 28810 7420 28816 7432
rect 28868 7420 28874 7472
rect 25777 7395 25835 7401
rect 25777 7361 25789 7395
rect 25823 7361 25835 7395
rect 25777 7355 25835 7361
rect 26053 7395 26111 7401
rect 26053 7361 26065 7395
rect 26099 7361 26111 7395
rect 26053 7355 26111 7361
rect 7239 7296 9260 7324
rect 9309 7327 9367 7333
rect 7239 7293 7251 7296
rect 7193 7287 7251 7293
rect 9309 7293 9321 7327
rect 9355 7293 9367 7327
rect 25792 7324 25820 7355
rect 30742 7324 30748 7336
rect 25792 7296 30748 7324
rect 9309 7287 9367 7293
rect 5442 7216 5448 7268
rect 5500 7256 5506 7268
rect 8294 7256 8300 7268
rect 5500 7228 8300 7256
rect 5500 7216 5506 7228
rect 8294 7216 8300 7228
rect 8352 7256 8358 7268
rect 9324 7256 9352 7287
rect 30742 7284 30748 7296
rect 30800 7284 30806 7336
rect 8352 7228 9352 7256
rect 8352 7216 8358 7228
rect 6546 7188 6552 7200
rect 6507 7160 6552 7188
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 10686 7188 10692 7200
rect 10647 7160 10692 7188
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 12158 7188 12164 7200
rect 12119 7160 12164 7188
rect 12158 7148 12164 7160
rect 12216 7148 12222 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 10410 6876 10416 6928
rect 10468 6916 10474 6928
rect 10468 6888 11100 6916
rect 10468 6876 10474 6888
rect 6086 6808 6092 6860
rect 6144 6848 6150 6860
rect 6917 6851 6975 6857
rect 6917 6848 6929 6851
rect 6144 6820 6929 6848
rect 6144 6808 6150 6820
rect 6917 6817 6929 6820
rect 6963 6817 6975 6851
rect 6917 6811 6975 6817
rect 7006 6808 7012 6860
rect 7064 6848 7070 6860
rect 7064 6820 7109 6848
rect 7064 6808 7070 6820
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 11072 6857 11100 6888
rect 10965 6851 11023 6857
rect 10965 6848 10977 6851
rect 10744 6820 10977 6848
rect 10744 6808 10750 6820
rect 10965 6817 10977 6820
rect 11011 6817 11023 6851
rect 10965 6811 11023 6817
rect 11057 6851 11115 6857
rect 11057 6817 11069 6851
rect 11103 6817 11115 6851
rect 11057 6811 11115 6817
rect 6546 6740 6552 6792
rect 6604 6780 6610 6792
rect 6825 6783 6883 6789
rect 6825 6780 6837 6783
rect 6604 6752 6837 6780
rect 6604 6740 6610 6752
rect 6825 6749 6837 6752
rect 6871 6749 6883 6783
rect 10870 6780 10876 6792
rect 10831 6752 10876 6780
rect 6825 6743 6883 6749
rect 10870 6740 10876 6752
rect 10928 6740 10934 6792
rect 14458 6780 14464 6792
rect 14419 6752 14464 6780
rect 14458 6740 14464 6752
rect 14516 6740 14522 6792
rect 14728 6783 14786 6789
rect 14728 6749 14740 6783
rect 14774 6780 14786 6783
rect 16298 6780 16304 6792
rect 14774 6752 16304 6780
rect 14774 6749 14786 6752
rect 14728 6743 14786 6749
rect 16298 6740 16304 6752
rect 16356 6740 16362 6792
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6780 24639 6783
rect 24670 6780 24676 6792
rect 24627 6752 24676 6780
rect 24627 6749 24639 6752
rect 24581 6743 24639 6749
rect 24670 6740 24676 6752
rect 24728 6740 24734 6792
rect 24848 6715 24906 6721
rect 24848 6681 24860 6715
rect 24894 6712 24906 6715
rect 25314 6712 25320 6724
rect 24894 6684 25320 6712
rect 24894 6681 24906 6684
rect 24848 6675 24906 6681
rect 25314 6672 25320 6684
rect 25372 6672 25378 6724
rect 6457 6647 6515 6653
rect 6457 6613 6469 6647
rect 6503 6644 6515 6647
rect 6638 6644 6644 6656
rect 6503 6616 6644 6644
rect 6503 6613 6515 6616
rect 6457 6607 6515 6613
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 10502 6644 10508 6656
rect 10463 6616 10508 6644
rect 10502 6604 10508 6616
rect 10560 6604 10566 6656
rect 15841 6647 15899 6653
rect 15841 6613 15853 6647
rect 15887 6644 15899 6647
rect 16666 6644 16672 6656
rect 15887 6616 16672 6644
rect 15887 6613 15899 6616
rect 15841 6607 15899 6613
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 25958 6644 25964 6656
rect 25919 6616 25964 6644
rect 25958 6604 25964 6616
rect 26016 6604 26022 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 12158 6440 12164 6452
rect 12119 6412 12164 6440
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 18874 6400 18880 6452
rect 18932 6440 18938 6452
rect 19889 6443 19947 6449
rect 19889 6440 19901 6443
rect 18932 6412 19901 6440
rect 18932 6400 18938 6412
rect 19889 6409 19901 6412
rect 19935 6409 19947 6443
rect 25314 6440 25320 6452
rect 25275 6412 25320 6440
rect 19889 6403 19947 6409
rect 25314 6400 25320 6412
rect 25372 6400 25378 6452
rect 25685 6443 25743 6449
rect 25685 6409 25697 6443
rect 25731 6440 25743 6443
rect 25958 6440 25964 6452
rect 25731 6412 25964 6440
rect 25731 6409 25743 6412
rect 25685 6403 25743 6409
rect 25958 6400 25964 6412
rect 26016 6400 26022 6452
rect 10502 6332 10508 6384
rect 10560 6372 10566 6384
rect 12069 6375 12127 6381
rect 12069 6372 12081 6375
rect 10560 6344 12081 6372
rect 10560 6332 10566 6344
rect 12069 6341 12081 6344
rect 12115 6341 12127 6375
rect 12069 6335 12127 6341
rect 18414 6332 18420 6384
rect 18472 6372 18478 6384
rect 18754 6375 18812 6381
rect 18754 6372 18766 6375
rect 18472 6344 18766 6372
rect 18472 6332 18478 6344
rect 18754 6341 18766 6344
rect 18800 6341 18812 6375
rect 27430 6372 27436 6384
rect 18754 6335 18812 6341
rect 25516 6344 27436 6372
rect 25516 6313 25544 6344
rect 27430 6332 27436 6344
rect 27488 6332 27494 6384
rect 25501 6307 25559 6313
rect 25501 6273 25513 6307
rect 25547 6273 25559 6307
rect 25501 6267 25559 6273
rect 25682 6264 25688 6316
rect 25740 6304 25746 6316
rect 25777 6307 25835 6313
rect 25777 6304 25789 6307
rect 25740 6276 25789 6304
rect 25740 6264 25746 6276
rect 25777 6273 25789 6276
rect 25823 6273 25835 6307
rect 25777 6267 25835 6273
rect 12250 6236 12256 6248
rect 12211 6208 12256 6236
rect 12250 6196 12256 6208
rect 12308 6196 12314 6248
rect 18509 6239 18567 6245
rect 18509 6205 18521 6239
rect 18555 6205 18567 6239
rect 18509 6199 18567 6205
rect 11698 6100 11704 6112
rect 11659 6072 11704 6100
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 18524 6100 18552 6199
rect 19426 6100 19432 6112
rect 18524 6072 19432 6100
rect 19426 6060 19432 6072
rect 19484 6060 19490 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 6733 5899 6791 5905
rect 6733 5865 6745 5899
rect 6779 5896 6791 5899
rect 7006 5896 7012 5908
rect 6779 5868 7012 5896
rect 6779 5865 6791 5868
rect 6733 5859 6791 5865
rect 7006 5856 7012 5868
rect 7064 5856 7070 5908
rect 11698 5856 11704 5908
rect 11756 5896 11762 5908
rect 21910 5896 21916 5908
rect 11756 5868 21916 5896
rect 11756 5856 11762 5868
rect 21910 5856 21916 5868
rect 21968 5856 21974 5908
rect 4614 5760 4620 5772
rect 4575 5732 4620 5760
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 4985 5763 5043 5769
rect 4985 5729 4997 5763
rect 5031 5760 5043 5763
rect 5031 5732 6960 5760
rect 5031 5729 5043 5732
rect 4985 5723 5043 5729
rect 5718 5584 5724 5636
rect 5776 5584 5782 5636
rect 6932 5556 6960 5732
rect 7024 5692 7052 5856
rect 27522 5720 27528 5772
rect 27580 5760 27586 5772
rect 27801 5763 27859 5769
rect 27801 5760 27813 5763
rect 27580 5732 27813 5760
rect 27580 5720 27586 5732
rect 27801 5729 27813 5732
rect 27847 5729 27859 5763
rect 27801 5723 27859 5729
rect 10137 5695 10195 5701
rect 10137 5692 10149 5695
rect 7024 5664 10149 5692
rect 10137 5661 10149 5664
rect 10183 5692 10195 5695
rect 10318 5692 10324 5704
rect 10183 5664 10324 5692
rect 10183 5661 10195 5664
rect 10137 5655 10195 5661
rect 10318 5652 10324 5664
rect 10376 5692 10382 5704
rect 12250 5692 12256 5704
rect 10376 5664 12256 5692
rect 10376 5652 10382 5664
rect 12250 5652 12256 5664
rect 12308 5652 12314 5704
rect 28074 5633 28080 5636
rect 28068 5587 28080 5633
rect 28132 5624 28138 5636
rect 28132 5596 28168 5624
rect 28074 5584 28080 5587
rect 28132 5584 28138 5596
rect 9766 5556 9772 5568
rect 6932 5528 9772 5556
rect 9766 5516 9772 5528
rect 9824 5556 9830 5568
rect 10229 5559 10287 5565
rect 10229 5556 10241 5559
rect 9824 5528 10241 5556
rect 9824 5516 9830 5528
rect 10229 5525 10241 5528
rect 10275 5525 10287 5559
rect 10229 5519 10287 5525
rect 28626 5516 28632 5568
rect 28684 5556 28690 5568
rect 29181 5559 29239 5565
rect 29181 5556 29193 5559
rect 28684 5528 29193 5556
rect 28684 5516 28690 5528
rect 29181 5525 29193 5528
rect 29227 5525 29239 5559
rect 29181 5519 29239 5525
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 10134 5352 10140 5364
rect 10095 5324 10140 5352
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 14458 5352 14464 5364
rect 14419 5324 14464 5352
rect 14458 5312 14464 5324
rect 14516 5312 14522 5364
rect 19426 5312 19432 5364
rect 19484 5352 19490 5364
rect 19521 5355 19579 5361
rect 19521 5352 19533 5355
rect 19484 5324 19533 5352
rect 19484 5312 19490 5324
rect 19521 5321 19533 5324
rect 19567 5321 19579 5355
rect 24670 5352 24676 5364
rect 24631 5324 24676 5352
rect 19521 5315 19579 5321
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 29914 5352 29920 5364
rect 29875 5324 29920 5352
rect 29914 5312 29920 5324
rect 29972 5312 29978 5364
rect 5534 5284 5540 5296
rect 5460 5256 5540 5284
rect 5460 5225 5488 5256
rect 5534 5244 5540 5256
rect 5592 5244 5598 5296
rect 5718 5284 5724 5296
rect 5679 5256 5724 5284
rect 5718 5244 5724 5256
rect 5776 5244 5782 5296
rect 12986 5284 12992 5296
rect 12947 5256 12992 5284
rect 12986 5244 12992 5256
rect 13044 5244 13050 5296
rect 18233 5287 18291 5293
rect 18233 5253 18245 5287
rect 18279 5284 18291 5287
rect 19334 5284 19340 5296
rect 18279 5256 19340 5284
rect 18279 5253 18291 5256
rect 18233 5247 18291 5253
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 23382 5284 23388 5296
rect 23343 5256 23388 5284
rect 23382 5244 23388 5256
rect 23440 5244 23446 5296
rect 28629 5287 28687 5293
rect 28629 5253 28641 5287
rect 28675 5284 28687 5287
rect 28810 5284 28816 5296
rect 28675 5256 28816 5284
rect 28675 5253 28687 5256
rect 28629 5247 28687 5253
rect 28810 5244 28816 5256
rect 28868 5244 28874 5296
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5185 5503 5219
rect 5626 5216 5632 5228
rect 5587 5188 5632 5216
rect 5445 5179 5503 5185
rect 5626 5176 5632 5188
rect 5684 5176 5690 5228
rect 9950 5216 9956 5228
rect 9911 5188 9956 5216
rect 9950 5176 9956 5188
rect 10008 5176 10014 5228
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5185 10195 5219
rect 10137 5179 10195 5185
rect 8202 5108 8208 5160
rect 8260 5148 8266 5160
rect 10152 5148 10180 5179
rect 17862 5176 17868 5228
rect 17920 5216 17926 5228
rect 22097 5219 22155 5225
rect 22097 5216 22109 5219
rect 17920 5188 22109 5216
rect 17920 5176 17926 5188
rect 22097 5185 22109 5188
rect 22143 5216 22155 5219
rect 22186 5216 22192 5228
rect 22143 5188 22192 5216
rect 22143 5185 22155 5188
rect 22097 5179 22155 5185
rect 22186 5176 22192 5188
rect 22244 5176 22250 5228
rect 8260 5120 10180 5148
rect 8260 5108 8266 5120
rect 22094 4972 22100 5024
rect 22152 5012 22158 5024
rect 22189 5015 22247 5021
rect 22189 5012 22201 5015
rect 22152 4984 22201 5012
rect 22152 4972 22158 4984
rect 22189 4981 22201 4984
rect 22235 4981 22247 5015
rect 22189 4975 22247 4981
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 10410 4768 10416 4820
rect 10468 4808 10474 4820
rect 11149 4811 11207 4817
rect 11149 4808 11161 4811
rect 10468 4780 11161 4808
rect 10468 4768 10474 4780
rect 11149 4777 11161 4780
rect 11195 4777 11207 4811
rect 11149 4771 11207 4777
rect 12710 4768 12716 4820
rect 12768 4808 12774 4820
rect 12768 4780 14228 4808
rect 12768 4768 12774 4780
rect 7837 4743 7895 4749
rect 7837 4709 7849 4743
rect 7883 4740 7895 4743
rect 9766 4740 9772 4752
rect 7883 4712 9628 4740
rect 7883 4709 7895 4712
rect 7837 4703 7895 4709
rect 5626 4632 5632 4684
rect 5684 4672 5690 4684
rect 9600 4681 9628 4712
rect 9692 4712 9772 4740
rect 9692 4681 9720 4712
rect 9766 4700 9772 4712
rect 9824 4700 9830 4752
rect 8481 4675 8539 4681
rect 5684 4644 6592 4672
rect 5684 4632 5690 4644
rect 6564 4616 6592 4644
rect 8481 4641 8493 4675
rect 8527 4641 8539 4675
rect 8481 4635 8539 4641
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4641 9643 4675
rect 9585 4635 9643 4641
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4641 9735 4675
rect 10428 4672 10456 4768
rect 10505 4743 10563 4749
rect 10505 4709 10517 4743
rect 10551 4740 10563 4743
rect 10551 4712 13492 4740
rect 10551 4709 10563 4712
rect 10505 4703 10563 4709
rect 10597 4675 10655 4681
rect 10597 4672 10609 4675
rect 9677 4635 9735 4641
rect 9784 4644 10609 4672
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 6362 4604 6368 4616
rect 5592 4576 6368 4604
rect 5592 4564 5598 4576
rect 6362 4564 6368 4576
rect 6420 4564 6426 4616
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 8202 4604 8208 4616
rect 6604 4576 6697 4604
rect 8163 4576 8208 4604
rect 6604 4564 6610 4576
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8496 4604 8524 4635
rect 9784 4604 9812 4644
rect 10597 4641 10609 4644
rect 10643 4641 10655 4675
rect 10597 4635 10655 4641
rect 10318 4604 10324 4616
rect 8496 4576 9812 4604
rect 10279 4576 10324 4604
rect 10318 4564 10324 4576
rect 10376 4564 10382 4616
rect 10413 4607 10471 4613
rect 10413 4573 10425 4607
rect 10459 4604 10471 4607
rect 10502 4604 10508 4616
rect 10459 4576 10508 4604
rect 10459 4573 10471 4576
rect 10413 4567 10471 4573
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 10686 4564 10692 4616
rect 10744 4604 10750 4616
rect 11057 4607 11115 4613
rect 11057 4604 11069 4607
rect 10744 4576 11069 4604
rect 10744 4564 10750 4576
rect 11057 4573 11069 4576
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 11333 4607 11391 4613
rect 11333 4573 11345 4607
rect 11379 4573 11391 4607
rect 12710 4604 12716 4616
rect 12671 4576 12716 4604
rect 11333 4567 11391 4573
rect 6733 4539 6791 4545
rect 6733 4505 6745 4539
rect 6779 4536 6791 4539
rect 6914 4536 6920 4548
rect 6779 4508 6920 4536
rect 6779 4505 6791 4508
rect 6733 4499 6791 4505
rect 6914 4496 6920 4508
rect 6972 4496 6978 4548
rect 7926 4496 7932 4548
rect 7984 4536 7990 4548
rect 8297 4539 8355 4545
rect 8297 4536 8309 4539
rect 7984 4508 8309 4536
rect 7984 4496 7990 4508
rect 8297 4505 8309 4508
rect 8343 4505 8355 4539
rect 8297 4499 8355 4505
rect 9493 4539 9551 4545
rect 9493 4505 9505 4539
rect 9539 4536 9551 4539
rect 10226 4536 10232 4548
rect 9539 4508 10232 4536
rect 9539 4505 9551 4508
rect 9493 4499 9551 4505
rect 10226 4496 10232 4508
rect 10284 4496 10290 4548
rect 10336 4536 10364 4564
rect 11348 4536 11376 4567
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 13464 4604 13492 4712
rect 14200 4672 14228 4780
rect 17494 4768 17500 4820
rect 17552 4808 17558 4820
rect 28905 4811 28963 4817
rect 28905 4808 28917 4811
rect 17552 4780 28917 4808
rect 17552 4768 17558 4780
rect 28905 4777 28917 4780
rect 28951 4777 28963 4811
rect 28905 4771 28963 4777
rect 14277 4743 14335 4749
rect 14277 4709 14289 4743
rect 14323 4740 14335 4743
rect 21545 4743 21603 4749
rect 14323 4712 18184 4740
rect 14323 4709 14335 4712
rect 14277 4703 14335 4709
rect 18156 4672 18184 4712
rect 21545 4709 21557 4743
rect 21591 4740 21603 4743
rect 22278 4740 22284 4752
rect 21591 4712 22284 4740
rect 21591 4709 21603 4712
rect 21545 4703 21603 4709
rect 22278 4700 22284 4712
rect 22336 4700 22342 4752
rect 28626 4740 28632 4752
rect 28587 4712 28632 4740
rect 28626 4700 28632 4712
rect 28684 4700 28690 4752
rect 28718 4700 28724 4752
rect 28776 4740 28782 4752
rect 28776 4712 28821 4740
rect 28776 4700 28782 4712
rect 22189 4675 22247 4681
rect 14200 4644 15056 4672
rect 18156 4644 22094 4672
rect 15028 4613 15056 4644
rect 14553 4607 14611 4613
rect 14553 4604 14565 4607
rect 13464 4576 14565 4604
rect 14553 4573 14565 4576
rect 14599 4573 14611 4607
rect 14553 4567 14611 4573
rect 15013 4607 15071 4613
rect 15013 4573 15025 4607
rect 15059 4573 15071 4607
rect 15013 4567 15071 4573
rect 15102 4564 15108 4616
rect 15160 4564 15166 4616
rect 17773 4607 17831 4613
rect 17773 4573 17785 4607
rect 17819 4604 17831 4607
rect 17862 4604 17868 4616
rect 17819 4576 17868 4604
rect 17819 4573 17831 4576
rect 17773 4567 17831 4573
rect 17862 4564 17868 4576
rect 17920 4604 17926 4616
rect 19613 4607 19671 4613
rect 19613 4604 19625 4607
rect 17920 4576 19625 4604
rect 17920 4564 17926 4576
rect 19613 4573 19625 4576
rect 19659 4573 19671 4607
rect 21910 4604 21916 4616
rect 21871 4576 21916 4604
rect 19613 4567 19671 4573
rect 21910 4564 21916 4576
rect 21968 4564 21974 4616
rect 22066 4604 22094 4644
rect 22189 4641 22201 4675
rect 22235 4672 22247 4675
rect 28810 4672 28816 4684
rect 22235 4644 23244 4672
rect 28771 4644 28816 4672
rect 22235 4641 22247 4644
rect 22189 4635 22247 4641
rect 23216 4616 23244 4644
rect 28810 4632 28816 4644
rect 28868 4632 28874 4684
rect 22925 4607 22983 4613
rect 22925 4604 22937 4607
rect 22066 4576 22937 4604
rect 22925 4573 22937 4576
rect 22971 4573 22983 4607
rect 23198 4604 23204 4616
rect 23159 4576 23204 4604
rect 22925 4567 22983 4573
rect 23198 4564 23204 4576
rect 23256 4564 23262 4616
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4604 24639 4607
rect 26421 4607 26479 4613
rect 26421 4604 26433 4607
rect 24627 4576 26433 4604
rect 24627 4573 24639 4576
rect 24581 4567 24639 4573
rect 26421 4573 26433 4576
rect 26467 4604 26479 4607
rect 27154 4604 27160 4616
rect 26467 4576 27160 4604
rect 26467 4573 26479 4576
rect 26421 4567 26479 4573
rect 27154 4564 27160 4576
rect 27212 4604 27218 4616
rect 27522 4604 27528 4616
rect 27212 4576 27528 4604
rect 27212 4564 27218 4576
rect 27522 4564 27528 4576
rect 27580 4564 27586 4616
rect 28261 4607 28319 4613
rect 28261 4604 28273 4607
rect 27816 4576 28273 4604
rect 14277 4539 14335 4545
rect 10336 4508 11376 4536
rect 12406 4508 13492 4536
rect 9122 4468 9128 4480
rect 9083 4440 9128 4468
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 11609 4471 11667 4477
rect 11609 4437 11621 4471
rect 11655 4468 11667 4471
rect 12406 4468 12434 4508
rect 11655 4440 12434 4468
rect 11655 4437 11667 4440
rect 11609 4431 11667 4437
rect 12618 4428 12624 4480
rect 12676 4468 12682 4480
rect 12805 4471 12863 4477
rect 12805 4468 12817 4471
rect 12676 4440 12817 4468
rect 12676 4428 12682 4440
rect 12805 4437 12817 4440
rect 12851 4437 12863 4471
rect 13464 4468 13492 4508
rect 14277 4505 14289 4539
rect 14323 4536 14335 4539
rect 15120 4536 15148 4564
rect 14323 4508 15148 4536
rect 26688 4539 26746 4545
rect 14323 4505 14335 4508
rect 14277 4499 14335 4505
rect 26688 4505 26700 4539
rect 26734 4536 26746 4539
rect 26786 4536 26792 4548
rect 26734 4508 26792 4536
rect 26734 4505 26746 4508
rect 26688 4499 26746 4505
rect 26786 4496 26792 4508
rect 26844 4496 26850 4548
rect 27816 4480 27844 4576
rect 28261 4573 28273 4576
rect 28307 4573 28319 4607
rect 28261 4567 28319 4573
rect 14461 4471 14519 4477
rect 14461 4468 14473 4471
rect 13464 4440 14473 4468
rect 12805 4431 12863 4437
rect 14461 4437 14473 4440
rect 14507 4437 14519 4471
rect 14461 4431 14519 4437
rect 14550 4428 14556 4480
rect 14608 4468 14614 4480
rect 15105 4471 15163 4477
rect 15105 4468 15117 4471
rect 14608 4440 15117 4468
rect 14608 4428 14614 4440
rect 15105 4437 15117 4440
rect 15151 4437 15163 4471
rect 15105 4431 15163 4437
rect 17678 4428 17684 4480
rect 17736 4468 17742 4480
rect 17865 4471 17923 4477
rect 17865 4468 17877 4471
rect 17736 4440 17877 4468
rect 17736 4428 17742 4440
rect 17865 4437 17877 4440
rect 17911 4437 17923 4471
rect 17865 4431 17923 4437
rect 19426 4428 19432 4480
rect 19484 4468 19490 4480
rect 19705 4471 19763 4477
rect 19705 4468 19717 4471
rect 19484 4440 19717 4468
rect 19484 4428 19490 4440
rect 19705 4437 19717 4440
rect 19751 4437 19763 4471
rect 19705 4431 19763 4437
rect 22005 4471 22063 4477
rect 22005 4437 22017 4471
rect 22051 4468 22063 4471
rect 22646 4468 22652 4480
rect 22051 4440 22652 4468
rect 22051 4437 22063 4440
rect 22005 4431 22063 4437
rect 22646 4428 22652 4440
rect 22704 4428 22710 4480
rect 22741 4471 22799 4477
rect 22741 4437 22753 4471
rect 22787 4468 22799 4471
rect 22830 4468 22836 4480
rect 22787 4440 22836 4468
rect 22787 4437 22799 4440
rect 22741 4431 22799 4437
rect 22830 4428 22836 4440
rect 22888 4428 22894 4480
rect 23109 4471 23167 4477
rect 23109 4437 23121 4471
rect 23155 4468 23167 4471
rect 23566 4468 23572 4480
rect 23155 4440 23572 4468
rect 23155 4437 23167 4440
rect 23109 4431 23167 4437
rect 23566 4428 23572 4440
rect 23624 4428 23630 4480
rect 23842 4428 23848 4480
rect 23900 4468 23906 4480
rect 24673 4471 24731 4477
rect 24673 4468 24685 4471
rect 23900 4440 24685 4468
rect 23900 4428 23906 4440
rect 24673 4437 24685 4440
rect 24719 4437 24731 4471
rect 27798 4468 27804 4480
rect 27759 4440 27804 4468
rect 24673 4431 24731 4437
rect 27798 4428 27804 4440
rect 27856 4428 27862 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 7926 4264 7932 4276
rect 7887 4236 7932 4264
rect 7926 4224 7932 4236
rect 7984 4224 7990 4276
rect 9950 4224 9956 4276
rect 10008 4264 10014 4276
rect 10686 4264 10692 4276
rect 10008 4236 10692 4264
rect 10008 4224 10014 4236
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 17862 4224 17868 4276
rect 17920 4224 17926 4276
rect 22646 4224 22652 4276
rect 22704 4264 22710 4276
rect 23014 4264 23020 4276
rect 22704 4236 23020 4264
rect 22704 4224 22710 4236
rect 23014 4224 23020 4236
rect 23072 4264 23078 4276
rect 23385 4267 23443 4273
rect 23385 4264 23397 4267
rect 23072 4236 23397 4264
rect 23072 4224 23078 4236
rect 23385 4233 23397 4236
rect 23431 4233 23443 4267
rect 23385 4227 23443 4233
rect 28537 4267 28595 4273
rect 28537 4233 28549 4267
rect 28583 4264 28595 4267
rect 28810 4264 28816 4276
rect 28583 4236 28816 4264
rect 28583 4233 28595 4236
rect 28537 4227 28595 4233
rect 28810 4224 28816 4236
rect 28868 4224 28874 4276
rect 10226 4156 10232 4208
rect 10284 4156 10290 4208
rect 17880 4196 17908 4224
rect 22278 4205 22284 4208
rect 16868 4168 17908 4196
rect 4706 4088 4712 4140
rect 4764 4128 4770 4140
rect 5902 4128 5908 4140
rect 4764 4100 5908 4128
rect 4764 4088 4770 4100
rect 5902 4088 5908 4100
rect 5960 4128 5966 4140
rect 6805 4131 6863 4137
rect 6805 4128 6817 4131
rect 5960 4100 6817 4128
rect 5960 4088 5966 4100
rect 6805 4097 6817 4100
rect 6851 4097 6863 4131
rect 8938 4128 8944 4140
rect 8899 4100 8944 4128
rect 6805 4091 6863 4097
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 12618 4128 12624 4140
rect 12579 4100 12624 4128
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 12888 4131 12946 4137
rect 12888 4097 12900 4131
rect 12934 4128 12946 4131
rect 14090 4128 14096 4140
rect 12934 4100 14096 4128
rect 12934 4097 12946 4100
rect 12888 4091 12946 4097
rect 14090 4088 14096 4100
rect 14148 4088 14154 4140
rect 14461 4131 14519 4137
rect 14461 4097 14473 4131
rect 14507 4128 14519 4131
rect 14550 4128 14556 4140
rect 14507 4100 14556 4128
rect 14507 4097 14519 4100
rect 14461 4091 14519 4097
rect 14550 4088 14556 4100
rect 14608 4088 14614 4140
rect 14734 4137 14740 4140
rect 14728 4091 14740 4137
rect 14792 4128 14798 4140
rect 16868 4137 16896 4168
rect 22272 4159 22284 4205
rect 22336 4196 22342 4208
rect 22336 4168 22372 4196
rect 27172 4168 27568 4196
rect 22278 4156 22284 4159
rect 22336 4156 22342 4168
rect 27172 4140 27200 4168
rect 16853 4131 16911 4137
rect 14792 4100 14828 4128
rect 14734 4088 14740 4091
rect 14792 4088 14798 4100
rect 16853 4097 16865 4131
rect 16899 4097 16911 4131
rect 17678 4128 17684 4140
rect 17639 4100 17684 4128
rect 16853 4091 16911 4097
rect 17678 4088 17684 4100
rect 17736 4088 17742 4140
rect 17948 4131 18006 4137
rect 17948 4097 17960 4131
rect 17994 4128 18006 4131
rect 18414 4128 18420 4140
rect 17994 4100 18420 4128
rect 17994 4097 18006 4100
rect 17948 4091 18006 4097
rect 18414 4088 18420 4100
rect 18472 4088 18478 4140
rect 19426 4088 19432 4140
rect 19484 4128 19490 4140
rect 19794 4137 19800 4140
rect 19521 4131 19579 4137
rect 19521 4128 19533 4131
rect 19484 4100 19533 4128
rect 19484 4088 19490 4100
rect 19521 4097 19533 4100
rect 19567 4097 19579 4131
rect 19521 4091 19579 4097
rect 19788 4091 19800 4137
rect 19852 4128 19858 4140
rect 22005 4131 22063 4137
rect 19852 4100 19888 4128
rect 19794 4088 19800 4091
rect 19852 4088 19858 4100
rect 22005 4097 22017 4131
rect 22051 4128 22063 4131
rect 22094 4128 22100 4140
rect 22051 4100 22100 4128
rect 22051 4097 22063 4100
rect 22005 4091 22063 4097
rect 22094 4088 22100 4100
rect 22152 4088 22158 4140
rect 23842 4128 23848 4140
rect 23803 4100 23848 4128
rect 23842 4088 23848 4100
rect 23900 4088 23906 4140
rect 24112 4131 24170 4137
rect 24112 4097 24124 4131
rect 24158 4128 24170 4131
rect 24578 4128 24584 4140
rect 24158 4100 24584 4128
rect 24158 4097 24170 4100
rect 24112 4091 24170 4097
rect 24578 4088 24584 4100
rect 24636 4088 24642 4140
rect 27154 4128 27160 4140
rect 27115 4100 27160 4128
rect 27154 4088 27160 4100
rect 27212 4088 27218 4140
rect 27413 4131 27471 4137
rect 27413 4128 27425 4131
rect 27264 4100 27425 4128
rect 6549 4063 6607 4069
rect 6549 4029 6561 4063
rect 6595 4029 6607 4063
rect 9214 4060 9220 4072
rect 9175 4032 9220 4060
rect 6549 4023 6607 4029
rect 6564 3924 6592 4023
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 26145 4063 26203 4069
rect 26145 4029 26157 4063
rect 26191 4060 26203 4063
rect 26418 4060 26424 4072
rect 26191 4032 26424 4060
rect 26191 4029 26203 4032
rect 26145 4023 26203 4029
rect 26418 4020 26424 4032
rect 26476 4020 26482 4072
rect 26605 4063 26663 4069
rect 26605 4029 26617 4063
rect 26651 4060 26663 4063
rect 27264 4060 27292 4100
rect 27413 4097 27425 4100
rect 27459 4097 27471 4131
rect 27540 4128 27568 4168
rect 28997 4131 29055 4137
rect 28997 4128 29009 4131
rect 27540 4100 29009 4128
rect 27413 4091 27471 4097
rect 28997 4097 29009 4100
rect 29043 4097 29055 4131
rect 28997 4091 29055 4097
rect 29086 4088 29092 4140
rect 29144 4128 29150 4140
rect 29253 4131 29311 4137
rect 29253 4128 29265 4131
rect 29144 4100 29265 4128
rect 29144 4088 29150 4100
rect 29253 4097 29265 4100
rect 29299 4097 29311 4131
rect 29253 4091 29311 4097
rect 26651 4032 27292 4060
rect 26651 4029 26663 4032
rect 26605 4023 26663 4029
rect 15841 3995 15899 4001
rect 15841 3961 15853 3995
rect 15887 3992 15899 3995
rect 17126 3992 17132 4004
rect 15887 3964 17132 3992
rect 15887 3961 15899 3964
rect 15841 3955 15899 3961
rect 17126 3952 17132 3964
rect 17184 3952 17190 4004
rect 26513 3995 26571 4001
rect 26513 3961 26525 3995
rect 26559 3961 26571 3995
rect 26513 3955 26571 3961
rect 8294 3924 8300 3936
rect 6564 3896 8300 3924
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 14001 3927 14059 3933
rect 14001 3893 14013 3927
rect 14047 3924 14059 3927
rect 14458 3924 14464 3936
rect 14047 3896 14464 3924
rect 14047 3893 14059 3896
rect 14001 3887 14059 3893
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 16574 3884 16580 3936
rect 16632 3924 16638 3936
rect 16945 3927 17003 3933
rect 16945 3924 16957 3927
rect 16632 3896 16957 3924
rect 16632 3884 16638 3896
rect 16945 3893 16957 3896
rect 16991 3893 17003 3927
rect 16945 3887 17003 3893
rect 19061 3927 19119 3933
rect 19061 3893 19073 3927
rect 19107 3924 19119 3927
rect 19334 3924 19340 3936
rect 19107 3896 19340 3924
rect 19107 3893 19119 3896
rect 19061 3887 19119 3893
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 20898 3924 20904 3936
rect 20859 3896 20904 3924
rect 20898 3884 20904 3896
rect 20956 3884 20962 3936
rect 25038 3884 25044 3936
rect 25096 3924 25102 3936
rect 25225 3927 25283 3933
rect 25225 3924 25237 3927
rect 25096 3896 25237 3924
rect 25096 3884 25102 3896
rect 25225 3893 25237 3896
rect 25271 3893 25283 3927
rect 26528 3924 26556 3955
rect 27430 3924 27436 3936
rect 26528 3896 27436 3924
rect 25225 3887 25283 3893
rect 27430 3884 27436 3896
rect 27488 3884 27494 3936
rect 28718 3884 28724 3936
rect 28776 3924 28782 3936
rect 30377 3927 30435 3933
rect 30377 3924 30389 3927
rect 28776 3896 30389 3924
rect 28776 3884 28782 3896
rect 30377 3893 30389 3896
rect 30423 3924 30435 3927
rect 32306 3924 32312 3936
rect 30423 3896 32312 3924
rect 30423 3893 30435 3896
rect 30377 3887 30435 3893
rect 32306 3884 32312 3896
rect 32364 3884 32370 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 6638 3680 6644 3732
rect 6696 3720 6702 3732
rect 7377 3723 7435 3729
rect 6696 3692 7328 3720
rect 6696 3680 6702 3692
rect 7300 3652 7328 3692
rect 7377 3689 7389 3723
rect 7423 3720 7435 3723
rect 8202 3720 8208 3732
rect 7423 3692 8208 3720
rect 7423 3689 7435 3692
rect 7377 3683 7435 3689
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 9508 3692 10456 3720
rect 9508 3652 9536 3692
rect 7300 3624 9536 3652
rect 10428 3652 10456 3692
rect 10502 3680 10508 3732
rect 10560 3720 10566 3732
rect 10873 3723 10931 3729
rect 10873 3720 10885 3723
rect 10560 3692 10885 3720
rect 10560 3680 10566 3692
rect 10873 3689 10885 3692
rect 10919 3689 10931 3723
rect 10873 3683 10931 3689
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 14829 3723 14887 3729
rect 14829 3720 14841 3723
rect 14792 3692 14841 3720
rect 14792 3680 14798 3692
rect 14829 3689 14841 3692
rect 14875 3689 14887 3723
rect 19794 3720 19800 3732
rect 14829 3683 14887 3689
rect 16592 3692 17632 3720
rect 19755 3692 19800 3720
rect 16592 3652 16620 3692
rect 10428 3624 16620 3652
rect 5902 3584 5908 3596
rect 5863 3556 5908 3584
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 9180 3556 9628 3584
rect 9180 3544 9186 3556
rect 5629 3519 5687 3525
rect 5629 3485 5641 3519
rect 5675 3485 5687 3519
rect 5629 3479 5687 3485
rect 5644 3380 5672 3479
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 9493 3519 9551 3525
rect 9493 3516 9505 3519
rect 8352 3488 9505 3516
rect 8352 3476 8358 3488
rect 9493 3485 9505 3488
rect 9539 3485 9551 3519
rect 9600 3516 9628 3556
rect 15102 3544 15108 3596
rect 15160 3584 15166 3596
rect 15381 3587 15439 3593
rect 15381 3584 15393 3587
rect 15160 3556 15393 3584
rect 15160 3544 15166 3556
rect 15381 3553 15393 3556
rect 15427 3553 15439 3587
rect 16574 3584 16580 3596
rect 16535 3556 16580 3584
rect 15381 3547 15439 3553
rect 16574 3544 16580 3556
rect 16632 3544 16638 3596
rect 17604 3516 17632 3692
rect 19794 3680 19800 3692
rect 19852 3680 19858 3732
rect 23198 3720 23204 3732
rect 22066 3692 23204 3720
rect 19058 3544 19064 3596
rect 19116 3584 19122 3596
rect 20441 3587 20499 3593
rect 20441 3584 20453 3587
rect 19116 3556 20453 3584
rect 19116 3544 19122 3556
rect 20441 3553 20453 3556
rect 20487 3584 20499 3587
rect 22066 3584 22094 3692
rect 23198 3680 23204 3692
rect 23256 3680 23262 3732
rect 23566 3680 23572 3732
rect 23624 3720 23630 3732
rect 23750 3720 23756 3732
rect 23624 3692 23756 3720
rect 23624 3680 23630 3692
rect 23750 3680 23756 3692
rect 23808 3720 23814 3732
rect 23937 3723 23995 3729
rect 23937 3720 23949 3723
rect 23808 3692 23949 3720
rect 23808 3680 23814 3692
rect 23937 3689 23949 3692
rect 23983 3689 23995 3723
rect 24578 3720 24584 3732
rect 24539 3692 24584 3720
rect 23937 3683 23995 3689
rect 24578 3680 24584 3692
rect 24636 3680 24642 3732
rect 26786 3720 26792 3732
rect 26747 3692 26792 3720
rect 26786 3680 26792 3692
rect 26844 3680 26850 3732
rect 27430 3680 27436 3732
rect 27488 3720 27494 3732
rect 27709 3723 27767 3729
rect 27709 3720 27721 3723
rect 27488 3692 27721 3720
rect 27488 3680 27494 3692
rect 27709 3689 27721 3692
rect 27755 3720 27767 3723
rect 27798 3720 27804 3732
rect 27755 3692 27804 3720
rect 27755 3689 27767 3692
rect 27709 3683 27767 3689
rect 27798 3680 27804 3692
rect 27856 3680 27862 3732
rect 28626 3680 28632 3732
rect 28684 3720 28690 3732
rect 29086 3720 29092 3732
rect 28684 3692 28948 3720
rect 29047 3692 29092 3720
rect 28684 3680 28690 3692
rect 28920 3664 28948 3692
rect 29086 3680 29092 3692
rect 29144 3680 29150 3732
rect 27617 3655 27675 3661
rect 27617 3652 27629 3655
rect 26620 3624 27629 3652
rect 25038 3584 25044 3596
rect 20487 3556 22094 3584
rect 24999 3556 25044 3584
rect 20487 3553 20499 3556
rect 20441 3547 20499 3553
rect 25038 3544 25044 3556
rect 25096 3544 25102 3596
rect 25225 3587 25283 3593
rect 25225 3553 25237 3587
rect 25271 3584 25283 3587
rect 25271 3556 25728 3584
rect 25271 3553 25283 3556
rect 25225 3547 25283 3553
rect 20165 3519 20223 3525
rect 20165 3516 20177 3519
rect 9600 3488 17264 3516
rect 17604 3488 20177 3516
rect 9493 3479 9551 3485
rect 6914 3408 6920 3460
rect 6972 3408 6978 3460
rect 9214 3408 9220 3460
rect 9272 3448 9278 3460
rect 9738 3451 9796 3457
rect 9738 3448 9750 3451
rect 9272 3420 9750 3448
rect 9272 3408 9278 3420
rect 9738 3417 9750 3420
rect 9784 3417 9796 3451
rect 9738 3411 9796 3417
rect 11054 3408 11060 3460
rect 11112 3448 11118 3460
rect 16850 3457 16856 3460
rect 15197 3451 15255 3457
rect 15197 3448 15209 3451
rect 11112 3420 15209 3448
rect 11112 3408 11118 3420
rect 15197 3417 15209 3420
rect 15243 3417 15255 3451
rect 15197 3411 15255 3417
rect 16844 3411 16856 3457
rect 16908 3448 16914 3460
rect 17236 3448 17264 3488
rect 20165 3485 20177 3488
rect 20211 3485 20223 3519
rect 20165 3479 20223 3485
rect 20257 3519 20315 3525
rect 20257 3485 20269 3519
rect 20303 3516 20315 3519
rect 20898 3516 20904 3528
rect 20303 3488 20904 3516
rect 20303 3485 20315 3488
rect 20257 3479 20315 3485
rect 20898 3476 20904 3488
rect 20956 3476 20962 3528
rect 22554 3516 22560 3528
rect 22515 3488 22560 3516
rect 22554 3476 22560 3488
rect 22612 3476 22618 3528
rect 22830 3525 22836 3528
rect 22824 3516 22836 3525
rect 22791 3488 22836 3516
rect 22824 3479 22836 3488
rect 22830 3476 22836 3479
rect 22888 3476 22894 3528
rect 23198 3476 23204 3528
rect 23256 3516 23262 3528
rect 25240 3516 25268 3547
rect 23256 3488 25268 3516
rect 23256 3476 23262 3488
rect 24949 3451 25007 3457
rect 24949 3448 24961 3451
rect 16908 3420 16944 3448
rect 17236 3420 24961 3448
rect 16850 3408 16856 3411
rect 16908 3408 16914 3420
rect 24949 3417 24961 3420
rect 24995 3448 25007 3451
rect 25593 3451 25651 3457
rect 25593 3448 25605 3451
rect 24995 3420 25605 3448
rect 24995 3417 25007 3420
rect 24949 3411 25007 3417
rect 25593 3417 25605 3420
rect 25639 3417 25651 3451
rect 25593 3411 25651 3417
rect 8938 3380 8944 3392
rect 5644 3352 8944 3380
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 15289 3383 15347 3389
rect 15289 3349 15301 3383
rect 15335 3380 15347 3383
rect 17126 3380 17132 3392
rect 15335 3352 17132 3380
rect 15335 3349 15347 3352
rect 15289 3343 15347 3349
rect 17126 3340 17132 3352
rect 17184 3340 17190 3392
rect 17954 3380 17960 3392
rect 17915 3352 17960 3380
rect 17954 3340 17960 3352
rect 18012 3340 18018 3392
rect 25700 3380 25728 3556
rect 26620 3525 26648 3624
rect 27617 3621 27629 3624
rect 27663 3652 27675 3655
rect 28718 3652 28724 3664
rect 27663 3624 28724 3652
rect 27663 3621 27675 3624
rect 27617 3615 27675 3621
rect 28718 3612 28724 3624
rect 28776 3612 28782 3664
rect 28902 3612 28908 3664
rect 28960 3652 28966 3664
rect 28960 3624 29053 3652
rect 28960 3612 28966 3624
rect 27801 3587 27859 3593
rect 27801 3553 27813 3587
rect 27847 3584 27859 3587
rect 27890 3584 27896 3596
rect 27847 3556 27896 3584
rect 27847 3553 27859 3556
rect 27801 3547 27859 3553
rect 27890 3544 27896 3556
rect 27948 3584 27954 3596
rect 28810 3584 28816 3596
rect 27948 3556 28816 3584
rect 27948 3544 27954 3556
rect 28810 3544 28816 3556
rect 28868 3544 28874 3596
rect 26605 3519 26663 3525
rect 26605 3485 26617 3519
rect 26651 3485 26663 3519
rect 26605 3479 26663 3485
rect 27249 3519 27307 3525
rect 27249 3485 27261 3519
rect 27295 3516 27307 3519
rect 28902 3516 28908 3528
rect 27295 3488 28908 3516
rect 27295 3485 27307 3488
rect 27249 3479 27307 3485
rect 28902 3476 28908 3488
rect 28960 3476 28966 3528
rect 26418 3448 26424 3460
rect 26379 3420 26424 3448
rect 26418 3408 26424 3420
rect 26476 3448 26482 3460
rect 28629 3451 28687 3457
rect 28629 3448 28641 3451
rect 26476 3420 28641 3448
rect 26476 3408 26482 3420
rect 28629 3417 28641 3420
rect 28675 3417 28687 3451
rect 28629 3411 28687 3417
rect 28077 3383 28135 3389
rect 28077 3380 28089 3383
rect 25700 3352 28089 3380
rect 28077 3349 28089 3352
rect 28123 3349 28135 3383
rect 28077 3343 28135 3349
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 1596 3148 2774 3176
rect 1596 3049 1624 3148
rect 2746 3108 2774 3148
rect 10134 3136 10140 3188
rect 10192 3176 10198 3188
rect 12710 3176 12716 3188
rect 10192 3148 12716 3176
rect 10192 3136 10198 3148
rect 12710 3136 12716 3148
rect 12768 3136 12774 3188
rect 14090 3176 14096 3188
rect 14051 3148 14096 3176
rect 14090 3136 14096 3148
rect 14148 3136 14154 3188
rect 14458 3136 14464 3188
rect 14516 3176 14522 3188
rect 14553 3179 14611 3185
rect 14553 3176 14565 3179
rect 14516 3148 14565 3176
rect 14516 3136 14522 3148
rect 14553 3145 14565 3148
rect 14599 3176 14611 3179
rect 15654 3176 15660 3188
rect 14599 3148 15660 3176
rect 14599 3145 14611 3148
rect 14553 3139 14611 3145
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 16850 3176 16856 3188
rect 16811 3148 16856 3176
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 17218 3176 17224 3188
rect 17179 3148 17224 3176
rect 17218 3136 17224 3148
rect 17276 3136 17282 3188
rect 17313 3179 17371 3185
rect 17313 3145 17325 3179
rect 17359 3176 17371 3179
rect 17954 3176 17960 3188
rect 17359 3148 17960 3176
rect 17359 3145 17371 3148
rect 17313 3139 17371 3145
rect 17954 3136 17960 3148
rect 18012 3136 18018 3188
rect 18414 3176 18420 3188
rect 18375 3148 18420 3176
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 22554 3136 22560 3188
rect 22612 3176 22618 3188
rect 22741 3179 22799 3185
rect 22741 3176 22753 3179
rect 22612 3148 22753 3176
rect 22612 3136 22618 3148
rect 22741 3145 22753 3148
rect 22787 3145 22799 3179
rect 22741 3139 22799 3145
rect 27985 3179 28043 3185
rect 27985 3145 27997 3179
rect 28031 3176 28043 3179
rect 28074 3176 28080 3188
rect 28031 3148 28080 3176
rect 28031 3145 28043 3148
rect 27985 3139 28043 3145
rect 28074 3136 28080 3148
rect 28132 3136 28138 3188
rect 8478 3108 8484 3120
rect 2746 3080 8484 3108
rect 8478 3068 8484 3080
rect 8536 3108 8542 3120
rect 8536 3080 12434 3108
rect 8536 3068 8542 3080
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 6362 3000 6368 3052
rect 6420 3040 6426 3052
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 6420 3012 9873 3040
rect 6420 3000 6426 3012
rect 9861 3009 9873 3012
rect 9907 3040 9919 3043
rect 9950 3040 9956 3052
rect 9907 3012 9956 3040
rect 9907 3009 9919 3012
rect 9861 3003 9919 3009
rect 9950 3000 9956 3012
rect 10008 3000 10014 3052
rect 10045 3043 10103 3049
rect 10045 3009 10057 3043
rect 10091 3009 10103 3043
rect 12406 3040 12434 3080
rect 14461 3043 14519 3049
rect 14461 3040 14473 3043
rect 12406 3012 14473 3040
rect 10045 3003 10103 3009
rect 14461 3009 14473 3012
rect 14507 3009 14519 3043
rect 18782 3040 18788 3052
rect 18743 3012 18788 3040
rect 14461 3003 14519 3009
rect 842 2932 848 2984
rect 900 2972 906 2984
rect 1765 2975 1823 2981
rect 1765 2972 1777 2975
rect 900 2944 1777 2972
rect 900 2932 906 2944
rect 1765 2941 1777 2944
rect 1811 2941 1823 2975
rect 1765 2935 1823 2941
rect 6546 2932 6552 2984
rect 6604 2972 6610 2984
rect 10060 2972 10088 3003
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 18877 3043 18935 3049
rect 18877 3009 18889 3043
rect 18923 3040 18935 3043
rect 19334 3040 19340 3052
rect 18923 3012 19340 3040
rect 18923 3009 18935 3012
rect 18877 3003 18935 3009
rect 19334 3000 19340 3012
rect 19392 3040 19398 3052
rect 20070 3040 20076 3052
rect 19392 3012 20076 3040
rect 19392 3000 19398 3012
rect 20070 3000 20076 3012
rect 20128 3000 20134 3052
rect 22186 3000 22192 3052
rect 22244 3040 22250 3052
rect 22649 3043 22707 3049
rect 22649 3040 22661 3043
rect 22244 3012 22661 3040
rect 22244 3000 22250 3012
rect 22649 3009 22661 3012
rect 22695 3009 22707 3043
rect 22649 3003 22707 3009
rect 10226 2972 10232 2984
rect 6604 2944 10088 2972
rect 10187 2944 10232 2972
rect 6604 2932 6610 2944
rect 10226 2932 10232 2944
rect 10284 2932 10290 2984
rect 14737 2975 14795 2981
rect 14737 2941 14749 2975
rect 14783 2972 14795 2975
rect 15102 2972 15108 2984
rect 14783 2944 15108 2972
rect 14783 2941 14795 2944
rect 14737 2935 14795 2941
rect 15102 2932 15108 2944
rect 15160 2972 15166 2984
rect 17497 2975 17555 2981
rect 17497 2972 17509 2975
rect 15160 2944 17509 2972
rect 15160 2932 15166 2944
rect 17497 2941 17509 2944
rect 17543 2972 17555 2975
rect 19058 2972 19064 2984
rect 17543 2944 19064 2972
rect 17543 2941 17555 2944
rect 17497 2935 17555 2941
rect 19058 2932 19064 2944
rect 19116 2932 19122 2984
rect 27525 2975 27583 2981
rect 27525 2941 27537 2975
rect 27571 2941 27583 2975
rect 27525 2935 27583 2941
rect 38105 2975 38163 2981
rect 38105 2941 38117 2975
rect 38151 2972 38163 2975
rect 39114 2972 39120 2984
rect 38151 2944 39120 2972
rect 38151 2941 38163 2944
rect 38105 2935 38163 2941
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 26418 2904 26424 2916
rect 9732 2876 26424 2904
rect 9732 2864 9738 2876
rect 26418 2864 26424 2876
rect 26476 2904 26482 2916
rect 27540 2904 27568 2935
rect 39114 2932 39120 2944
rect 39172 2932 39178 2984
rect 27890 2904 27896 2916
rect 26476 2876 27568 2904
rect 27851 2876 27896 2904
rect 26476 2864 26482 2876
rect 27890 2864 27896 2876
rect 27948 2864 27954 2916
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 6362 2592 6368 2644
rect 6420 2632 6426 2644
rect 18782 2632 18788 2644
rect 6420 2604 18788 2632
rect 6420 2592 6426 2604
rect 18782 2592 18788 2604
rect 18840 2592 18846 2644
rect 11054 2564 11060 2576
rect 2424 2536 11060 2564
rect 2424 2437 2452 2536
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 11146 2524 11152 2576
rect 11204 2524 11210 2576
rect 11164 2496 11192 2524
rect 3988 2468 11192 2496
rect 3988 2437 4016 2468
rect 28902 2456 28908 2508
rect 28960 2496 28966 2508
rect 28960 2468 30696 2496
rect 28960 2456 28966 2468
rect 2409 2431 2467 2437
rect 2409 2397 2421 2431
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 5353 2431 5411 2437
rect 5353 2397 5365 2431
rect 5399 2428 5411 2431
rect 6362 2428 6368 2440
rect 5399 2400 6368 2428
rect 5399 2397 5411 2400
rect 5353 2391 5411 2397
rect 6362 2388 6368 2400
rect 6420 2388 6426 2440
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 7009 2431 7067 2437
rect 7009 2428 7021 2431
rect 6788 2400 7021 2428
rect 6788 2388 6794 2400
rect 7009 2397 7021 2400
rect 7055 2397 7067 2431
rect 7009 2391 7067 2397
rect 8202 2388 8208 2440
rect 8260 2428 8266 2440
rect 8481 2431 8539 2437
rect 8481 2428 8493 2431
rect 8260 2400 8493 2428
rect 8260 2388 8266 2400
rect 8481 2397 8493 2400
rect 8527 2397 8539 2431
rect 8481 2391 8539 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 9732 2400 9965 2428
rect 9732 2388 9738 2400
rect 9953 2397 9965 2400
rect 9999 2397 10011 2431
rect 9953 2391 10011 2397
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11204 2400 11897 2428
rect 11204 2388 11210 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 12618 2388 12624 2440
rect 12676 2428 12682 2440
rect 12897 2431 12955 2437
rect 12897 2428 12909 2431
rect 12676 2400 12909 2428
rect 12676 2388 12682 2400
rect 12897 2397 12909 2400
rect 12943 2397 12955 2431
rect 12897 2391 12955 2397
rect 14090 2388 14096 2440
rect 14148 2428 14154 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 14148 2400 14473 2428
rect 14148 2388 14154 2400
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 15654 2428 15660 2440
rect 15615 2400 15660 2428
rect 14461 2391 14519 2397
rect 15654 2388 15660 2400
rect 15712 2388 15718 2440
rect 17126 2428 17132 2440
rect 17087 2400 17132 2428
rect 17126 2388 17132 2400
rect 17184 2388 17190 2440
rect 17954 2388 17960 2440
rect 18012 2428 18018 2440
rect 18417 2431 18475 2437
rect 18417 2428 18429 2431
rect 18012 2400 18429 2428
rect 18012 2388 18018 2400
rect 18417 2397 18429 2400
rect 18463 2397 18475 2431
rect 20070 2428 20076 2440
rect 20031 2400 20076 2428
rect 18417 2391 18475 2397
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 20898 2388 20904 2440
rect 20956 2428 20962 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 20956 2400 22017 2428
rect 20956 2388 20962 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 23014 2428 23020 2440
rect 22975 2400 23020 2428
rect 22005 2391 22063 2397
rect 23014 2388 23020 2400
rect 23072 2388 23078 2440
rect 23750 2388 23756 2440
rect 23808 2428 23814 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 23808 2400 24593 2428
rect 23808 2388 23814 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 25038 2388 25044 2440
rect 25096 2428 25102 2440
rect 25961 2431 26019 2437
rect 25961 2428 25973 2431
rect 25096 2400 25973 2428
rect 25096 2388 25102 2400
rect 25961 2397 25973 2400
rect 26007 2397 26019 2431
rect 27430 2428 27436 2440
rect 27391 2400 27436 2428
rect 25961 2391 26019 2397
rect 27430 2388 27436 2400
rect 27488 2388 27494 2440
rect 27890 2388 27896 2440
rect 27948 2428 27954 2440
rect 30668 2437 30696 2468
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 27948 2400 29745 2428
rect 27948 2388 27954 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30653 2431 30711 2437
rect 30653 2397 30665 2431
rect 30699 2397 30711 2431
rect 32306 2428 32312 2440
rect 32267 2400 32312 2428
rect 30653 2391 30711 2397
rect 32306 2388 32312 2400
rect 32364 2388 32370 2440
rect 33226 2388 33232 2440
rect 33284 2428 33290 2440
rect 33505 2431 33563 2437
rect 33505 2428 33517 2431
rect 33284 2400 33517 2428
rect 33284 2388 33290 2400
rect 33505 2397 33517 2400
rect 33551 2397 33563 2431
rect 33505 2391 33563 2397
rect 34698 2388 34704 2440
rect 34756 2428 34762 2440
rect 35069 2431 35127 2437
rect 35069 2428 35081 2431
rect 34756 2400 35081 2428
rect 34756 2388 34762 2400
rect 35069 2397 35081 2400
rect 35115 2397 35127 2431
rect 35069 2391 35127 2397
rect 36170 2388 36176 2440
rect 36228 2428 36234 2440
rect 36449 2431 36507 2437
rect 36449 2428 36461 2431
rect 36228 2400 36461 2428
rect 36228 2388 36234 2400
rect 36449 2397 36461 2400
rect 36495 2397 36507 2431
rect 36449 2391 36507 2397
rect 37642 2388 37648 2440
rect 37700 2428 37706 2440
rect 37921 2431 37979 2437
rect 37921 2428 37933 2431
rect 37700 2400 37933 2428
rect 37700 2388 37706 2400
rect 37921 2397 37933 2400
rect 37967 2397 37979 2431
rect 37921 2391 37979 2397
rect 2314 2320 2320 2372
rect 2372 2360 2378 2372
rect 2685 2363 2743 2369
rect 2685 2360 2697 2363
rect 2372 2332 2697 2360
rect 2372 2320 2378 2332
rect 2685 2329 2697 2332
rect 2731 2329 2743 2363
rect 2685 2323 2743 2329
rect 3786 2320 3792 2372
rect 3844 2360 3850 2372
rect 4249 2363 4307 2369
rect 4249 2360 4261 2363
rect 3844 2332 4261 2360
rect 3844 2320 3850 2332
rect 4249 2329 4261 2332
rect 4295 2329 4307 2363
rect 4249 2323 4307 2329
rect 5258 2320 5264 2372
rect 5316 2360 5322 2372
rect 5629 2363 5687 2369
rect 5629 2360 5641 2363
rect 5316 2332 5641 2360
rect 5316 2320 5322 2332
rect 5629 2329 5641 2332
rect 5675 2329 5687 2363
rect 5629 2323 5687 2329
rect 15562 2320 15568 2372
rect 15620 2360 15626 2372
rect 15933 2363 15991 2369
rect 15933 2360 15945 2363
rect 15620 2332 15945 2360
rect 15620 2320 15626 2332
rect 15933 2329 15945 2332
rect 15979 2329 15991 2363
rect 15933 2323 15991 2329
rect 17034 2320 17040 2372
rect 17092 2360 17098 2372
rect 17405 2363 17463 2369
rect 17405 2360 17417 2363
rect 17092 2332 17417 2360
rect 17092 2320 17098 2332
rect 17405 2329 17417 2332
rect 17451 2329 17463 2363
rect 17405 2323 17463 2329
rect 18506 2320 18512 2372
rect 18564 2360 18570 2372
rect 18693 2363 18751 2369
rect 18693 2360 18705 2363
rect 18564 2332 18705 2360
rect 18564 2320 18570 2332
rect 18693 2329 18705 2332
rect 18739 2329 18751 2363
rect 18693 2323 18751 2329
rect 19978 2320 19984 2372
rect 20036 2360 20042 2372
rect 20349 2363 20407 2369
rect 20349 2360 20361 2363
rect 20036 2332 20361 2360
rect 20036 2320 20042 2332
rect 20349 2329 20361 2332
rect 20395 2329 20407 2363
rect 20349 2323 20407 2329
rect 21450 2320 21456 2372
rect 21508 2360 21514 2372
rect 22281 2363 22339 2369
rect 22281 2360 22293 2363
rect 21508 2332 22293 2360
rect 21508 2320 21514 2332
rect 22281 2329 22293 2332
rect 22327 2329 22339 2363
rect 22281 2323 22339 2329
rect 22922 2320 22928 2372
rect 22980 2360 22986 2372
rect 23293 2363 23351 2369
rect 23293 2360 23305 2363
rect 22980 2332 23305 2360
rect 22980 2320 22986 2332
rect 23293 2329 23305 2332
rect 23339 2329 23351 2363
rect 23293 2323 23351 2329
rect 24394 2320 24400 2372
rect 24452 2360 24458 2372
rect 24857 2363 24915 2369
rect 24857 2360 24869 2363
rect 24452 2332 24869 2360
rect 24452 2320 24458 2332
rect 24857 2329 24869 2332
rect 24903 2329 24915 2363
rect 24857 2323 24915 2329
rect 25866 2320 25872 2372
rect 25924 2360 25930 2372
rect 26237 2363 26295 2369
rect 26237 2360 26249 2363
rect 25924 2332 26249 2360
rect 25924 2320 25930 2332
rect 26237 2329 26249 2332
rect 26283 2329 26295 2363
rect 26237 2323 26295 2329
rect 27338 2320 27344 2372
rect 27396 2360 27402 2372
rect 27709 2363 27767 2369
rect 27709 2360 27721 2363
rect 27396 2332 27721 2360
rect 27396 2320 27402 2332
rect 27709 2329 27721 2332
rect 27755 2329 27767 2363
rect 27709 2323 27767 2329
rect 28810 2320 28816 2372
rect 28868 2360 28874 2372
rect 30009 2363 30067 2369
rect 30009 2360 30021 2363
rect 28868 2332 30021 2360
rect 28868 2320 28874 2332
rect 30009 2329 30021 2332
rect 30055 2329 30067 2363
rect 30009 2323 30067 2329
rect 30282 2320 30288 2372
rect 30340 2360 30346 2372
rect 30929 2363 30987 2369
rect 30929 2360 30941 2363
rect 30340 2332 30941 2360
rect 30340 2320 30346 2332
rect 30929 2329 30941 2332
rect 30975 2329 30987 2363
rect 30929 2323 30987 2329
rect 31754 2320 31760 2372
rect 31812 2360 31818 2372
rect 32585 2363 32643 2369
rect 32585 2360 32597 2363
rect 31812 2332 32597 2360
rect 31812 2320 31818 2332
rect 32585 2329 32597 2332
rect 32631 2329 32643 2363
rect 32585 2323 32643 2329
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 17224 37408 17276 37460
rect 14280 37340 14332 37392
rect 14924 37340 14976 37392
rect 5448 37315 5500 37324
rect 5448 37281 5457 37315
rect 5457 37281 5491 37315
rect 5491 37281 5500 37315
rect 5448 37272 5500 37281
rect 13452 37272 13504 37324
rect 37188 37272 37240 37324
rect 5080 37204 5132 37256
rect 8392 37204 8444 37256
rect 11704 37204 11756 37256
rect 15200 37247 15252 37256
rect 15200 37213 15209 37247
rect 15209 37213 15243 37247
rect 15243 37213 15252 37247
rect 15200 37204 15252 37213
rect 18328 37204 18380 37256
rect 24952 37204 25004 37256
rect 28264 37204 28316 37256
rect 31760 37204 31812 37256
rect 34796 37204 34848 37256
rect 38200 37204 38252 37256
rect 22100 37179 22152 37188
rect 22100 37145 22109 37179
rect 22109 37145 22143 37179
rect 22143 37145 22152 37179
rect 22100 37136 22152 37145
rect 15292 37111 15344 37120
rect 15292 37077 15301 37111
rect 15301 37077 15335 37111
rect 15335 37077 15344 37111
rect 15292 37068 15344 37077
rect 18604 37111 18656 37120
rect 18604 37077 18613 37111
rect 18613 37077 18647 37111
rect 18647 37077 18656 37111
rect 18604 37068 18656 37077
rect 22192 37111 22244 37120
rect 22192 37077 22201 37111
rect 22201 37077 22235 37111
rect 22235 37077 22244 37111
rect 22192 37068 22244 37077
rect 25228 37111 25280 37120
rect 25228 37077 25237 37111
rect 25237 37077 25271 37111
rect 25271 37077 25280 37111
rect 25228 37068 25280 37077
rect 34520 37068 34572 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 13452 36864 13504 36916
rect 22192 36864 22244 36916
rect 19432 36796 19484 36848
rect 18696 36728 18748 36780
rect 20076 36728 20128 36780
rect 25136 36771 25188 36780
rect 25136 36737 25145 36771
rect 25145 36737 25179 36771
rect 25179 36737 25188 36771
rect 25136 36728 25188 36737
rect 25504 36728 25556 36780
rect 26148 36771 26200 36780
rect 26148 36737 26157 36771
rect 26157 36737 26191 36771
rect 26191 36737 26200 36771
rect 26148 36728 26200 36737
rect 14464 36703 14516 36712
rect 14464 36669 14473 36703
rect 14473 36669 14507 36703
rect 14507 36669 14516 36703
rect 14464 36660 14516 36669
rect 25044 36703 25096 36712
rect 25044 36669 25053 36703
rect 25053 36669 25087 36703
rect 25087 36669 25096 36703
rect 25044 36660 25096 36669
rect 31024 36728 31076 36780
rect 31208 36660 31260 36712
rect 26056 36592 26108 36644
rect 13820 36567 13872 36576
rect 13820 36533 13829 36567
rect 13829 36533 13863 36567
rect 13863 36533 13872 36567
rect 13820 36524 13872 36533
rect 25872 36524 25924 36576
rect 30104 36567 30156 36576
rect 30104 36533 30113 36567
rect 30113 36533 30147 36567
rect 30147 36533 30156 36567
rect 30104 36524 30156 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 26148 36320 26200 36372
rect 30380 36320 30432 36372
rect 31024 36363 31076 36372
rect 31024 36329 31033 36363
rect 31033 36329 31067 36363
rect 31067 36329 31076 36363
rect 31024 36320 31076 36329
rect 14188 36252 14240 36304
rect 15752 36252 15804 36304
rect 14924 36227 14976 36236
rect 14924 36193 14933 36227
rect 14933 36193 14967 36227
rect 14967 36193 14976 36227
rect 14924 36184 14976 36193
rect 17224 36227 17276 36236
rect 17224 36193 17233 36227
rect 17233 36193 17267 36227
rect 17267 36193 17276 36227
rect 17224 36184 17276 36193
rect 18604 36184 18656 36236
rect 25872 36227 25924 36236
rect 25872 36193 25881 36227
rect 25881 36193 25915 36227
rect 25915 36193 25924 36227
rect 25872 36184 25924 36193
rect 26056 36227 26108 36236
rect 26056 36193 26065 36227
rect 26065 36193 26099 36227
rect 26099 36193 26108 36227
rect 26056 36184 26108 36193
rect 17408 36116 17460 36168
rect 24768 36159 24820 36168
rect 24768 36125 24777 36159
rect 24777 36125 24811 36159
rect 24811 36125 24820 36159
rect 24768 36116 24820 36125
rect 33232 36227 33284 36236
rect 33232 36193 33241 36227
rect 33241 36193 33275 36227
rect 33275 36193 33284 36227
rect 33232 36184 33284 36193
rect 14464 36048 14516 36100
rect 17776 36048 17828 36100
rect 15292 35980 15344 36032
rect 29092 36116 29144 36168
rect 26148 36048 26200 36100
rect 29460 36048 29512 36100
rect 30380 36116 30432 36168
rect 31392 36116 31444 36168
rect 33416 36116 33468 36168
rect 34520 36116 34572 36168
rect 37188 36159 37240 36168
rect 37188 36125 37197 36159
rect 37197 36125 37231 36159
rect 37231 36125 37240 36159
rect 37188 36116 37240 36125
rect 30472 36048 30524 36100
rect 29184 36023 29236 36032
rect 29184 35989 29193 36023
rect 29193 35989 29227 36023
rect 29227 35989 29236 36023
rect 29184 35980 29236 35989
rect 30288 35980 30340 36032
rect 30840 36023 30892 36032
rect 30840 35989 30865 36023
rect 30865 35989 30892 36023
rect 30840 35980 30892 35989
rect 34060 35980 34112 36032
rect 34244 36023 34296 36032
rect 34244 35989 34253 36023
rect 34253 35989 34287 36023
rect 34287 35989 34296 36023
rect 34244 35980 34296 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 14280 35819 14332 35828
rect 14280 35785 14289 35819
rect 14289 35785 14323 35819
rect 14323 35785 14332 35819
rect 14280 35776 14332 35785
rect 22836 35708 22888 35760
rect 18788 35683 18840 35692
rect 18788 35649 18797 35683
rect 18797 35649 18831 35683
rect 18831 35649 18840 35683
rect 18788 35640 18840 35649
rect 19432 35683 19484 35692
rect 19432 35649 19441 35683
rect 19441 35649 19475 35683
rect 19475 35649 19484 35683
rect 19432 35640 19484 35649
rect 21180 35640 21232 35692
rect 14464 35615 14516 35624
rect 14464 35581 14473 35615
rect 14473 35581 14507 35615
rect 14507 35581 14516 35615
rect 14464 35572 14516 35581
rect 20536 35572 20588 35624
rect 22008 35640 22060 35692
rect 25136 35776 25188 35828
rect 30472 35776 30524 35828
rect 23112 35708 23164 35760
rect 25228 35708 25280 35760
rect 30288 35751 30340 35760
rect 23204 35683 23256 35692
rect 23204 35649 23213 35683
rect 23213 35649 23247 35683
rect 23247 35649 23256 35683
rect 23204 35640 23256 35649
rect 23388 35683 23440 35692
rect 23388 35649 23397 35683
rect 23397 35649 23431 35683
rect 23431 35649 23440 35683
rect 23388 35640 23440 35649
rect 29460 35640 29512 35692
rect 30288 35717 30297 35751
rect 30297 35717 30331 35751
rect 30331 35717 30340 35751
rect 30288 35708 30340 35717
rect 30380 35640 30432 35692
rect 30472 35640 30524 35692
rect 31392 35751 31444 35760
rect 31392 35717 31401 35751
rect 31401 35717 31435 35751
rect 31435 35717 31444 35751
rect 31392 35708 31444 35717
rect 22652 35615 22704 35624
rect 22652 35581 22661 35615
rect 22661 35581 22695 35615
rect 22695 35581 22704 35615
rect 22652 35572 22704 35581
rect 23756 35572 23808 35624
rect 24768 35572 24820 35624
rect 24952 35615 25004 35624
rect 24952 35581 24961 35615
rect 24961 35581 24995 35615
rect 24995 35581 25004 35615
rect 24952 35572 25004 35581
rect 25504 35615 25556 35624
rect 25504 35581 25513 35615
rect 25513 35581 25547 35615
rect 25547 35581 25556 35615
rect 25504 35572 25556 35581
rect 23480 35547 23532 35556
rect 23480 35513 23489 35547
rect 23489 35513 23523 35547
rect 23523 35513 23532 35547
rect 23480 35504 23532 35513
rect 24216 35504 24268 35556
rect 29000 35572 29052 35624
rect 30840 35572 30892 35624
rect 32956 35683 33008 35692
rect 32956 35649 32965 35683
rect 32965 35649 32999 35683
rect 32999 35649 33008 35683
rect 32956 35640 33008 35649
rect 32128 35572 32180 35624
rect 34428 35640 34480 35692
rect 29644 35504 29696 35556
rect 33600 35504 33652 35556
rect 14096 35436 14148 35488
rect 25504 35436 25556 35488
rect 31208 35479 31260 35488
rect 31208 35445 31217 35479
rect 31217 35445 31251 35479
rect 31251 35445 31260 35479
rect 31208 35436 31260 35445
rect 33140 35479 33192 35488
rect 33140 35445 33149 35479
rect 33149 35445 33183 35479
rect 33183 35445 33192 35479
rect 33140 35436 33192 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 20076 35275 20128 35284
rect 20076 35241 20085 35275
rect 20085 35241 20119 35275
rect 20119 35241 20128 35275
rect 20076 35232 20128 35241
rect 20352 35207 20404 35216
rect 20352 35173 20361 35207
rect 20361 35173 20395 35207
rect 20395 35173 20404 35207
rect 20352 35164 20404 35173
rect 20628 35232 20680 35284
rect 22652 35232 22704 35284
rect 23204 35275 23256 35284
rect 23204 35241 23213 35275
rect 23213 35241 23247 35275
rect 23247 35241 23256 35275
rect 23204 35232 23256 35241
rect 25044 35232 25096 35284
rect 30840 35232 30892 35284
rect 20720 35164 20772 35216
rect 29552 35164 29604 35216
rect 18696 35071 18748 35080
rect 18696 35037 18705 35071
rect 18705 35037 18739 35071
rect 18739 35037 18748 35071
rect 18696 35028 18748 35037
rect 20260 35071 20312 35080
rect 20260 35037 20269 35071
rect 20269 35037 20303 35071
rect 20303 35037 20312 35071
rect 20260 35028 20312 35037
rect 20812 35028 20864 35080
rect 21180 35071 21232 35080
rect 21180 35037 21189 35071
rect 21189 35037 21223 35071
rect 21223 35037 21232 35071
rect 21180 35028 21232 35037
rect 19064 34960 19116 35012
rect 20168 34960 20220 35012
rect 20076 34892 20128 34944
rect 20352 34892 20404 34944
rect 21916 35028 21968 35080
rect 22468 35071 22520 35080
rect 22468 35037 22477 35071
rect 22477 35037 22511 35071
rect 22511 35037 22520 35071
rect 22468 35028 22520 35037
rect 22652 35071 22704 35080
rect 22652 35037 22661 35071
rect 22661 35037 22695 35071
rect 22695 35037 22704 35071
rect 23388 35096 23440 35148
rect 29000 35096 29052 35148
rect 30012 35096 30064 35148
rect 30104 35096 30156 35148
rect 22652 35028 22704 35037
rect 23296 35071 23348 35080
rect 23296 35037 23305 35071
rect 23305 35037 23339 35071
rect 23339 35037 23348 35071
rect 23296 35028 23348 35037
rect 23480 35028 23532 35080
rect 24492 34960 24544 35012
rect 24768 35003 24820 35012
rect 24768 34969 24777 35003
rect 24777 34969 24811 35003
rect 24811 34969 24820 35003
rect 24768 34960 24820 34969
rect 25780 35028 25832 35080
rect 26792 35071 26844 35080
rect 26792 35037 26801 35071
rect 26801 35037 26835 35071
rect 26835 35037 26844 35071
rect 26792 35028 26844 35037
rect 29184 35028 29236 35080
rect 32128 35071 32180 35080
rect 32128 35037 32137 35071
rect 32137 35037 32171 35071
rect 32171 35037 32180 35071
rect 32128 35028 32180 35037
rect 32312 35096 32364 35148
rect 32956 35096 33008 35148
rect 33416 35096 33468 35148
rect 22468 34892 22520 34944
rect 23296 34892 23348 34944
rect 24676 34892 24728 34944
rect 30012 34892 30064 34944
rect 30840 34960 30892 35012
rect 33048 34960 33100 35012
rect 34060 35028 34112 35080
rect 33600 34960 33652 35012
rect 32956 34892 33008 34944
rect 35992 34935 36044 34944
rect 35992 34901 36001 34935
rect 36001 34901 36035 34935
rect 36035 34901 36044 34935
rect 35992 34892 36044 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 22652 34688 22704 34740
rect 30380 34688 30432 34740
rect 33232 34688 33284 34740
rect 20076 34620 20128 34672
rect 17408 34595 17460 34604
rect 17408 34561 17417 34595
rect 17417 34561 17451 34595
rect 17451 34561 17460 34595
rect 17408 34552 17460 34561
rect 18144 34595 18196 34604
rect 18144 34561 18153 34595
rect 18153 34561 18187 34595
rect 18187 34561 18196 34595
rect 18144 34552 18196 34561
rect 17224 34484 17276 34536
rect 18880 34552 18932 34604
rect 20260 34595 20312 34604
rect 20260 34561 20269 34595
rect 20269 34561 20303 34595
rect 20303 34561 20312 34595
rect 20260 34552 20312 34561
rect 20352 34595 20404 34604
rect 20352 34561 20361 34595
rect 20361 34561 20395 34595
rect 20395 34561 20404 34595
rect 20352 34552 20404 34561
rect 20628 34552 20680 34604
rect 21180 34620 21232 34672
rect 21364 34595 21416 34604
rect 21364 34561 21373 34595
rect 21373 34561 21407 34595
rect 21407 34561 21416 34595
rect 21364 34552 21416 34561
rect 22008 34595 22060 34604
rect 22008 34561 22017 34595
rect 22017 34561 22051 34595
rect 22051 34561 22060 34595
rect 22008 34552 22060 34561
rect 23756 34620 23808 34672
rect 24216 34595 24268 34604
rect 24216 34561 24225 34595
rect 24225 34561 24259 34595
rect 24259 34561 24268 34595
rect 24216 34552 24268 34561
rect 24492 34552 24544 34604
rect 25044 34620 25096 34672
rect 24676 34552 24728 34604
rect 32404 34620 32456 34672
rect 33048 34620 33100 34672
rect 29552 34552 29604 34604
rect 30840 34552 30892 34604
rect 32312 34595 32364 34604
rect 32312 34561 32321 34595
rect 32321 34561 32355 34595
rect 32355 34561 32364 34595
rect 32312 34552 32364 34561
rect 33140 34595 33192 34604
rect 33140 34561 33149 34595
rect 33149 34561 33183 34595
rect 33183 34561 33192 34595
rect 33140 34552 33192 34561
rect 22100 34484 22152 34536
rect 22192 34416 22244 34468
rect 23296 34484 23348 34536
rect 26424 34484 26476 34536
rect 32128 34484 32180 34536
rect 32772 34484 32824 34536
rect 24216 34416 24268 34468
rect 33876 34416 33928 34468
rect 21548 34348 21600 34400
rect 25688 34348 25740 34400
rect 32404 34391 32456 34400
rect 32404 34357 32413 34391
rect 32413 34357 32447 34391
rect 32447 34357 32456 34391
rect 32404 34348 32456 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 20720 34144 20772 34196
rect 32772 34187 32824 34196
rect 32772 34153 32781 34187
rect 32781 34153 32815 34187
rect 32815 34153 32824 34187
rect 32772 34144 32824 34153
rect 18880 34076 18932 34128
rect 21548 34076 21600 34128
rect 26792 34119 26844 34128
rect 26792 34085 26801 34119
rect 26801 34085 26835 34119
rect 26835 34085 26844 34119
rect 26792 34076 26844 34085
rect 17224 33983 17276 33992
rect 17224 33949 17233 33983
rect 17233 33949 17267 33983
rect 17267 33949 17276 33983
rect 17224 33940 17276 33949
rect 17408 33983 17460 33992
rect 17408 33949 17417 33983
rect 17417 33949 17451 33983
rect 17451 33949 17460 33983
rect 18788 34008 18840 34060
rect 20628 34008 20680 34060
rect 17408 33940 17460 33949
rect 18052 33983 18104 33992
rect 18052 33949 18061 33983
rect 18061 33949 18095 33983
rect 18095 33949 18104 33983
rect 18052 33940 18104 33949
rect 18144 33872 18196 33924
rect 18328 33940 18380 33992
rect 21364 33983 21416 33992
rect 21364 33949 21373 33983
rect 21373 33949 21407 33983
rect 21407 33949 21416 33983
rect 21364 33940 21416 33949
rect 24768 34008 24820 34060
rect 21916 33983 21968 33992
rect 21916 33949 21925 33983
rect 21925 33949 21959 33983
rect 21959 33949 21968 33983
rect 21916 33940 21968 33949
rect 22192 33983 22244 33992
rect 22192 33949 22201 33983
rect 22201 33949 22235 33983
rect 22235 33949 22244 33983
rect 22192 33940 22244 33949
rect 24952 33940 25004 33992
rect 23020 33872 23072 33924
rect 25688 33940 25740 33992
rect 26424 33983 26476 33992
rect 26148 33872 26200 33924
rect 26424 33949 26433 33983
rect 26433 33949 26467 33983
rect 26467 33949 26476 33983
rect 26424 33940 26476 33949
rect 31668 33940 31720 33992
rect 27252 33872 27304 33924
rect 32496 33915 32548 33924
rect 32496 33881 32505 33915
rect 32505 33881 32539 33915
rect 32539 33881 32548 33915
rect 32496 33872 32548 33881
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 25044 33643 25096 33652
rect 17408 33532 17460 33584
rect 25044 33609 25053 33643
rect 25053 33609 25087 33643
rect 25087 33609 25096 33643
rect 25044 33600 25096 33609
rect 32312 33600 32364 33652
rect 18696 33532 18748 33584
rect 17224 33507 17276 33516
rect 17224 33473 17233 33507
rect 17233 33473 17267 33507
rect 17267 33473 17276 33507
rect 17224 33464 17276 33473
rect 17500 33507 17552 33516
rect 17500 33473 17509 33507
rect 17509 33473 17543 33507
rect 17543 33473 17552 33507
rect 17500 33464 17552 33473
rect 17592 33464 17644 33516
rect 18052 33464 18104 33516
rect 20628 33532 20680 33584
rect 19064 33507 19116 33516
rect 19064 33473 19073 33507
rect 19073 33473 19107 33507
rect 19107 33473 19116 33507
rect 19064 33464 19116 33473
rect 26424 33507 26476 33516
rect 26424 33473 26433 33507
rect 26433 33473 26467 33507
rect 26467 33473 26476 33507
rect 26424 33464 26476 33473
rect 27896 33507 27948 33516
rect 18144 33439 18196 33448
rect 18144 33405 18153 33439
rect 18153 33405 18187 33439
rect 18187 33405 18196 33439
rect 18144 33396 18196 33405
rect 25412 33439 25464 33448
rect 17500 33328 17552 33380
rect 25412 33405 25421 33439
rect 25421 33405 25455 33439
rect 25455 33405 25464 33439
rect 25412 33396 25464 33405
rect 25964 33396 26016 33448
rect 27896 33473 27905 33507
rect 27905 33473 27939 33507
rect 27939 33473 27948 33507
rect 27896 33464 27948 33473
rect 28908 33532 28960 33584
rect 29552 33464 29604 33516
rect 29736 33507 29788 33516
rect 29736 33473 29745 33507
rect 29745 33473 29779 33507
rect 29779 33473 29788 33507
rect 29736 33464 29788 33473
rect 32404 33532 32456 33584
rect 32496 33464 32548 33516
rect 31668 33396 31720 33448
rect 24952 33328 25004 33380
rect 27436 33260 27488 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 17224 33056 17276 33108
rect 24768 33056 24820 33108
rect 25780 33099 25832 33108
rect 25780 33065 25789 33099
rect 25789 33065 25823 33099
rect 25823 33065 25832 33099
rect 25780 33056 25832 33065
rect 27896 33056 27948 33108
rect 19340 32988 19392 33040
rect 23112 32988 23164 33040
rect 25412 32988 25464 33040
rect 26148 32988 26200 33040
rect 26240 32988 26292 33040
rect 18144 32963 18196 32972
rect 18144 32929 18153 32963
rect 18153 32929 18187 32963
rect 18187 32929 18196 32963
rect 18144 32920 18196 32929
rect 17684 32784 17736 32836
rect 23020 32852 23072 32904
rect 24860 32895 24912 32904
rect 24860 32861 24869 32895
rect 24869 32861 24903 32895
rect 24903 32861 24912 32895
rect 24860 32852 24912 32861
rect 25320 32895 25372 32904
rect 25320 32861 25329 32895
rect 25329 32861 25363 32895
rect 25363 32861 25372 32895
rect 25320 32852 25372 32861
rect 25964 32895 26016 32904
rect 25964 32861 25973 32895
rect 25973 32861 26007 32895
rect 26007 32861 26016 32895
rect 25964 32852 26016 32861
rect 26148 32852 26200 32904
rect 29736 32988 29788 33040
rect 27160 32895 27212 32904
rect 27160 32861 27169 32895
rect 27169 32861 27203 32895
rect 27203 32861 27212 32895
rect 27160 32852 27212 32861
rect 27252 32895 27304 32904
rect 27252 32861 27261 32895
rect 27261 32861 27295 32895
rect 27295 32861 27304 32895
rect 27436 32895 27488 32904
rect 27252 32852 27304 32861
rect 27436 32861 27445 32895
rect 27445 32861 27479 32895
rect 27479 32861 27488 32895
rect 27436 32852 27488 32861
rect 27528 32895 27580 32904
rect 27528 32861 27537 32895
rect 27537 32861 27571 32895
rect 27571 32861 27580 32895
rect 28080 32895 28132 32904
rect 27528 32852 27580 32861
rect 28080 32861 28089 32895
rect 28089 32861 28123 32895
rect 28123 32861 28132 32895
rect 28080 32852 28132 32861
rect 28632 32895 28684 32904
rect 28632 32861 28641 32895
rect 28641 32861 28675 32895
rect 28675 32861 28684 32895
rect 28632 32852 28684 32861
rect 26424 32784 26476 32836
rect 21272 32716 21324 32768
rect 22008 32716 22060 32768
rect 27252 32716 27304 32768
rect 27804 32716 27856 32768
rect 28632 32716 28684 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 17500 32555 17552 32564
rect 17500 32521 17509 32555
rect 17509 32521 17543 32555
rect 17543 32521 17552 32555
rect 17500 32512 17552 32521
rect 17592 32512 17644 32564
rect 26148 32512 26200 32564
rect 27528 32512 27580 32564
rect 18328 32487 18380 32496
rect 18328 32453 18337 32487
rect 18337 32453 18371 32487
rect 18371 32453 18380 32487
rect 18328 32444 18380 32453
rect 18880 32444 18932 32496
rect 21364 32444 21416 32496
rect 23020 32444 23072 32496
rect 23388 32444 23440 32496
rect 20812 32419 20864 32428
rect 20812 32385 20821 32419
rect 20821 32385 20855 32419
rect 20855 32385 20864 32419
rect 20812 32376 20864 32385
rect 21272 32376 21324 32428
rect 23112 32419 23164 32428
rect 23112 32385 23121 32419
rect 23121 32385 23155 32419
rect 23155 32385 23164 32419
rect 23112 32376 23164 32385
rect 24952 32444 25004 32496
rect 27344 32419 27396 32428
rect 27344 32385 27353 32419
rect 27353 32385 27387 32419
rect 27387 32385 27396 32419
rect 27344 32376 27396 32385
rect 28816 32419 28868 32428
rect 17868 32351 17920 32360
rect 17868 32317 17877 32351
rect 17877 32317 17911 32351
rect 17911 32317 17920 32351
rect 17868 32308 17920 32317
rect 18328 32308 18380 32360
rect 19156 32308 19208 32360
rect 26424 32240 26476 32292
rect 28816 32385 28825 32419
rect 28825 32385 28859 32419
rect 28859 32385 28868 32419
rect 28816 32376 28868 32385
rect 28356 32308 28408 32360
rect 29644 32376 29696 32428
rect 34428 32512 34480 32564
rect 34520 32444 34572 32496
rect 32956 32308 33008 32360
rect 35992 32376 36044 32428
rect 35348 32351 35400 32360
rect 31668 32240 31720 32292
rect 17868 32172 17920 32224
rect 33508 32172 33560 32224
rect 35348 32317 35357 32351
rect 35357 32317 35391 32351
rect 35391 32317 35400 32351
rect 35348 32308 35400 32317
rect 34612 32215 34664 32224
rect 34612 32181 34621 32215
rect 34621 32181 34655 32215
rect 34655 32181 34664 32215
rect 34612 32172 34664 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 17592 31968 17644 32020
rect 23204 31968 23256 32020
rect 17684 31943 17736 31952
rect 17684 31909 17693 31943
rect 17693 31909 17727 31943
rect 17727 31909 17736 31943
rect 17684 31900 17736 31909
rect 23388 31943 23440 31952
rect 23388 31909 23397 31943
rect 23397 31909 23431 31943
rect 23431 31909 23440 31943
rect 23388 31900 23440 31909
rect 24860 31968 24912 32020
rect 28080 31900 28132 31952
rect 17224 31832 17276 31884
rect 23112 31875 23164 31884
rect 5448 31764 5500 31816
rect 17408 31764 17460 31816
rect 17592 31764 17644 31816
rect 23112 31841 23121 31875
rect 23121 31841 23155 31875
rect 23155 31841 23164 31875
rect 23112 31832 23164 31841
rect 27712 31875 27764 31884
rect 27712 31841 27721 31875
rect 27721 31841 27755 31875
rect 27755 31841 27764 31875
rect 27712 31832 27764 31841
rect 33232 31832 33284 31884
rect 27160 31764 27212 31816
rect 27804 31807 27856 31816
rect 27804 31773 27813 31807
rect 27813 31773 27847 31807
rect 27847 31773 27856 31807
rect 27804 31764 27856 31773
rect 33508 31807 33560 31816
rect 33508 31773 33517 31807
rect 33517 31773 33551 31807
rect 33551 31773 33560 31807
rect 33508 31764 33560 31773
rect 34796 31832 34848 31884
rect 35440 31875 35492 31884
rect 35440 31841 35449 31875
rect 35449 31841 35483 31875
rect 35483 31841 35492 31875
rect 35440 31832 35492 31841
rect 33784 31764 33836 31816
rect 15108 31696 15160 31748
rect 34612 31764 34664 31816
rect 34060 31628 34112 31680
rect 34152 31628 34204 31680
rect 34612 31628 34664 31680
rect 35348 31628 35400 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 13820 31424 13872 31476
rect 17868 31424 17920 31476
rect 6736 31288 6788 31340
rect 12624 31331 12676 31340
rect 12624 31297 12633 31331
rect 12633 31297 12667 31331
rect 12667 31297 12676 31331
rect 12624 31288 12676 31297
rect 5540 31263 5592 31272
rect 5540 31229 5549 31263
rect 5549 31229 5583 31263
rect 5583 31229 5592 31263
rect 5540 31220 5592 31229
rect 15108 31331 15160 31340
rect 15108 31297 15117 31331
rect 15117 31297 15151 31331
rect 15151 31297 15160 31331
rect 17132 31331 17184 31340
rect 15108 31288 15160 31297
rect 17132 31297 17141 31331
rect 17141 31297 17175 31331
rect 17175 31297 17184 31331
rect 17132 31288 17184 31297
rect 20720 31356 20772 31408
rect 31024 31356 31076 31408
rect 34520 31399 34572 31408
rect 34520 31365 34529 31399
rect 34529 31365 34563 31399
rect 34563 31365 34572 31399
rect 34520 31356 34572 31365
rect 19984 31331 20036 31340
rect 15844 31220 15896 31272
rect 18880 31220 18932 31272
rect 19248 31220 19300 31272
rect 19984 31297 19993 31331
rect 19993 31297 20027 31331
rect 20027 31297 20036 31331
rect 19984 31288 20036 31297
rect 20536 31331 20588 31340
rect 20536 31297 20545 31331
rect 20545 31297 20579 31331
rect 20579 31297 20588 31331
rect 20536 31288 20588 31297
rect 22284 31288 22336 31340
rect 23572 31288 23624 31340
rect 30472 31288 30524 31340
rect 30656 31331 30708 31340
rect 30656 31297 30665 31331
rect 30665 31297 30699 31331
rect 30699 31297 30708 31331
rect 34060 31331 34112 31340
rect 30656 31288 30708 31297
rect 34060 31297 34069 31331
rect 34069 31297 34103 31331
rect 34103 31297 34112 31331
rect 34060 31288 34112 31297
rect 34152 31331 34204 31340
rect 34152 31297 34161 31331
rect 34161 31297 34195 31331
rect 34195 31297 34204 31331
rect 34152 31288 34204 31297
rect 20260 31263 20312 31272
rect 20260 31229 20269 31263
rect 20269 31229 20303 31263
rect 20303 31229 20312 31263
rect 20260 31220 20312 31229
rect 33784 31263 33836 31272
rect 33784 31229 33793 31263
rect 33793 31229 33827 31263
rect 33827 31229 33836 31263
rect 33784 31220 33836 31229
rect 6828 31152 6880 31204
rect 23204 31195 23256 31204
rect 23204 31161 23213 31195
rect 23213 31161 23247 31195
rect 23247 31161 23256 31195
rect 23204 31152 23256 31161
rect 34428 31152 34480 31204
rect 5448 31127 5500 31136
rect 5448 31093 5457 31127
rect 5457 31093 5491 31127
rect 5491 31093 5500 31127
rect 5448 31084 5500 31093
rect 12072 31084 12124 31136
rect 22376 31127 22428 31136
rect 22376 31093 22385 31127
rect 22385 31093 22419 31127
rect 22419 31093 22428 31127
rect 22376 31084 22428 31093
rect 29828 31084 29880 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 29644 30880 29696 30932
rect 14372 30855 14424 30864
rect 14372 30821 14381 30855
rect 14381 30821 14415 30855
rect 14415 30821 14424 30855
rect 14372 30812 14424 30821
rect 18236 30812 18288 30864
rect 19984 30812 20036 30864
rect 5264 30744 5316 30796
rect 10324 30744 10376 30796
rect 19248 30744 19300 30796
rect 4620 30719 4672 30728
rect 4620 30685 4629 30719
rect 4629 30685 4663 30719
rect 4663 30685 4672 30719
rect 4620 30676 4672 30685
rect 8484 30676 8536 30728
rect 12072 30676 12124 30728
rect 14556 30719 14608 30728
rect 6000 30651 6052 30660
rect 6000 30617 6009 30651
rect 6009 30617 6043 30651
rect 6043 30617 6052 30651
rect 6000 30608 6052 30617
rect 9772 30608 9824 30660
rect 14556 30685 14565 30719
rect 14565 30685 14599 30719
rect 14599 30685 14608 30719
rect 14556 30676 14608 30685
rect 15108 30676 15160 30728
rect 18144 30719 18196 30728
rect 18144 30685 18153 30719
rect 18153 30685 18187 30719
rect 18187 30685 18196 30719
rect 18144 30676 18196 30685
rect 18420 30719 18472 30728
rect 18420 30685 18429 30719
rect 18429 30685 18463 30719
rect 18463 30685 18472 30719
rect 18420 30676 18472 30685
rect 21180 30812 21232 30864
rect 29920 30812 29972 30864
rect 20812 30744 20864 30796
rect 20904 30719 20956 30728
rect 15844 30608 15896 30660
rect 20904 30685 20913 30719
rect 20913 30685 20947 30719
rect 20947 30685 20956 30719
rect 20904 30676 20956 30685
rect 29736 30744 29788 30796
rect 34152 30880 34204 30932
rect 35440 30855 35492 30864
rect 30472 30744 30524 30796
rect 20720 30608 20772 30660
rect 28080 30608 28132 30660
rect 30196 30719 30248 30728
rect 30196 30685 30205 30719
rect 30205 30685 30239 30719
rect 30239 30685 30248 30719
rect 30196 30676 30248 30685
rect 30564 30676 30616 30728
rect 31024 30719 31076 30728
rect 31024 30685 31033 30719
rect 31033 30685 31067 30719
rect 31067 30685 31076 30719
rect 31024 30676 31076 30685
rect 34612 30744 34664 30796
rect 34796 30744 34848 30796
rect 33876 30676 33928 30728
rect 35440 30821 35449 30855
rect 35449 30821 35483 30855
rect 35483 30821 35492 30855
rect 35440 30812 35492 30821
rect 33416 30608 33468 30660
rect 33692 30608 33744 30660
rect 9404 30540 9456 30592
rect 17960 30583 18012 30592
rect 17960 30549 17969 30583
rect 17969 30549 18003 30583
rect 18003 30549 18012 30583
rect 17960 30540 18012 30549
rect 18328 30583 18380 30592
rect 18328 30549 18337 30583
rect 18337 30549 18371 30583
rect 18371 30549 18380 30583
rect 18328 30540 18380 30549
rect 29184 30583 29236 30592
rect 29184 30549 29193 30583
rect 29193 30549 29227 30583
rect 29227 30549 29236 30583
rect 29184 30540 29236 30549
rect 29276 30540 29328 30592
rect 29920 30540 29972 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4620 30336 4672 30388
rect 18788 30336 18840 30388
rect 19064 30336 19116 30388
rect 5448 30311 5500 30320
rect 5448 30277 5457 30311
rect 5457 30277 5491 30311
rect 5491 30277 5500 30311
rect 5448 30268 5500 30277
rect 6736 30311 6788 30320
rect 6736 30277 6745 30311
rect 6745 30277 6779 30311
rect 6779 30277 6788 30311
rect 6736 30268 6788 30277
rect 7104 30268 7156 30320
rect 6368 30200 6420 30252
rect 6460 30200 6512 30252
rect 6828 30243 6880 30252
rect 6828 30209 6837 30243
rect 6837 30209 6871 30243
rect 6871 30209 6880 30243
rect 6828 30200 6880 30209
rect 8392 30200 8444 30252
rect 9772 30268 9824 30320
rect 14372 30268 14424 30320
rect 18144 30268 18196 30320
rect 20720 30336 20772 30388
rect 10968 30243 11020 30252
rect 6000 30132 6052 30184
rect 6644 30132 6696 30184
rect 8852 30132 8904 30184
rect 10968 30209 10977 30243
rect 10977 30209 11011 30243
rect 11011 30209 11020 30243
rect 10968 30200 11020 30209
rect 10784 30132 10836 30184
rect 11152 30064 11204 30116
rect 5724 29996 5776 30048
rect 6920 29996 6972 30048
rect 11060 30039 11112 30048
rect 11060 30005 11069 30039
rect 11069 30005 11103 30039
rect 11103 30005 11112 30039
rect 11060 29996 11112 30005
rect 12716 30132 12768 30184
rect 14096 30132 14148 30184
rect 15200 30200 15252 30252
rect 16672 30200 16724 30252
rect 17132 30243 17184 30252
rect 17132 30209 17141 30243
rect 17141 30209 17175 30243
rect 17175 30209 17184 30243
rect 17132 30200 17184 30209
rect 17408 30200 17460 30252
rect 17960 30200 18012 30252
rect 22284 30268 22336 30320
rect 29184 30268 29236 30320
rect 20720 30243 20772 30252
rect 20720 30209 20729 30243
rect 20729 30209 20763 30243
rect 20763 30209 20772 30243
rect 20720 30200 20772 30209
rect 21272 30243 21324 30252
rect 21272 30209 21281 30243
rect 21281 30209 21315 30243
rect 21315 30209 21324 30243
rect 21272 30200 21324 30209
rect 24308 30243 24360 30252
rect 24308 30209 24317 30243
rect 24317 30209 24351 30243
rect 24351 30209 24360 30243
rect 24308 30200 24360 30209
rect 24952 30200 25004 30252
rect 28172 30243 28224 30252
rect 28172 30209 28181 30243
rect 28181 30209 28215 30243
rect 28215 30209 28224 30243
rect 28172 30200 28224 30209
rect 29276 30200 29328 30252
rect 29920 30268 29972 30320
rect 18696 30132 18748 30184
rect 18880 30132 18932 30184
rect 20260 30132 20312 30184
rect 22376 30132 22428 30184
rect 25320 30132 25372 30184
rect 25964 30132 26016 30184
rect 28080 30132 28132 30184
rect 29828 30243 29880 30252
rect 29828 30209 29837 30243
rect 29837 30209 29871 30243
rect 29871 30209 29880 30243
rect 29828 30200 29880 30209
rect 30564 30243 30616 30252
rect 30564 30209 30573 30243
rect 30573 30209 30607 30243
rect 30607 30209 30616 30243
rect 30564 30200 30616 30209
rect 31024 30268 31076 30320
rect 32220 30200 32272 30252
rect 32956 30243 33008 30252
rect 32404 30132 32456 30184
rect 32956 30209 32965 30243
rect 32965 30209 32999 30243
rect 32999 30209 33008 30243
rect 32956 30200 33008 30209
rect 33140 30200 33192 30252
rect 33876 30336 33928 30388
rect 33692 30268 33744 30320
rect 18604 30064 18656 30116
rect 14832 29996 14884 30048
rect 23940 29996 23992 30048
rect 27988 29996 28040 30048
rect 28356 30064 28408 30116
rect 29736 29996 29788 30048
rect 33324 30064 33376 30116
rect 34428 30200 34480 30252
rect 34244 29996 34296 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 6460 29835 6512 29844
rect 6460 29801 6469 29835
rect 6469 29801 6503 29835
rect 6503 29801 6512 29835
rect 6460 29792 6512 29801
rect 6644 29792 6696 29844
rect 6736 29792 6788 29844
rect 6828 29792 6880 29844
rect 5356 29656 5408 29708
rect 7104 29724 7156 29776
rect 8024 29724 8076 29776
rect 10784 29792 10836 29844
rect 18420 29792 18472 29844
rect 8300 29767 8352 29776
rect 8300 29733 8309 29767
rect 8309 29733 8343 29767
rect 8343 29733 8352 29767
rect 8300 29724 8352 29733
rect 9680 29724 9732 29776
rect 4988 29588 5040 29640
rect 5540 29588 5592 29640
rect 9772 29656 9824 29708
rect 8484 29631 8536 29640
rect 6092 29520 6144 29572
rect 8484 29597 8493 29631
rect 8493 29597 8527 29631
rect 8527 29597 8536 29631
rect 8484 29588 8536 29597
rect 9312 29631 9364 29640
rect 5172 29452 5224 29504
rect 5448 29452 5500 29504
rect 8024 29520 8076 29572
rect 9312 29597 9321 29631
rect 9321 29597 9355 29631
rect 9355 29597 9364 29631
rect 9312 29588 9364 29597
rect 10968 29724 11020 29776
rect 11152 29767 11204 29776
rect 11152 29733 11161 29767
rect 11161 29733 11195 29767
rect 11195 29733 11204 29767
rect 11152 29724 11204 29733
rect 10324 29631 10376 29640
rect 10324 29597 10333 29631
rect 10333 29597 10367 29631
rect 10367 29597 10376 29631
rect 10324 29588 10376 29597
rect 10968 29588 11020 29640
rect 13820 29656 13872 29708
rect 10232 29520 10284 29572
rect 14464 29588 14516 29640
rect 14832 29631 14884 29640
rect 14832 29597 14841 29631
rect 14841 29597 14875 29631
rect 14875 29597 14884 29631
rect 14832 29588 14884 29597
rect 14924 29520 14976 29572
rect 13360 29452 13412 29504
rect 14280 29452 14332 29504
rect 14464 29452 14516 29504
rect 15108 29452 15160 29504
rect 15752 29631 15804 29640
rect 15752 29597 15761 29631
rect 15761 29597 15795 29631
rect 15795 29597 15804 29631
rect 15752 29588 15804 29597
rect 18144 29656 18196 29708
rect 18236 29588 18288 29640
rect 18788 29656 18840 29708
rect 19984 29724 20036 29776
rect 20168 29724 20220 29776
rect 24952 29835 25004 29844
rect 22100 29724 22152 29776
rect 23572 29724 23624 29776
rect 24952 29801 24961 29835
rect 24961 29801 24995 29835
rect 24995 29801 25004 29835
rect 24952 29792 25004 29801
rect 29276 29792 29328 29844
rect 30196 29792 30248 29844
rect 30564 29792 30616 29844
rect 20904 29699 20956 29708
rect 19340 29588 19392 29640
rect 20904 29665 20913 29699
rect 20913 29665 20947 29699
rect 20947 29665 20956 29699
rect 20904 29656 20956 29665
rect 23756 29699 23808 29708
rect 23756 29665 23765 29699
rect 23765 29665 23799 29699
rect 23799 29665 23808 29699
rect 23756 29656 23808 29665
rect 23940 29699 23992 29708
rect 23940 29665 23949 29699
rect 23949 29665 23983 29699
rect 23983 29665 23992 29699
rect 23940 29656 23992 29665
rect 18328 29452 18380 29504
rect 19984 29631 20036 29640
rect 19984 29597 19993 29631
rect 19993 29597 20027 29631
rect 20027 29597 20036 29631
rect 19984 29588 20036 29597
rect 20076 29520 20128 29572
rect 20352 29520 20404 29572
rect 23480 29588 23532 29640
rect 23664 29631 23716 29640
rect 23664 29597 23673 29631
rect 23673 29597 23707 29631
rect 23707 29597 23716 29631
rect 23664 29588 23716 29597
rect 23848 29631 23900 29640
rect 23848 29597 23857 29631
rect 23857 29597 23891 29631
rect 23891 29597 23900 29631
rect 25596 29724 25648 29776
rect 24584 29656 24636 29708
rect 26056 29699 26108 29708
rect 23848 29588 23900 29597
rect 23388 29520 23440 29572
rect 22836 29452 22888 29504
rect 24676 29520 24728 29572
rect 26056 29665 26065 29699
rect 26065 29665 26099 29699
rect 26099 29665 26108 29699
rect 26056 29656 26108 29665
rect 28356 29724 28408 29776
rect 33232 29792 33284 29844
rect 25964 29631 26016 29640
rect 25964 29597 25973 29631
rect 25973 29597 26007 29631
rect 26007 29597 26016 29631
rect 25964 29588 26016 29597
rect 27988 29588 28040 29640
rect 29184 29656 29236 29708
rect 29736 29631 29788 29640
rect 28724 29520 28776 29572
rect 29736 29597 29745 29631
rect 29745 29597 29779 29631
rect 29779 29597 29788 29631
rect 29736 29588 29788 29597
rect 31668 29520 31720 29572
rect 25872 29452 25924 29504
rect 27712 29452 27764 29504
rect 27804 29452 27856 29504
rect 29552 29452 29604 29504
rect 29828 29452 29880 29504
rect 32956 29724 33008 29776
rect 32220 29631 32272 29640
rect 32220 29597 32229 29631
rect 32229 29597 32263 29631
rect 32263 29597 32272 29631
rect 32220 29588 32272 29597
rect 32404 29631 32456 29640
rect 32404 29597 32413 29631
rect 32413 29597 32447 29631
rect 32447 29597 32456 29631
rect 32404 29588 32456 29597
rect 33140 29631 33192 29640
rect 33140 29597 33149 29631
rect 33149 29597 33183 29631
rect 33183 29597 33192 29631
rect 33140 29588 33192 29597
rect 33232 29631 33284 29640
rect 33232 29597 33241 29631
rect 33241 29597 33275 29631
rect 33275 29597 33284 29631
rect 33232 29588 33284 29597
rect 33692 29588 33744 29640
rect 33324 29520 33376 29572
rect 33508 29452 33560 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 5080 29248 5132 29300
rect 6000 29248 6052 29300
rect 6368 29248 6420 29300
rect 8392 29291 8444 29300
rect 5172 29180 5224 29232
rect 4988 29155 5040 29164
rect 4988 29121 4997 29155
rect 4997 29121 5031 29155
rect 5031 29121 5040 29155
rect 4988 29112 5040 29121
rect 5448 29155 5500 29164
rect 5448 29121 5457 29155
rect 5457 29121 5491 29155
rect 5491 29121 5500 29155
rect 5448 29112 5500 29121
rect 5540 29112 5592 29164
rect 8116 29180 8168 29232
rect 6920 29155 6972 29164
rect 6920 29121 6929 29155
rect 6929 29121 6963 29155
rect 6963 29121 6972 29155
rect 8392 29257 8401 29291
rect 8401 29257 8435 29291
rect 8435 29257 8444 29291
rect 8392 29248 8444 29257
rect 9312 29248 9364 29300
rect 10324 29248 10376 29300
rect 18788 29291 18840 29300
rect 18788 29257 18797 29291
rect 18797 29257 18831 29291
rect 18831 29257 18840 29291
rect 18788 29248 18840 29257
rect 14464 29180 14516 29232
rect 6920 29112 6972 29121
rect 6092 29044 6144 29096
rect 7748 29044 7800 29096
rect 9220 29087 9272 29096
rect 5356 29019 5408 29028
rect 5356 28985 5365 29019
rect 5365 28985 5399 29019
rect 5399 28985 5408 29019
rect 5356 28976 5408 28985
rect 5264 28908 5316 28960
rect 7932 28976 7984 29028
rect 9220 29053 9229 29087
rect 9229 29053 9263 29087
rect 9263 29053 9272 29087
rect 9220 29044 9272 29053
rect 14280 29112 14332 29164
rect 19432 29248 19484 29300
rect 20260 29248 20312 29300
rect 23756 29291 23808 29300
rect 23756 29257 23765 29291
rect 23765 29257 23799 29291
rect 23799 29257 23808 29291
rect 23756 29248 23808 29257
rect 23940 29291 23992 29300
rect 23940 29257 23949 29291
rect 23949 29257 23983 29291
rect 23983 29257 23992 29291
rect 23940 29248 23992 29257
rect 24768 29248 24820 29300
rect 24860 29248 24912 29300
rect 25872 29248 25924 29300
rect 28080 29291 28132 29300
rect 19156 29155 19208 29164
rect 19156 29121 19165 29155
rect 19165 29121 19199 29155
rect 19199 29121 19208 29155
rect 19156 29112 19208 29121
rect 18604 29044 18656 29096
rect 13820 28976 13872 29028
rect 14924 28976 14976 29028
rect 17408 28976 17460 29028
rect 19248 29087 19300 29096
rect 19248 29053 19257 29087
rect 19257 29053 19291 29087
rect 19291 29053 19300 29087
rect 19248 29044 19300 29053
rect 20076 29044 20128 29096
rect 20352 29155 20404 29164
rect 20352 29121 20361 29155
rect 20361 29121 20395 29155
rect 20395 29121 20404 29155
rect 22376 29180 22428 29232
rect 23664 29180 23716 29232
rect 25596 29223 25648 29232
rect 20352 29112 20404 29121
rect 20628 29112 20680 29164
rect 24676 29112 24728 29164
rect 24952 29112 25004 29164
rect 25596 29189 25605 29223
rect 25605 29189 25639 29223
rect 25639 29189 25648 29223
rect 25596 29180 25648 29189
rect 28080 29257 28089 29291
rect 28089 29257 28123 29291
rect 28123 29257 28132 29291
rect 28080 29248 28132 29257
rect 25872 29155 25924 29164
rect 25872 29121 25881 29155
rect 25881 29121 25915 29155
rect 25915 29121 25924 29155
rect 25872 29112 25924 29121
rect 21272 29044 21324 29096
rect 10600 28908 10652 28960
rect 20168 28976 20220 29028
rect 20444 29019 20496 29028
rect 20444 28985 20453 29019
rect 20453 28985 20487 29019
rect 20487 28985 20496 29019
rect 22836 29019 22888 29028
rect 20444 28976 20496 28985
rect 22836 28985 22845 29019
rect 22845 28985 22879 29019
rect 22879 28985 22888 29019
rect 22836 28976 22888 28985
rect 23940 29044 23992 29096
rect 24032 29087 24084 29096
rect 24032 29053 24041 29087
rect 24041 29053 24075 29087
rect 24075 29053 24084 29087
rect 24032 29044 24084 29053
rect 24492 29044 24544 29096
rect 26056 29044 26108 29096
rect 19340 28908 19392 28960
rect 22376 28908 22428 28960
rect 24308 28976 24360 29028
rect 28724 29155 28776 29164
rect 28724 29121 28733 29155
rect 28733 29121 28767 29155
rect 28767 29121 28776 29155
rect 28724 29112 28776 29121
rect 29184 29044 29236 29096
rect 29276 29087 29328 29096
rect 29276 29053 29285 29087
rect 29285 29053 29319 29087
rect 29319 29053 29328 29087
rect 29276 29044 29328 29053
rect 24860 28908 24912 28960
rect 31116 28976 31168 29028
rect 33324 28976 33376 29028
rect 29092 28908 29144 28960
rect 29276 28908 29328 28960
rect 29736 28908 29788 28960
rect 33232 28908 33284 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 9220 28747 9272 28756
rect 9220 28713 9229 28747
rect 9229 28713 9263 28747
rect 9263 28713 9272 28747
rect 9220 28704 9272 28713
rect 10232 28704 10284 28756
rect 5540 28611 5592 28620
rect 5540 28577 5549 28611
rect 5549 28577 5583 28611
rect 5583 28577 5592 28611
rect 5540 28568 5592 28577
rect 6092 28611 6144 28620
rect 6092 28577 6101 28611
rect 6101 28577 6135 28611
rect 6135 28577 6144 28611
rect 6092 28568 6144 28577
rect 8300 28568 8352 28620
rect 6920 28500 6972 28552
rect 9404 28543 9456 28552
rect 9404 28509 9413 28543
rect 9413 28509 9447 28543
rect 9447 28509 9456 28543
rect 9404 28500 9456 28509
rect 9680 28543 9732 28552
rect 9680 28509 9715 28543
rect 9715 28509 9732 28543
rect 9864 28543 9916 28552
rect 9680 28500 9732 28509
rect 9864 28509 9873 28543
rect 9873 28509 9907 28543
rect 9907 28509 9916 28543
rect 9864 28500 9916 28509
rect 10324 28500 10376 28552
rect 11060 28704 11112 28756
rect 14924 28747 14976 28756
rect 14924 28713 14933 28747
rect 14933 28713 14967 28747
rect 14967 28713 14976 28747
rect 14924 28704 14976 28713
rect 19248 28704 19300 28756
rect 19984 28704 20036 28756
rect 20444 28704 20496 28756
rect 23940 28747 23992 28756
rect 23940 28713 23949 28747
rect 23949 28713 23983 28747
rect 23983 28713 23992 28747
rect 23940 28704 23992 28713
rect 29920 28747 29972 28756
rect 29920 28713 29929 28747
rect 29929 28713 29963 28747
rect 29963 28713 29972 28747
rect 29920 28704 29972 28713
rect 10784 28636 10836 28688
rect 27344 28636 27396 28688
rect 28264 28679 28316 28688
rect 28264 28645 28273 28679
rect 28273 28645 28307 28679
rect 28307 28645 28316 28679
rect 28264 28636 28316 28645
rect 29184 28636 29236 28688
rect 33508 28679 33560 28688
rect 33508 28645 33517 28679
rect 33517 28645 33551 28679
rect 33551 28645 33560 28679
rect 33508 28636 33560 28645
rect 34336 28568 34388 28620
rect 10600 28543 10652 28552
rect 10600 28509 10609 28543
rect 10609 28509 10643 28543
rect 10643 28509 10652 28543
rect 10600 28500 10652 28509
rect 6828 28432 6880 28484
rect 14740 28500 14792 28552
rect 18420 28500 18472 28552
rect 22744 28543 22796 28552
rect 22744 28509 22753 28543
rect 22753 28509 22787 28543
rect 22787 28509 22796 28543
rect 22744 28500 22796 28509
rect 19156 28432 19208 28484
rect 23572 28500 23624 28552
rect 24400 28500 24452 28552
rect 27712 28500 27764 28552
rect 33048 28500 33100 28552
rect 33416 28500 33468 28552
rect 5724 28407 5776 28416
rect 5724 28373 5733 28407
rect 5733 28373 5767 28407
rect 5767 28373 5776 28407
rect 5724 28364 5776 28373
rect 22560 28364 22612 28416
rect 24676 28432 24728 28484
rect 28724 28432 28776 28484
rect 29736 28475 29788 28484
rect 29736 28441 29745 28475
rect 29745 28441 29779 28475
rect 29779 28441 29788 28475
rect 29736 28432 29788 28441
rect 33324 28432 33376 28484
rect 25044 28364 25096 28416
rect 27620 28364 27672 28416
rect 28356 28364 28408 28416
rect 28816 28407 28868 28416
rect 28816 28373 28825 28407
rect 28825 28373 28859 28407
rect 28859 28373 28868 28407
rect 28816 28364 28868 28373
rect 29552 28364 29604 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 5264 28203 5316 28212
rect 5264 28169 5289 28203
rect 5289 28169 5316 28203
rect 5264 28160 5316 28169
rect 9864 28160 9916 28212
rect 19984 28160 20036 28212
rect 24768 28203 24820 28212
rect 5080 28135 5132 28144
rect 5080 28101 5089 28135
rect 5089 28101 5123 28135
rect 5123 28101 5132 28135
rect 5080 28092 5132 28101
rect 6920 28092 6972 28144
rect 16672 28092 16724 28144
rect 22560 28135 22612 28144
rect 22560 28101 22569 28135
rect 22569 28101 22603 28135
rect 22603 28101 22612 28135
rect 22560 28092 22612 28101
rect 24768 28169 24777 28203
rect 24777 28169 24811 28203
rect 24811 28169 24820 28203
rect 24768 28160 24820 28169
rect 29092 28203 29144 28212
rect 29092 28169 29101 28203
rect 29101 28169 29135 28203
rect 29135 28169 29144 28203
rect 29092 28160 29144 28169
rect 29920 28160 29972 28212
rect 5632 28024 5684 28076
rect 6828 28024 6880 28076
rect 8392 28024 8444 28076
rect 10324 28024 10376 28076
rect 16488 28024 16540 28076
rect 16764 28024 16816 28076
rect 22192 28067 22244 28076
rect 22192 28033 22201 28067
rect 22201 28033 22235 28067
rect 22235 28033 22244 28067
rect 22192 28024 22244 28033
rect 22376 28067 22428 28076
rect 22376 28033 22385 28067
rect 22385 28033 22419 28067
rect 22419 28033 22428 28067
rect 22376 28024 22428 28033
rect 24400 28067 24452 28076
rect 24400 28033 24409 28067
rect 24409 28033 24443 28067
rect 24443 28033 24452 28067
rect 24400 28024 24452 28033
rect 27620 28024 27672 28076
rect 28172 28067 28224 28076
rect 28172 28033 28181 28067
rect 28181 28033 28215 28067
rect 28215 28033 28224 28067
rect 28172 28024 28224 28033
rect 28448 28067 28500 28076
rect 28448 28033 28457 28067
rect 28457 28033 28491 28067
rect 28491 28033 28500 28067
rect 28448 28024 28500 28033
rect 28816 28024 28868 28076
rect 29276 28067 29328 28076
rect 29276 28033 29285 28067
rect 29285 28033 29319 28067
rect 29319 28033 29328 28067
rect 29276 28024 29328 28033
rect 29552 28067 29604 28076
rect 29552 28033 29561 28067
rect 29561 28033 29595 28067
rect 29595 28033 29604 28067
rect 29552 28024 29604 28033
rect 31116 28024 31168 28076
rect 33048 28092 33100 28144
rect 16028 27956 16080 28008
rect 22100 27888 22152 27940
rect 5172 27820 5224 27872
rect 5448 27863 5500 27872
rect 5448 27829 5457 27863
rect 5457 27829 5491 27863
rect 5491 27829 5500 27863
rect 5448 27820 5500 27829
rect 7748 27863 7800 27872
rect 7748 27829 7757 27863
rect 7757 27829 7791 27863
rect 7791 27829 7800 27863
rect 7748 27820 7800 27829
rect 15752 27820 15804 27872
rect 17040 27863 17092 27872
rect 17040 27829 17049 27863
rect 17049 27829 17083 27863
rect 17083 27829 17092 27863
rect 17040 27820 17092 27829
rect 28172 27820 28224 27872
rect 31852 28024 31904 28076
rect 33416 28067 33468 28076
rect 31484 27888 31536 27940
rect 31760 27956 31812 28008
rect 33416 28033 33425 28067
rect 33425 28033 33459 28067
rect 33459 28033 33468 28067
rect 33416 28024 33468 28033
rect 33140 27956 33192 28008
rect 33692 28024 33744 28076
rect 34336 28067 34388 28076
rect 34336 28033 34345 28067
rect 34345 28033 34379 28067
rect 34379 28033 34388 28067
rect 34336 28024 34388 28033
rect 33784 27999 33836 28008
rect 33784 27965 33793 27999
rect 33793 27965 33827 27999
rect 33827 27965 33836 27999
rect 33784 27956 33836 27965
rect 33048 27888 33100 27940
rect 32036 27820 32088 27872
rect 32312 27863 32364 27872
rect 32312 27829 32321 27863
rect 32321 27829 32355 27863
rect 32355 27829 32364 27863
rect 32312 27820 32364 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 5724 27548 5776 27600
rect 6920 27548 6972 27600
rect 18144 27548 18196 27600
rect 19432 27548 19484 27600
rect 29552 27616 29604 27668
rect 26240 27548 26292 27600
rect 27344 27548 27396 27600
rect 4528 27523 4580 27532
rect 4528 27489 4537 27523
rect 4537 27489 4571 27523
rect 4571 27489 4580 27523
rect 4528 27480 4580 27489
rect 14372 27480 14424 27532
rect 22744 27480 22796 27532
rect 24400 27480 24452 27532
rect 7104 27455 7156 27464
rect 7104 27421 7113 27455
rect 7113 27421 7147 27455
rect 7147 27421 7156 27455
rect 7104 27412 7156 27421
rect 14280 27412 14332 27464
rect 14464 27455 14516 27464
rect 14464 27421 14473 27455
rect 14473 27421 14507 27455
rect 14507 27421 14516 27455
rect 14464 27412 14516 27421
rect 14740 27455 14792 27464
rect 14740 27421 14749 27455
rect 14749 27421 14783 27455
rect 14783 27421 14792 27455
rect 14740 27412 14792 27421
rect 15476 27412 15528 27464
rect 16856 27412 16908 27464
rect 18512 27455 18564 27464
rect 4620 27344 4672 27396
rect 5448 27344 5500 27396
rect 18512 27421 18521 27455
rect 18521 27421 18555 27455
rect 18555 27421 18564 27455
rect 18512 27412 18564 27421
rect 18696 27344 18748 27396
rect 19984 27412 20036 27464
rect 22468 27412 22520 27464
rect 24032 27412 24084 27464
rect 28448 27523 28500 27532
rect 28448 27489 28457 27523
rect 28457 27489 28491 27523
rect 28491 27489 28500 27523
rect 28448 27480 28500 27489
rect 25320 27455 25372 27464
rect 25320 27421 25329 27455
rect 25329 27421 25363 27455
rect 25363 27421 25372 27455
rect 25320 27412 25372 27421
rect 20628 27344 20680 27396
rect 27712 27412 27764 27464
rect 28264 27412 28316 27464
rect 4712 27276 4764 27328
rect 17224 27276 17276 27328
rect 18052 27319 18104 27328
rect 18052 27285 18061 27319
rect 18061 27285 18095 27319
rect 18095 27285 18104 27319
rect 18052 27276 18104 27285
rect 18420 27319 18472 27328
rect 18420 27285 18429 27319
rect 18429 27285 18463 27319
rect 18463 27285 18472 27319
rect 18420 27276 18472 27285
rect 19340 27276 19392 27328
rect 24768 27319 24820 27328
rect 24768 27285 24777 27319
rect 24777 27285 24811 27319
rect 24811 27285 24820 27319
rect 24768 27276 24820 27285
rect 27620 27344 27672 27396
rect 28356 27387 28408 27396
rect 28356 27353 28365 27387
rect 28365 27353 28399 27387
rect 28399 27353 28408 27387
rect 28356 27344 28408 27353
rect 28724 27412 28776 27464
rect 32680 27548 32732 27600
rect 31484 27480 31536 27532
rect 33416 27616 33468 27668
rect 32036 27455 32088 27464
rect 32036 27421 32045 27455
rect 32045 27421 32079 27455
rect 32079 27421 32088 27455
rect 32036 27412 32088 27421
rect 32956 27455 33008 27464
rect 32956 27421 32965 27455
rect 32965 27421 32999 27455
rect 32999 27421 33008 27455
rect 32956 27412 33008 27421
rect 33048 27412 33100 27464
rect 32312 27344 32364 27396
rect 32772 27344 32824 27396
rect 31392 27276 31444 27328
rect 31668 27276 31720 27328
rect 33048 27276 33100 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 16120 27072 16172 27124
rect 18144 27072 18196 27124
rect 18420 27072 18472 27124
rect 22192 27072 22244 27124
rect 23388 27072 23440 27124
rect 25320 27072 25372 27124
rect 28724 27072 28776 27124
rect 32956 27072 33008 27124
rect 5080 27004 5132 27056
rect 15844 27047 15896 27056
rect 15844 27013 15853 27047
rect 15853 27013 15887 27047
rect 15887 27013 15896 27047
rect 15844 27004 15896 27013
rect 15936 27004 15988 27056
rect 4620 26979 4672 26988
rect 4620 26945 4629 26979
rect 4629 26945 4663 26979
rect 4663 26945 4672 26979
rect 4620 26936 4672 26945
rect 5632 26936 5684 26988
rect 13820 26936 13872 26988
rect 14280 26979 14332 26988
rect 4528 26868 4580 26920
rect 12532 26868 12584 26920
rect 13360 26911 13412 26920
rect 13360 26877 13369 26911
rect 13369 26877 13403 26911
rect 13403 26877 13412 26911
rect 13360 26868 13412 26877
rect 3148 26800 3200 26852
rect 5724 26800 5776 26852
rect 14280 26945 14289 26979
rect 14289 26945 14323 26979
rect 14323 26945 14332 26979
rect 14280 26936 14332 26945
rect 16948 26936 17000 26988
rect 18052 27004 18104 27056
rect 19432 26979 19484 26988
rect 19432 26945 19441 26979
rect 19441 26945 19475 26979
rect 19475 26945 19484 26979
rect 19432 26936 19484 26945
rect 14004 26911 14056 26920
rect 14004 26877 14013 26911
rect 14013 26877 14047 26911
rect 14047 26877 14056 26911
rect 14188 26911 14240 26920
rect 14004 26868 14056 26877
rect 14188 26877 14197 26911
rect 14197 26877 14231 26911
rect 14231 26877 14240 26911
rect 14188 26868 14240 26877
rect 19616 26868 19668 26920
rect 4620 26732 4672 26784
rect 10600 26732 10652 26784
rect 14004 26732 14056 26784
rect 14924 26732 14976 26784
rect 16120 26732 16172 26784
rect 16304 26732 16356 26784
rect 20076 26800 20128 26852
rect 18420 26732 18472 26784
rect 22100 26936 22152 26988
rect 22376 26936 22428 26988
rect 24216 26936 24268 26988
rect 32496 27004 32548 27056
rect 24768 26979 24820 26988
rect 24768 26945 24777 26979
rect 24777 26945 24811 26979
rect 24811 26945 24820 26979
rect 24768 26936 24820 26945
rect 24860 26936 24912 26988
rect 25136 26979 25188 26988
rect 25136 26945 25145 26979
rect 25145 26945 25179 26979
rect 25179 26945 25188 26979
rect 25136 26936 25188 26945
rect 27620 26936 27672 26988
rect 27896 26979 27948 26988
rect 27896 26945 27905 26979
rect 27905 26945 27939 26979
rect 27939 26945 27948 26979
rect 27896 26936 27948 26945
rect 27988 26979 28040 26988
rect 27988 26945 27997 26979
rect 27997 26945 28031 26979
rect 28031 26945 28040 26979
rect 28172 26979 28224 26988
rect 27988 26936 28040 26945
rect 28172 26945 28181 26979
rect 28181 26945 28215 26979
rect 28215 26945 28224 26979
rect 28172 26936 28224 26945
rect 28632 26936 28684 26988
rect 31392 26979 31444 26988
rect 31392 26945 31401 26979
rect 31401 26945 31435 26979
rect 31435 26945 31444 26979
rect 31392 26936 31444 26945
rect 31852 26936 31904 26988
rect 32588 26979 32640 26988
rect 32588 26945 32597 26979
rect 32597 26945 32631 26979
rect 32631 26945 32640 26979
rect 32588 26936 32640 26945
rect 23480 26868 23532 26920
rect 32864 26868 32916 26920
rect 33416 26911 33468 26920
rect 33416 26877 33425 26911
rect 33425 26877 33459 26911
rect 33459 26877 33468 26911
rect 33416 26868 33468 26877
rect 24860 26800 24912 26852
rect 25136 26800 25188 26852
rect 27436 26800 27488 26852
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 8484 26528 8536 26580
rect 4620 26435 4672 26444
rect 4620 26401 4629 26435
rect 4629 26401 4663 26435
rect 4663 26401 4672 26435
rect 4620 26392 4672 26401
rect 5816 26460 5868 26512
rect 3148 26256 3200 26308
rect 3976 26231 4028 26240
rect 3976 26197 3985 26231
rect 3985 26197 4019 26231
rect 4019 26197 4028 26231
rect 3976 26188 4028 26197
rect 4252 26367 4304 26376
rect 4252 26333 4261 26367
rect 4261 26333 4295 26367
rect 4295 26333 4304 26367
rect 4252 26324 4304 26333
rect 4712 26324 4764 26376
rect 4988 26324 5040 26376
rect 5356 26367 5408 26376
rect 4620 26256 4672 26308
rect 5080 26299 5132 26308
rect 5080 26265 5089 26299
rect 5089 26265 5123 26299
rect 5123 26265 5132 26299
rect 5080 26256 5132 26265
rect 5356 26333 5365 26367
rect 5365 26333 5399 26367
rect 5399 26333 5408 26367
rect 5356 26324 5408 26333
rect 8944 26324 8996 26376
rect 9588 26367 9640 26376
rect 9588 26333 9597 26367
rect 9597 26333 9631 26367
rect 9631 26333 9640 26367
rect 9588 26324 9640 26333
rect 10140 26324 10192 26376
rect 12072 26367 12124 26376
rect 12072 26333 12081 26367
rect 12081 26333 12115 26367
rect 12115 26333 12124 26367
rect 12072 26324 12124 26333
rect 12532 26528 12584 26580
rect 34336 26528 34388 26580
rect 20260 26460 20312 26512
rect 20536 26460 20588 26512
rect 14924 26435 14976 26444
rect 14924 26401 14933 26435
rect 14933 26401 14967 26435
rect 14967 26401 14976 26435
rect 14924 26392 14976 26401
rect 12440 26324 12492 26376
rect 13820 26324 13872 26376
rect 14372 26367 14424 26376
rect 14372 26333 14381 26367
rect 14381 26333 14415 26367
rect 14415 26333 14424 26367
rect 14372 26324 14424 26333
rect 16304 26367 16356 26376
rect 16304 26333 16313 26367
rect 16313 26333 16347 26367
rect 16347 26333 16356 26367
rect 16304 26324 16356 26333
rect 20352 26324 20404 26376
rect 20628 26392 20680 26444
rect 21364 26367 21416 26376
rect 21364 26333 21373 26367
rect 21373 26333 21407 26367
rect 21407 26333 21416 26367
rect 21364 26324 21416 26333
rect 21548 26367 21600 26376
rect 21548 26333 21557 26367
rect 21557 26333 21591 26367
rect 21591 26333 21600 26367
rect 21548 26324 21600 26333
rect 22376 26367 22428 26376
rect 22376 26333 22385 26367
rect 22385 26333 22419 26367
rect 22419 26333 22428 26367
rect 22376 26324 22428 26333
rect 22468 26367 22520 26376
rect 22468 26333 22477 26367
rect 22477 26333 22511 26367
rect 22511 26333 22520 26367
rect 23480 26392 23532 26444
rect 23756 26392 23808 26444
rect 22468 26324 22520 26333
rect 6920 26256 6972 26308
rect 9864 26256 9916 26308
rect 19984 26256 20036 26308
rect 4988 26188 5040 26240
rect 9496 26231 9548 26240
rect 9496 26197 9505 26231
rect 9505 26197 9539 26231
rect 9539 26197 9548 26231
rect 9496 26188 9548 26197
rect 10232 26231 10284 26240
rect 10232 26197 10241 26231
rect 10241 26197 10275 26231
rect 10275 26197 10284 26231
rect 10232 26188 10284 26197
rect 17592 26231 17644 26240
rect 17592 26197 17601 26231
rect 17601 26197 17635 26231
rect 17635 26197 17644 26231
rect 17592 26188 17644 26197
rect 20536 26194 20588 26246
rect 22008 26188 22060 26240
rect 24032 26324 24084 26376
rect 24216 26460 24268 26512
rect 27896 26460 27948 26512
rect 27988 26460 28040 26512
rect 32588 26503 32640 26512
rect 24860 26367 24912 26376
rect 24860 26333 24869 26367
rect 24869 26333 24903 26367
rect 24903 26333 24912 26367
rect 24860 26324 24912 26333
rect 28080 26392 28132 26444
rect 32588 26469 32597 26503
rect 32597 26469 32631 26503
rect 32631 26469 32640 26503
rect 32588 26460 32640 26469
rect 33416 26460 33468 26512
rect 26240 26324 26292 26376
rect 26608 26324 26660 26376
rect 33048 26392 33100 26444
rect 27528 26256 27580 26308
rect 31300 26231 31352 26240
rect 31300 26197 31309 26231
rect 31309 26197 31343 26231
rect 31343 26197 31352 26231
rect 31300 26188 31352 26197
rect 32864 26367 32916 26376
rect 32864 26333 32873 26367
rect 32873 26333 32907 26367
rect 32907 26333 32916 26367
rect 32864 26324 32916 26333
rect 31852 26256 31904 26308
rect 32680 26256 32732 26308
rect 32588 26188 32640 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4252 25984 4304 26036
rect 3148 25916 3200 25968
rect 5264 25916 5316 25968
rect 10784 25984 10836 26036
rect 12440 26027 12492 26036
rect 12440 25993 12449 26027
rect 12449 25993 12483 26027
rect 12483 25993 12492 26027
rect 12440 25984 12492 25993
rect 19340 25984 19392 26036
rect 20352 25984 20404 26036
rect 8944 25959 8996 25968
rect 8944 25925 8953 25959
rect 8953 25925 8987 25959
rect 8987 25925 8996 25959
rect 8944 25916 8996 25925
rect 3056 25823 3108 25832
rect 3056 25789 3065 25823
rect 3065 25789 3099 25823
rect 3099 25789 3108 25823
rect 3056 25780 3108 25789
rect 3976 25848 4028 25900
rect 5356 25891 5408 25900
rect 5356 25857 5365 25891
rect 5365 25857 5399 25891
rect 5399 25857 5408 25891
rect 5356 25848 5408 25857
rect 5724 25891 5776 25900
rect 5724 25857 5733 25891
rect 5733 25857 5767 25891
rect 5767 25857 5776 25891
rect 5724 25848 5776 25857
rect 5816 25891 5868 25900
rect 5816 25857 5825 25891
rect 5825 25857 5859 25891
rect 5859 25857 5868 25891
rect 5816 25848 5868 25857
rect 7104 25848 7156 25900
rect 7564 25848 7616 25900
rect 9864 25891 9916 25900
rect 5080 25780 5132 25832
rect 8576 25780 8628 25832
rect 9864 25857 9873 25891
rect 9873 25857 9907 25891
rect 9907 25857 9916 25891
rect 9864 25848 9916 25857
rect 10048 25891 10100 25900
rect 10048 25857 10057 25891
rect 10057 25857 10091 25891
rect 10091 25857 10100 25891
rect 10048 25848 10100 25857
rect 16028 25916 16080 25968
rect 17132 25916 17184 25968
rect 9496 25712 9548 25764
rect 10232 25780 10284 25832
rect 13820 25848 13872 25900
rect 15660 25891 15712 25900
rect 15660 25857 15669 25891
rect 15669 25857 15703 25891
rect 15703 25857 15712 25891
rect 15660 25848 15712 25857
rect 17868 25848 17920 25900
rect 24860 25848 24912 25900
rect 30932 25848 30984 25900
rect 31024 25891 31076 25900
rect 31024 25857 31033 25891
rect 31033 25857 31067 25891
rect 31067 25857 31076 25891
rect 31208 25891 31260 25900
rect 31024 25848 31076 25857
rect 31208 25857 31217 25891
rect 31217 25857 31251 25891
rect 31251 25857 31260 25891
rect 31208 25848 31260 25857
rect 32312 25848 32364 25900
rect 16948 25780 17000 25832
rect 21272 25780 21324 25832
rect 23572 25780 23624 25832
rect 4068 25644 4120 25696
rect 8300 25644 8352 25696
rect 9680 25644 9732 25696
rect 20260 25644 20312 25696
rect 29920 25687 29972 25696
rect 29920 25653 29929 25687
rect 29929 25653 29963 25687
rect 29963 25653 29972 25687
rect 29920 25644 29972 25653
rect 30840 25687 30892 25696
rect 30840 25653 30849 25687
rect 30849 25653 30883 25687
rect 30883 25653 30892 25687
rect 30840 25644 30892 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 4620 25440 4672 25492
rect 5080 25440 5132 25492
rect 7840 25440 7892 25492
rect 9588 25440 9640 25492
rect 10508 25440 10560 25492
rect 3516 25372 3568 25424
rect 4160 25372 4212 25424
rect 4988 25372 5040 25424
rect 5356 25304 5408 25356
rect 8576 25347 8628 25356
rect 4068 25236 4120 25288
rect 4712 25236 4764 25288
rect 4620 25168 4672 25220
rect 5172 25279 5224 25288
rect 5172 25245 5181 25279
rect 5181 25245 5215 25279
rect 5215 25245 5224 25279
rect 8576 25313 8585 25347
rect 8585 25313 8619 25347
rect 8619 25313 8628 25347
rect 8576 25304 8628 25313
rect 9680 25347 9732 25356
rect 9680 25313 9689 25347
rect 9689 25313 9723 25347
rect 9723 25313 9732 25347
rect 9680 25304 9732 25313
rect 5172 25236 5224 25245
rect 7840 25279 7892 25288
rect 7840 25245 7849 25279
rect 7849 25245 7883 25279
rect 7883 25245 7892 25279
rect 8300 25279 8352 25288
rect 7840 25236 7892 25245
rect 8300 25245 8309 25279
rect 8309 25245 8343 25279
rect 8343 25245 8352 25279
rect 8300 25236 8352 25245
rect 10048 25236 10100 25288
rect 10600 25279 10652 25288
rect 5264 25168 5316 25220
rect 4160 25100 4212 25152
rect 7748 25100 7800 25152
rect 9128 25143 9180 25152
rect 9128 25109 9137 25143
rect 9137 25109 9171 25143
rect 9171 25109 9180 25143
rect 9128 25100 9180 25109
rect 9680 25168 9732 25220
rect 10600 25245 10609 25279
rect 10609 25245 10643 25279
rect 10643 25245 10652 25279
rect 10600 25236 10652 25245
rect 10692 25236 10744 25288
rect 16488 25440 16540 25492
rect 16948 25483 17000 25492
rect 16948 25449 16957 25483
rect 16957 25449 16991 25483
rect 16991 25449 17000 25483
rect 16948 25440 17000 25449
rect 17868 25483 17920 25492
rect 17868 25449 17877 25483
rect 17877 25449 17911 25483
rect 17911 25449 17920 25483
rect 17868 25440 17920 25449
rect 14464 25372 14516 25424
rect 14648 25304 14700 25356
rect 16764 25304 16816 25356
rect 12624 25236 12676 25288
rect 13452 25279 13504 25288
rect 13452 25245 13461 25279
rect 13461 25245 13495 25279
rect 13495 25245 13504 25279
rect 13452 25236 13504 25245
rect 18052 25279 18104 25288
rect 18052 25245 18061 25279
rect 18061 25245 18095 25279
rect 18095 25245 18104 25279
rect 18052 25236 18104 25245
rect 18512 25236 18564 25288
rect 19248 25236 19300 25288
rect 20168 25304 20220 25356
rect 20628 25304 20680 25356
rect 23756 25304 23808 25356
rect 10784 25168 10836 25220
rect 12900 25168 12952 25220
rect 16580 25168 16632 25220
rect 17592 25168 17644 25220
rect 19340 25168 19392 25220
rect 20260 25236 20312 25288
rect 22284 25236 22336 25288
rect 29920 25236 29972 25288
rect 31300 25236 31352 25288
rect 31852 25440 31904 25492
rect 23480 25168 23532 25220
rect 23664 25168 23716 25220
rect 27620 25211 27672 25220
rect 27620 25177 27654 25211
rect 27654 25177 27672 25211
rect 27620 25168 27672 25177
rect 14648 25100 14700 25152
rect 20076 25100 20128 25152
rect 28724 25143 28776 25152
rect 28724 25109 28733 25143
rect 28733 25109 28767 25143
rect 28767 25109 28776 25143
rect 28724 25100 28776 25109
rect 32588 25143 32640 25152
rect 32588 25109 32597 25143
rect 32597 25109 32631 25143
rect 32631 25109 32640 25143
rect 32588 25100 32640 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 9864 24939 9916 24948
rect 9864 24905 9873 24939
rect 9873 24905 9907 24939
rect 9907 24905 9916 24939
rect 9864 24896 9916 24905
rect 10508 24939 10560 24948
rect 10508 24905 10517 24939
rect 10517 24905 10551 24939
rect 10551 24905 10560 24939
rect 10508 24896 10560 24905
rect 17132 24896 17184 24948
rect 3056 24828 3108 24880
rect 15660 24828 15712 24880
rect 16488 24828 16540 24880
rect 4712 24760 4764 24812
rect 7932 24760 7984 24812
rect 9128 24760 9180 24812
rect 5172 24556 5224 24608
rect 8208 24556 8260 24608
rect 9588 24692 9640 24744
rect 9128 24624 9180 24676
rect 12624 24760 12676 24812
rect 12900 24803 12952 24812
rect 12900 24769 12909 24803
rect 12909 24769 12943 24803
rect 12943 24769 12952 24803
rect 12900 24760 12952 24769
rect 13452 24760 13504 24812
rect 19340 24828 19392 24880
rect 20444 24828 20496 24880
rect 22284 24828 22336 24880
rect 24860 24896 24912 24948
rect 25780 24828 25832 24880
rect 32312 24828 32364 24880
rect 16856 24803 16908 24812
rect 16856 24769 16865 24803
rect 16865 24769 16899 24803
rect 16899 24769 16908 24803
rect 16856 24760 16908 24769
rect 17040 24803 17092 24812
rect 17040 24769 17049 24803
rect 17049 24769 17083 24803
rect 17083 24769 17092 24803
rect 17040 24760 17092 24769
rect 17224 24803 17276 24812
rect 17224 24769 17233 24803
rect 17233 24769 17267 24803
rect 17267 24769 17276 24803
rect 17224 24760 17276 24769
rect 18696 24760 18748 24812
rect 22376 24760 22428 24812
rect 22836 24803 22888 24812
rect 22836 24769 22845 24803
rect 22845 24769 22879 24803
rect 22879 24769 22888 24803
rect 22836 24760 22888 24769
rect 22928 24803 22980 24812
rect 22928 24769 22937 24803
rect 22937 24769 22971 24803
rect 22971 24769 22980 24803
rect 22928 24760 22980 24769
rect 24584 24760 24636 24812
rect 29736 24803 29788 24812
rect 29736 24769 29745 24803
rect 29745 24769 29779 24803
rect 29779 24769 29788 24803
rect 29736 24760 29788 24769
rect 32404 24760 32456 24812
rect 23664 24735 23716 24744
rect 23664 24701 23673 24735
rect 23673 24701 23707 24735
rect 23707 24701 23716 24735
rect 23664 24692 23716 24701
rect 27804 24692 27856 24744
rect 30932 24624 30984 24676
rect 9220 24599 9272 24608
rect 9220 24565 9229 24599
rect 9229 24565 9263 24599
rect 9263 24565 9272 24599
rect 9220 24556 9272 24565
rect 9588 24556 9640 24608
rect 23388 24556 23440 24608
rect 28908 24556 28960 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 16672 24352 16724 24404
rect 22836 24352 22888 24404
rect 24032 24395 24084 24404
rect 24032 24361 24041 24395
rect 24041 24361 24075 24395
rect 24075 24361 24084 24395
rect 24032 24352 24084 24361
rect 27620 24352 27672 24404
rect 31208 24352 31260 24404
rect 24860 24284 24912 24336
rect 29828 24284 29880 24336
rect 26424 24259 26476 24268
rect 26424 24225 26433 24259
rect 26433 24225 26467 24259
rect 26467 24225 26476 24259
rect 26424 24216 26476 24225
rect 27344 24216 27396 24268
rect 27620 24216 27672 24268
rect 15476 24191 15528 24200
rect 15476 24157 15485 24191
rect 15485 24157 15519 24191
rect 15519 24157 15528 24191
rect 15476 24148 15528 24157
rect 15752 24191 15804 24200
rect 15752 24157 15786 24191
rect 15786 24157 15804 24191
rect 22652 24191 22704 24200
rect 15752 24148 15804 24157
rect 22652 24157 22661 24191
rect 22661 24157 22695 24191
rect 22695 24157 22704 24191
rect 22652 24148 22704 24157
rect 24492 24148 24544 24200
rect 24676 24191 24728 24200
rect 24676 24157 24685 24191
rect 24685 24157 24719 24191
rect 24719 24157 24728 24191
rect 24676 24148 24728 24157
rect 25964 24148 26016 24200
rect 28080 24216 28132 24268
rect 20720 24080 20772 24132
rect 22192 24123 22244 24132
rect 22192 24089 22201 24123
rect 22201 24089 22235 24123
rect 22235 24089 22244 24123
rect 22192 24080 22244 24089
rect 22468 24080 22520 24132
rect 22744 24012 22796 24064
rect 27804 24148 27856 24200
rect 32496 24148 32548 24200
rect 26148 24080 26200 24132
rect 28724 24080 28776 24132
rect 30840 24080 30892 24132
rect 31760 24012 31812 24064
rect 32404 24012 32456 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 22468 23851 22520 23860
rect 22468 23817 22477 23851
rect 22477 23817 22511 23851
rect 22511 23817 22520 23851
rect 22468 23808 22520 23817
rect 23480 23808 23532 23860
rect 29736 23808 29788 23860
rect 14372 23740 14424 23792
rect 21364 23740 21416 23792
rect 12716 23715 12768 23724
rect 12716 23681 12725 23715
rect 12725 23681 12759 23715
rect 12759 23681 12768 23715
rect 12716 23672 12768 23681
rect 20260 23672 20312 23724
rect 20536 23672 20588 23724
rect 14188 23604 14240 23656
rect 19800 23604 19852 23656
rect 22744 23604 22796 23656
rect 24676 23740 24728 23792
rect 22928 23715 22980 23724
rect 22928 23681 22934 23715
rect 22934 23681 22968 23715
rect 22968 23681 22980 23715
rect 22928 23672 22980 23681
rect 25228 23672 25280 23724
rect 26424 23672 26476 23724
rect 27436 23672 27488 23724
rect 26240 23604 26292 23656
rect 32956 23604 33008 23656
rect 35992 23715 36044 23724
rect 35992 23681 36001 23715
rect 36001 23681 36035 23715
rect 36035 23681 36044 23715
rect 35992 23672 36044 23681
rect 34612 23604 34664 23656
rect 17040 23536 17092 23588
rect 20536 23536 20588 23588
rect 8024 23468 8076 23520
rect 19984 23468 20036 23520
rect 36084 23468 36136 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 4160 23264 4212 23316
rect 4620 23264 4672 23316
rect 7840 23264 7892 23316
rect 14372 23307 14424 23316
rect 14372 23273 14381 23307
rect 14381 23273 14415 23307
rect 14415 23273 14424 23307
rect 14372 23264 14424 23273
rect 20352 23264 20404 23316
rect 20628 23264 20680 23316
rect 4712 23196 4764 23248
rect 4804 23196 4856 23248
rect 11888 23196 11940 23248
rect 3608 23128 3660 23180
rect 3240 23060 3292 23112
rect 10968 23128 11020 23180
rect 17776 23196 17828 23248
rect 20168 23196 20220 23248
rect 19800 23128 19852 23180
rect 20076 23171 20128 23180
rect 20076 23137 20085 23171
rect 20085 23137 20119 23171
rect 20119 23137 20128 23171
rect 23664 23264 23716 23316
rect 25228 23264 25280 23316
rect 26056 23264 26108 23316
rect 32496 23307 32548 23316
rect 32496 23273 32505 23307
rect 32505 23273 32539 23307
rect 32539 23273 32548 23307
rect 32496 23264 32548 23273
rect 25964 23239 26016 23248
rect 25964 23205 25973 23239
rect 25973 23205 26007 23239
rect 26007 23205 26016 23239
rect 25964 23196 26016 23205
rect 20076 23128 20128 23137
rect 22928 23128 22980 23180
rect 36176 23196 36228 23248
rect 4160 23035 4212 23044
rect 4160 23001 4169 23035
rect 4169 23001 4203 23035
rect 4203 23001 4212 23035
rect 4160 22992 4212 23001
rect 5356 23060 5408 23112
rect 12992 23103 13044 23112
rect 12992 23069 13001 23103
rect 13001 23069 13035 23103
rect 13035 23069 13044 23103
rect 12992 23060 13044 23069
rect 13176 23103 13228 23112
rect 13176 23069 13185 23103
rect 13185 23069 13219 23103
rect 13219 23069 13228 23103
rect 13176 23060 13228 23069
rect 14280 23103 14332 23112
rect 7656 23035 7708 23044
rect 7656 23001 7665 23035
rect 7665 23001 7699 23035
rect 7699 23001 7708 23035
rect 7656 22992 7708 23001
rect 7932 23035 7984 23044
rect 7932 23001 7941 23035
rect 7941 23001 7975 23035
rect 7975 23001 7984 23035
rect 7932 22992 7984 23001
rect 12808 22992 12860 23044
rect 14280 23069 14289 23103
rect 14289 23069 14323 23103
rect 14323 23069 14332 23103
rect 14280 23060 14332 23069
rect 14372 23060 14424 23112
rect 14556 23060 14608 23112
rect 19340 23060 19392 23112
rect 14188 22992 14240 23044
rect 15844 22992 15896 23044
rect 17592 22992 17644 23044
rect 20628 23060 20680 23112
rect 20996 23103 21048 23112
rect 20996 23069 21005 23103
rect 21005 23069 21039 23103
rect 21039 23069 21048 23103
rect 20996 23060 21048 23069
rect 22192 23060 22244 23112
rect 23572 23103 23624 23112
rect 4344 22967 4396 22976
rect 4344 22933 4353 22967
rect 4353 22933 4387 22967
rect 4387 22933 4396 22967
rect 4344 22924 4396 22933
rect 7564 22924 7616 22976
rect 7748 22924 7800 22976
rect 19984 22967 20036 22976
rect 19984 22933 19993 22967
rect 19993 22933 20027 22967
rect 20027 22933 20036 22967
rect 19984 22924 20036 22933
rect 22560 22924 22612 22976
rect 23572 23069 23581 23103
rect 23581 23069 23615 23103
rect 23615 23069 23624 23103
rect 23572 23060 23624 23069
rect 35992 23128 36044 23180
rect 24032 23060 24084 23112
rect 24584 23103 24636 23112
rect 24584 23069 24593 23103
rect 24593 23069 24627 23103
rect 24627 23069 24636 23103
rect 24584 23060 24636 23069
rect 30932 23060 30984 23112
rect 36360 23060 36412 23112
rect 25872 22992 25924 23044
rect 26516 23035 26568 23044
rect 26516 23001 26525 23035
rect 26525 23001 26559 23035
rect 26559 23001 26568 23035
rect 26516 22992 26568 23001
rect 26148 22924 26200 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 2964 22720 3016 22772
rect 4344 22720 4396 22772
rect 7656 22720 7708 22772
rect 8300 22720 8352 22772
rect 8392 22720 8444 22772
rect 11888 22720 11940 22772
rect 14372 22720 14424 22772
rect 16856 22720 16908 22772
rect 3516 22695 3568 22704
rect 3516 22661 3525 22695
rect 3525 22661 3559 22695
rect 3559 22661 3568 22695
rect 3516 22652 3568 22661
rect 8024 22695 8076 22704
rect 8024 22661 8033 22695
rect 8033 22661 8067 22695
rect 8067 22661 8076 22695
rect 8024 22652 8076 22661
rect 4620 22584 4672 22636
rect 5724 22584 5776 22636
rect 7012 22627 7064 22636
rect 7012 22593 7021 22627
rect 7021 22593 7055 22627
rect 7055 22593 7064 22627
rect 7012 22584 7064 22593
rect 7380 22627 7432 22636
rect 7380 22593 7389 22627
rect 7389 22593 7423 22627
rect 7423 22593 7432 22627
rect 7380 22584 7432 22593
rect 8208 22627 8260 22636
rect 8208 22593 8214 22627
rect 8214 22593 8260 22627
rect 8208 22584 8260 22593
rect 14280 22652 14332 22704
rect 15476 22652 15528 22704
rect 17592 22695 17644 22704
rect 17592 22661 17601 22695
rect 17601 22661 17635 22695
rect 17635 22661 17644 22695
rect 17592 22652 17644 22661
rect 18880 22652 18932 22704
rect 19984 22652 20036 22704
rect 3608 22516 3660 22568
rect 8392 22559 8444 22568
rect 8392 22525 8401 22559
rect 8401 22525 8435 22559
rect 8435 22525 8444 22559
rect 8392 22516 8444 22525
rect 9588 22516 9640 22568
rect 7104 22448 7156 22500
rect 11888 22627 11940 22636
rect 11888 22593 11897 22627
rect 11897 22593 11931 22627
rect 11931 22593 11940 22627
rect 11888 22584 11940 22593
rect 16580 22584 16632 22636
rect 19064 22627 19116 22636
rect 19064 22593 19073 22627
rect 19073 22593 19107 22627
rect 19107 22593 19116 22627
rect 19064 22584 19116 22593
rect 20628 22720 20680 22772
rect 25872 22763 25924 22772
rect 25872 22729 25881 22763
rect 25881 22729 25915 22763
rect 25915 22729 25924 22763
rect 25872 22720 25924 22729
rect 26240 22763 26292 22772
rect 26240 22729 26249 22763
rect 26249 22729 26283 22763
rect 26283 22729 26292 22763
rect 26240 22720 26292 22729
rect 27528 22720 27580 22772
rect 36360 22763 36412 22772
rect 36360 22729 36369 22763
rect 36369 22729 36403 22763
rect 36403 22729 36412 22763
rect 36360 22720 36412 22729
rect 21088 22652 21140 22704
rect 20444 22627 20496 22636
rect 20444 22593 20453 22627
rect 20453 22593 20487 22627
rect 20487 22593 20496 22627
rect 20444 22584 20496 22593
rect 24860 22584 24912 22636
rect 25780 22584 25832 22636
rect 31024 22652 31076 22704
rect 26332 22627 26384 22636
rect 26332 22593 26341 22627
rect 26341 22593 26375 22627
rect 26375 22593 26384 22627
rect 26332 22584 26384 22593
rect 27620 22584 27672 22636
rect 12072 22559 12124 22568
rect 12072 22525 12081 22559
rect 12081 22525 12115 22559
rect 12115 22525 12124 22559
rect 12072 22516 12124 22525
rect 27896 22584 27948 22636
rect 28172 22627 28224 22636
rect 28172 22593 28181 22627
rect 28181 22593 28215 22627
rect 28215 22593 28224 22627
rect 29920 22627 29972 22636
rect 28172 22584 28224 22593
rect 29920 22593 29929 22627
rect 29929 22593 29963 22627
rect 29963 22593 29972 22627
rect 29920 22584 29972 22593
rect 30932 22584 30984 22636
rect 33324 22627 33376 22636
rect 33324 22593 33333 22627
rect 33333 22593 33367 22627
rect 33367 22593 33376 22627
rect 33324 22584 33376 22593
rect 33416 22627 33468 22636
rect 33416 22593 33425 22627
rect 33425 22593 33459 22627
rect 33459 22593 33468 22627
rect 33416 22584 33468 22593
rect 18880 22448 18932 22500
rect 29552 22516 29604 22568
rect 36084 22584 36136 22636
rect 36268 22627 36320 22636
rect 36268 22593 36277 22627
rect 36277 22593 36311 22627
rect 36311 22593 36320 22627
rect 36268 22584 36320 22593
rect 27988 22448 28040 22500
rect 30748 22448 30800 22500
rect 35900 22516 35952 22568
rect 35992 22448 36044 22500
rect 7748 22380 7800 22432
rect 8576 22380 8628 22432
rect 9772 22423 9824 22432
rect 9772 22389 9781 22423
rect 9781 22389 9815 22423
rect 9815 22389 9824 22423
rect 9772 22380 9824 22389
rect 12992 22380 13044 22432
rect 14004 22380 14056 22432
rect 17960 22423 18012 22432
rect 17960 22389 17969 22423
rect 17969 22389 18003 22423
rect 18003 22389 18012 22423
rect 17960 22380 18012 22389
rect 18788 22423 18840 22432
rect 18788 22389 18797 22423
rect 18797 22389 18831 22423
rect 18831 22389 18840 22423
rect 18788 22380 18840 22389
rect 19984 22423 20036 22432
rect 19984 22389 19993 22423
rect 19993 22389 20027 22423
rect 20027 22389 20036 22423
rect 19984 22380 20036 22389
rect 24768 22380 24820 22432
rect 27620 22380 27672 22432
rect 34520 22380 34572 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3240 22219 3292 22228
rect 3240 22185 3249 22219
rect 3249 22185 3283 22219
rect 3283 22185 3292 22219
rect 3240 22176 3292 22185
rect 3608 22176 3660 22228
rect 7932 22176 7984 22228
rect 7564 22108 7616 22160
rect 4620 22040 4672 22092
rect 8392 22108 8444 22160
rect 9772 22108 9824 22160
rect 12716 22176 12768 22228
rect 16212 22176 16264 22228
rect 19064 22176 19116 22228
rect 8576 22040 8628 22092
rect 2964 21904 3016 21956
rect 4436 21972 4488 22024
rect 4804 21972 4856 22024
rect 4252 21904 4304 21956
rect 1860 21836 1912 21888
rect 7288 22015 7340 22024
rect 7288 21981 7297 22015
rect 7297 21981 7331 22015
rect 7331 21981 7340 22015
rect 7288 21972 7340 21981
rect 8300 22015 8352 22024
rect 8300 21981 8309 22015
rect 8309 21981 8343 22015
rect 8343 21981 8352 22015
rect 8300 21972 8352 21981
rect 8484 22015 8536 22024
rect 8484 21981 8493 22015
rect 8493 21981 8527 22015
rect 8527 21981 8536 22015
rect 8484 21972 8536 21981
rect 9312 22015 9364 22024
rect 9312 21981 9321 22015
rect 9321 21981 9355 22015
rect 9355 21981 9364 22015
rect 9312 21972 9364 21981
rect 16856 22108 16908 22160
rect 24860 22151 24912 22160
rect 24860 22117 24869 22151
rect 24869 22117 24903 22151
rect 24903 22117 24912 22151
rect 24860 22108 24912 22117
rect 26516 22176 26568 22228
rect 27804 22219 27856 22228
rect 27804 22185 27813 22219
rect 27813 22185 27847 22219
rect 27847 22185 27856 22219
rect 27804 22176 27856 22185
rect 29920 22176 29972 22228
rect 33324 22176 33376 22228
rect 34612 22108 34664 22160
rect 10968 22083 11020 22092
rect 7472 21904 7524 21956
rect 8024 21904 8076 21956
rect 10968 22049 10977 22083
rect 10977 22049 11011 22083
rect 11011 22049 11020 22083
rect 10968 22040 11020 22049
rect 9680 22015 9732 22024
rect 9680 21981 9689 22015
rect 9689 21981 9723 22015
rect 9723 21981 9732 22015
rect 9680 21972 9732 21981
rect 12072 21972 12124 22024
rect 14372 22015 14424 22024
rect 14372 21981 14381 22015
rect 14381 21981 14415 22015
rect 14415 21981 14424 22015
rect 14372 21972 14424 21981
rect 15568 21972 15620 22024
rect 16672 22040 16724 22092
rect 16212 22015 16264 22024
rect 16212 21981 16221 22015
rect 16221 21981 16255 22015
rect 16255 21981 16264 22015
rect 16212 21972 16264 21981
rect 16304 21972 16356 22024
rect 19340 22040 19392 22092
rect 26608 22040 26660 22092
rect 27712 22083 27764 22092
rect 27712 22049 27721 22083
rect 27721 22049 27755 22083
rect 27755 22049 27764 22083
rect 27712 22040 27764 22049
rect 29552 22040 29604 22092
rect 32956 22083 33008 22092
rect 19432 22015 19484 22024
rect 14832 21947 14884 21956
rect 14832 21913 14841 21947
rect 14841 21913 14875 21947
rect 14875 21913 14884 21947
rect 14832 21904 14884 21913
rect 16580 21904 16632 21956
rect 16948 21904 17000 21956
rect 6920 21836 6972 21888
rect 8208 21836 8260 21888
rect 9772 21836 9824 21888
rect 9864 21836 9916 21888
rect 19432 21981 19441 22015
rect 19441 21981 19475 22015
rect 19475 21981 19484 22015
rect 19432 21972 19484 21981
rect 19984 21972 20036 22024
rect 20260 21972 20312 22024
rect 24676 21972 24728 22024
rect 26240 22015 26292 22024
rect 26240 21981 26249 22015
rect 26249 21981 26283 22015
rect 26283 21981 26292 22015
rect 26240 21972 26292 21981
rect 27620 22015 27672 22024
rect 17592 21904 17644 21956
rect 18328 21836 18380 21888
rect 21916 21904 21968 21956
rect 27620 21981 27629 22015
rect 27629 21981 27663 22015
rect 27663 21981 27672 22015
rect 27620 21972 27672 21981
rect 30748 22015 30800 22024
rect 28080 21904 28132 21956
rect 28908 21904 28960 21956
rect 30748 21981 30757 22015
rect 30757 21981 30791 22015
rect 30791 21981 30800 22015
rect 30748 21972 30800 21981
rect 30932 22015 30984 22024
rect 30932 21981 30941 22015
rect 30941 21981 30975 22015
rect 30975 21981 30984 22015
rect 30932 21972 30984 21981
rect 32956 22049 32965 22083
rect 32965 22049 32999 22083
rect 32999 22049 33008 22083
rect 32956 22040 33008 22049
rect 33416 21972 33468 22024
rect 34520 21972 34572 22024
rect 35348 21904 35400 21956
rect 37188 21972 37240 22024
rect 38016 22015 38068 22024
rect 38016 21981 38025 22015
rect 38025 21981 38059 22015
rect 38059 21981 38068 22015
rect 38016 21972 38068 21981
rect 36728 21904 36780 21956
rect 21088 21836 21140 21888
rect 21364 21836 21416 21888
rect 21456 21836 21508 21888
rect 35072 21879 35124 21888
rect 35072 21845 35081 21879
rect 35081 21845 35115 21879
rect 35115 21845 35124 21879
rect 35072 21836 35124 21845
rect 37188 21836 37240 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 7012 21632 7064 21684
rect 7380 21632 7432 21684
rect 9312 21632 9364 21684
rect 14372 21632 14424 21684
rect 20720 21632 20772 21684
rect 20812 21632 20864 21684
rect 21456 21632 21508 21684
rect 24492 21675 24544 21684
rect 24492 21641 24501 21675
rect 24501 21641 24535 21675
rect 24535 21641 24544 21675
rect 24492 21632 24544 21641
rect 1860 21539 1912 21548
rect 1860 21505 1869 21539
rect 1869 21505 1903 21539
rect 1903 21505 1912 21539
rect 1860 21496 1912 21505
rect 4252 21539 4304 21548
rect 4252 21505 4261 21539
rect 4261 21505 4295 21539
rect 4295 21505 4304 21539
rect 4252 21496 4304 21505
rect 4436 21539 4488 21548
rect 4436 21505 4445 21539
rect 4445 21505 4479 21539
rect 4479 21505 4488 21539
rect 4436 21496 4488 21505
rect 5080 21496 5132 21548
rect 7748 21564 7800 21616
rect 8116 21564 8168 21616
rect 9864 21564 9916 21616
rect 15660 21564 15712 21616
rect 7472 21539 7524 21548
rect 7472 21505 7481 21539
rect 7481 21505 7515 21539
rect 7515 21505 7524 21539
rect 7472 21496 7524 21505
rect 7564 21496 7616 21548
rect 9128 21496 9180 21548
rect 10232 21496 10284 21548
rect 10692 21496 10744 21548
rect 10876 21539 10928 21548
rect 10876 21505 10885 21539
rect 10885 21505 10919 21539
rect 10919 21505 10928 21539
rect 10876 21496 10928 21505
rect 12072 21539 12124 21548
rect 2780 21428 2832 21480
rect 4804 21428 4856 21480
rect 5448 21428 5500 21480
rect 7288 21428 7340 21480
rect 9404 21471 9456 21480
rect 9404 21437 9413 21471
rect 9413 21437 9447 21471
rect 9447 21437 9456 21471
rect 9404 21428 9456 21437
rect 12072 21505 12081 21539
rect 12081 21505 12115 21539
rect 12115 21505 12124 21539
rect 12072 21496 12124 21505
rect 14004 21496 14056 21548
rect 14832 21496 14884 21548
rect 16028 21539 16080 21548
rect 16028 21505 16037 21539
rect 16037 21505 16071 21539
rect 16071 21505 16080 21539
rect 16028 21496 16080 21505
rect 16580 21564 16632 21616
rect 17224 21564 17276 21616
rect 17960 21564 18012 21616
rect 20444 21564 20496 21616
rect 23388 21607 23440 21616
rect 16488 21496 16540 21548
rect 21272 21539 21324 21548
rect 12532 21428 12584 21480
rect 13176 21428 13228 21480
rect 20812 21428 20864 21480
rect 21272 21505 21281 21539
rect 21281 21505 21315 21539
rect 21315 21505 21324 21539
rect 21272 21496 21324 21505
rect 23388 21573 23422 21607
rect 23422 21573 23440 21607
rect 23388 21564 23440 21573
rect 21548 21496 21600 21548
rect 27988 21539 28040 21548
rect 27988 21505 27997 21539
rect 27997 21505 28031 21539
rect 28031 21505 28040 21539
rect 27988 21496 28040 21505
rect 28172 21539 28224 21548
rect 28172 21505 28181 21539
rect 28181 21505 28215 21539
rect 28215 21505 28224 21539
rect 28172 21496 28224 21505
rect 35072 21632 35124 21684
rect 36636 21564 36688 21616
rect 38016 21564 38068 21616
rect 35900 21496 35952 21548
rect 14924 21360 14976 21412
rect 22376 21428 22428 21480
rect 22560 21428 22612 21480
rect 29736 21428 29788 21480
rect 34520 21428 34572 21480
rect 34796 21428 34848 21480
rect 35348 21428 35400 21480
rect 35808 21428 35860 21480
rect 36176 21428 36228 21480
rect 2872 21292 2924 21344
rect 3148 21292 3200 21344
rect 8300 21292 8352 21344
rect 9220 21335 9272 21344
rect 9220 21301 9229 21335
rect 9229 21301 9263 21335
rect 9263 21301 9272 21335
rect 9220 21292 9272 21301
rect 11980 21292 12032 21344
rect 13176 21292 13228 21344
rect 16120 21292 16172 21344
rect 16212 21292 16264 21344
rect 18052 21292 18104 21344
rect 19340 21292 19392 21344
rect 20904 21335 20956 21344
rect 20904 21301 20913 21335
rect 20913 21301 20947 21335
rect 20947 21301 20956 21335
rect 20904 21292 20956 21301
rect 29828 21292 29880 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 6920 21088 6972 21140
rect 10876 21088 10928 21140
rect 12072 21088 12124 21140
rect 23664 21088 23716 21140
rect 24584 21088 24636 21140
rect 36084 21088 36136 21140
rect 4620 21020 4672 21072
rect 35348 21063 35400 21072
rect 35348 21029 35357 21063
rect 35357 21029 35391 21063
rect 35391 21029 35400 21063
rect 35348 21020 35400 21029
rect 7104 20952 7156 21004
rect 2780 20927 2832 20936
rect 2780 20893 2789 20927
rect 2789 20893 2823 20927
rect 2823 20893 2832 20927
rect 7472 20952 7524 21004
rect 2780 20884 2832 20893
rect 7564 20927 7616 20936
rect 2964 20816 3016 20868
rect 7564 20893 7573 20927
rect 7573 20893 7607 20927
rect 7607 20893 7616 20927
rect 7564 20884 7616 20893
rect 9864 20952 9916 21004
rect 12440 20952 12492 21004
rect 13452 20952 13504 21004
rect 14556 20952 14608 21004
rect 14924 20995 14976 21004
rect 14924 20961 14933 20995
rect 14933 20961 14967 20995
rect 14967 20961 14976 20995
rect 14924 20952 14976 20961
rect 17592 20952 17644 21004
rect 22560 20995 22612 21004
rect 22560 20961 22569 20995
rect 22569 20961 22603 20995
rect 22603 20961 22612 20995
rect 22560 20952 22612 20961
rect 28908 20952 28960 21004
rect 9772 20927 9824 20936
rect 9772 20893 9781 20927
rect 9781 20893 9815 20927
rect 9815 20893 9824 20927
rect 9772 20884 9824 20893
rect 11980 20927 12032 20936
rect 5448 20816 5500 20868
rect 7012 20816 7064 20868
rect 9036 20816 9088 20868
rect 11980 20893 11989 20927
rect 11989 20893 12023 20927
rect 12023 20893 12032 20927
rect 11980 20884 12032 20893
rect 13912 20884 13964 20936
rect 14464 20884 14516 20936
rect 24768 20884 24820 20936
rect 29828 20884 29880 20936
rect 34796 20952 34848 21004
rect 35808 20952 35860 21004
rect 36636 20995 36688 21004
rect 36176 20927 36228 20936
rect 36176 20893 36199 20927
rect 36199 20893 36228 20927
rect 5264 20748 5316 20800
rect 9404 20748 9456 20800
rect 16488 20816 16540 20868
rect 36176 20884 36228 20893
rect 36636 20961 36645 20995
rect 36645 20961 36679 20995
rect 36679 20961 36688 20995
rect 36636 20952 36688 20961
rect 35900 20816 35952 20868
rect 36728 20816 36780 20868
rect 10416 20791 10468 20800
rect 10416 20757 10425 20791
rect 10425 20757 10459 20791
rect 10459 20757 10468 20791
rect 10416 20748 10468 20757
rect 29000 20748 29052 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 2780 20587 2832 20596
rect 2780 20553 2789 20587
rect 2789 20553 2823 20587
rect 2823 20553 2832 20587
rect 2780 20544 2832 20553
rect 6920 20587 6972 20596
rect 6920 20553 6938 20587
rect 6938 20553 6972 20587
rect 6920 20544 6972 20553
rect 12072 20544 12124 20596
rect 16948 20544 17000 20596
rect 18328 20544 18380 20596
rect 19432 20544 19484 20596
rect 20996 20544 21048 20596
rect 7564 20476 7616 20528
rect 19340 20476 19392 20528
rect 20812 20519 20864 20528
rect 20812 20485 20821 20519
rect 20821 20485 20855 20519
rect 20855 20485 20864 20519
rect 20812 20476 20864 20485
rect 21272 20476 21324 20528
rect 21640 20476 21692 20528
rect 26608 20476 26660 20528
rect 29552 20476 29604 20528
rect 2872 20408 2924 20460
rect 4712 20408 4764 20460
rect 7380 20408 7432 20460
rect 9036 20451 9088 20460
rect 9036 20417 9045 20451
rect 9045 20417 9079 20451
rect 9079 20417 9088 20451
rect 9036 20408 9088 20417
rect 9680 20408 9732 20460
rect 12440 20408 12492 20460
rect 14832 20408 14884 20460
rect 15568 20451 15620 20460
rect 15568 20417 15577 20451
rect 15577 20417 15611 20451
rect 15611 20417 15620 20451
rect 15568 20408 15620 20417
rect 15660 20451 15712 20460
rect 15660 20417 15669 20451
rect 15669 20417 15703 20451
rect 15703 20417 15712 20451
rect 15660 20408 15712 20417
rect 8208 20272 8260 20324
rect 12532 20340 12584 20392
rect 13636 20340 13688 20392
rect 16304 20340 16356 20392
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 20168 20408 20220 20460
rect 20536 20451 20588 20460
rect 20536 20417 20546 20451
rect 20546 20417 20580 20451
rect 20580 20417 20588 20451
rect 20720 20451 20772 20460
rect 20536 20408 20588 20417
rect 20720 20417 20729 20451
rect 20729 20417 20763 20451
rect 20763 20417 20772 20451
rect 20720 20408 20772 20417
rect 21456 20408 21508 20460
rect 23388 20408 23440 20460
rect 16856 20272 16908 20324
rect 7472 20204 7524 20256
rect 7748 20247 7800 20256
rect 7748 20213 7757 20247
rect 7757 20213 7791 20247
rect 7791 20213 7800 20247
rect 7748 20204 7800 20213
rect 13820 20204 13872 20256
rect 18052 20204 18104 20256
rect 23572 20204 23624 20256
rect 25964 20408 26016 20460
rect 26332 20451 26384 20460
rect 26332 20417 26341 20451
rect 26341 20417 26375 20451
rect 26375 20417 26384 20451
rect 26332 20408 26384 20417
rect 27620 20408 27672 20460
rect 24032 20383 24084 20392
rect 24032 20349 24041 20383
rect 24041 20349 24075 20383
rect 24075 20349 24084 20383
rect 24032 20340 24084 20349
rect 23756 20272 23808 20324
rect 29552 20272 29604 20324
rect 30748 20451 30800 20460
rect 30748 20417 30757 20451
rect 30757 20417 30791 20451
rect 30791 20417 30800 20451
rect 30748 20408 30800 20417
rect 31760 20476 31812 20528
rect 31116 20340 31168 20392
rect 32312 20340 32364 20392
rect 38108 20383 38160 20392
rect 38108 20349 38117 20383
rect 38117 20349 38151 20383
rect 38151 20349 38160 20383
rect 38108 20340 38160 20349
rect 25872 20247 25924 20256
rect 25872 20213 25881 20247
rect 25881 20213 25915 20247
rect 25915 20213 25924 20247
rect 25872 20204 25924 20213
rect 30012 20204 30064 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 17224 20043 17276 20052
rect 17224 20009 17233 20043
rect 17233 20009 17267 20043
rect 17267 20009 17276 20043
rect 17224 20000 17276 20009
rect 20536 20000 20588 20052
rect 20812 20043 20864 20052
rect 20812 20009 20821 20043
rect 20821 20009 20855 20043
rect 20855 20009 20864 20043
rect 20812 20000 20864 20009
rect 22008 20000 22060 20052
rect 12900 19796 12952 19848
rect 13176 19796 13228 19848
rect 14556 19796 14608 19848
rect 19432 19907 19484 19916
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 24860 20000 24912 20052
rect 22192 19932 22244 19984
rect 13636 19660 13688 19712
rect 15660 19796 15712 19848
rect 16120 19839 16172 19848
rect 16120 19805 16154 19839
rect 16154 19805 16172 19839
rect 16120 19796 16172 19805
rect 20904 19796 20956 19848
rect 21272 19839 21324 19848
rect 21272 19805 21281 19839
rect 21281 19805 21315 19839
rect 21315 19805 21324 19839
rect 21272 19796 21324 19805
rect 21364 19839 21416 19848
rect 21364 19805 21374 19839
rect 21374 19805 21408 19839
rect 21408 19805 21416 19839
rect 21640 19839 21692 19848
rect 21364 19796 21416 19805
rect 21640 19805 21649 19839
rect 21649 19805 21683 19839
rect 21683 19805 21692 19839
rect 21640 19796 21692 19805
rect 22468 19864 22520 19916
rect 23664 19839 23716 19848
rect 23664 19805 23673 19839
rect 23673 19805 23707 19839
rect 23707 19805 23716 19839
rect 23664 19796 23716 19805
rect 28172 20000 28224 20052
rect 28356 20043 28408 20052
rect 28356 20009 28365 20043
rect 28365 20009 28399 20043
rect 28399 20009 28408 20043
rect 28356 20000 28408 20009
rect 28632 20043 28684 20052
rect 28632 20009 28641 20043
rect 28641 20009 28675 20043
rect 28675 20009 28684 20043
rect 28632 20000 28684 20009
rect 30748 20000 30800 20052
rect 33324 20000 33376 20052
rect 34796 20000 34848 20052
rect 36268 20000 36320 20052
rect 30012 19907 30064 19916
rect 30012 19873 30021 19907
rect 30021 19873 30055 19907
rect 30055 19873 30064 19907
rect 30012 19864 30064 19873
rect 33324 19864 33376 19916
rect 26056 19839 26108 19848
rect 17040 19728 17092 19780
rect 21180 19728 21232 19780
rect 21456 19728 21508 19780
rect 23848 19728 23900 19780
rect 26056 19805 26065 19839
rect 26065 19805 26099 19839
rect 26099 19805 26108 19839
rect 26056 19796 26108 19805
rect 28264 19839 28316 19848
rect 28264 19805 28273 19839
rect 28273 19805 28307 19839
rect 28307 19805 28316 19839
rect 28264 19796 28316 19805
rect 29000 19796 29052 19848
rect 29644 19796 29696 19848
rect 32312 19839 32364 19848
rect 26884 19728 26936 19780
rect 32312 19805 32321 19839
rect 32321 19805 32355 19839
rect 32355 19805 32364 19839
rect 32312 19796 32364 19805
rect 36176 19864 36228 19916
rect 32496 19728 32548 19780
rect 35348 19796 35400 19848
rect 35992 19839 36044 19848
rect 35992 19805 36001 19839
rect 36001 19805 36035 19839
rect 36035 19805 36044 19839
rect 35992 19796 36044 19805
rect 36544 19839 36596 19848
rect 36544 19805 36553 19839
rect 36553 19805 36587 19839
rect 36587 19805 36596 19839
rect 36544 19796 36596 19805
rect 36912 19796 36964 19848
rect 36452 19728 36504 19780
rect 16304 19660 16356 19712
rect 22928 19660 22980 19712
rect 23388 19660 23440 19712
rect 27528 19660 27580 19712
rect 31208 19660 31260 19712
rect 32220 19703 32272 19712
rect 32220 19669 32229 19703
rect 32229 19669 32263 19703
rect 32263 19669 32272 19703
rect 32220 19660 32272 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 7104 19456 7156 19508
rect 14004 19499 14056 19508
rect 14004 19465 14013 19499
rect 14013 19465 14047 19499
rect 14047 19465 14056 19499
rect 14004 19456 14056 19465
rect 22100 19456 22152 19508
rect 23848 19499 23900 19508
rect 23848 19465 23857 19499
rect 23857 19465 23891 19499
rect 23891 19465 23900 19499
rect 23848 19456 23900 19465
rect 26608 19499 26660 19508
rect 26608 19465 26617 19499
rect 26617 19465 26651 19499
rect 26651 19465 26660 19499
rect 26608 19456 26660 19465
rect 35900 19456 35952 19508
rect 4804 19363 4856 19372
rect 4804 19329 4813 19363
rect 4813 19329 4847 19363
rect 4847 19329 4856 19363
rect 4804 19320 4856 19329
rect 5080 19363 5132 19372
rect 5080 19329 5089 19363
rect 5089 19329 5123 19363
rect 5123 19329 5132 19363
rect 5080 19320 5132 19329
rect 6736 19363 6788 19372
rect 6736 19329 6745 19363
rect 6745 19329 6779 19363
rect 6779 19329 6788 19363
rect 6736 19320 6788 19329
rect 6920 19320 6972 19372
rect 25872 19388 25924 19440
rect 26884 19388 26936 19440
rect 32220 19388 32272 19440
rect 8944 19320 8996 19372
rect 13452 19320 13504 19372
rect 14556 19320 14608 19372
rect 15384 19320 15436 19372
rect 18788 19320 18840 19372
rect 22008 19320 22060 19372
rect 23204 19320 23256 19372
rect 7012 19295 7064 19304
rect 7012 19261 7021 19295
rect 7021 19261 7055 19295
rect 7055 19261 7064 19295
rect 7012 19252 7064 19261
rect 15200 19252 15252 19304
rect 25228 19295 25280 19304
rect 25228 19261 25237 19295
rect 25237 19261 25271 19295
rect 25271 19261 25280 19295
rect 25228 19252 25280 19261
rect 4896 19159 4948 19168
rect 4896 19125 4905 19159
rect 4905 19125 4939 19159
rect 4939 19125 4948 19159
rect 4896 19116 4948 19125
rect 6092 19116 6144 19168
rect 7748 19116 7800 19168
rect 18144 19159 18196 19168
rect 18144 19125 18153 19159
rect 18153 19125 18187 19159
rect 18187 19125 18196 19159
rect 18144 19116 18196 19125
rect 25872 19116 25924 19168
rect 27620 19363 27672 19372
rect 27620 19329 27629 19363
rect 27629 19329 27663 19363
rect 27663 19329 27672 19363
rect 27620 19320 27672 19329
rect 36176 19363 36228 19372
rect 36176 19329 36185 19363
rect 36185 19329 36219 19363
rect 36219 19329 36228 19363
rect 36176 19320 36228 19329
rect 36912 19320 36964 19372
rect 29644 19295 29696 19304
rect 29644 19261 29653 19295
rect 29653 19261 29687 19295
rect 29687 19261 29696 19295
rect 29644 19252 29696 19261
rect 31208 19252 31260 19304
rect 36084 19252 36136 19304
rect 36544 19184 36596 19236
rect 27160 19159 27212 19168
rect 27160 19125 27169 19159
rect 27169 19125 27203 19159
rect 27203 19125 27212 19159
rect 27160 19116 27212 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 4712 18912 4764 18964
rect 7012 18912 7064 18964
rect 12992 18912 13044 18964
rect 13452 18955 13504 18964
rect 13452 18921 13461 18955
rect 13461 18921 13495 18955
rect 13495 18921 13504 18955
rect 13452 18912 13504 18921
rect 23204 18955 23256 18964
rect 14740 18844 14792 18896
rect 4620 18776 4672 18828
rect 18512 18844 18564 18896
rect 23204 18921 23213 18955
rect 23213 18921 23247 18955
rect 23247 18921 23256 18955
rect 23204 18912 23256 18921
rect 26240 18912 26292 18964
rect 26884 18955 26936 18964
rect 26884 18921 26893 18955
rect 26893 18921 26927 18955
rect 26927 18921 26936 18955
rect 26884 18912 26936 18921
rect 28264 18912 28316 18964
rect 27528 18844 27580 18896
rect 36084 18887 36136 18896
rect 2872 18708 2924 18760
rect 2964 18751 3016 18760
rect 2964 18717 2973 18751
rect 2973 18717 3007 18751
rect 3007 18717 3016 18751
rect 3976 18751 4028 18760
rect 2964 18708 3016 18717
rect 3976 18717 3985 18751
rect 3985 18717 4019 18751
rect 4019 18717 4028 18751
rect 3976 18708 4028 18717
rect 7104 18708 7156 18760
rect 10600 18708 10652 18760
rect 2136 18572 2188 18624
rect 4896 18640 4948 18692
rect 6736 18683 6788 18692
rect 6736 18649 6745 18683
rect 6745 18649 6779 18683
rect 6779 18649 6788 18683
rect 6736 18640 6788 18649
rect 10692 18640 10744 18692
rect 17224 18640 17276 18692
rect 17868 18708 17920 18760
rect 20260 18776 20312 18828
rect 36084 18853 36093 18887
rect 36093 18853 36127 18887
rect 36127 18853 36136 18887
rect 36084 18844 36136 18853
rect 22376 18708 22428 18760
rect 23664 18751 23716 18760
rect 18696 18640 18748 18692
rect 21916 18640 21968 18692
rect 22192 18683 22244 18692
rect 22192 18649 22201 18683
rect 22201 18649 22235 18683
rect 22235 18649 22244 18683
rect 22192 18640 22244 18649
rect 4436 18572 4488 18624
rect 5724 18615 5776 18624
rect 5724 18581 5733 18615
rect 5733 18581 5767 18615
rect 5767 18581 5776 18615
rect 5724 18572 5776 18581
rect 9128 18572 9180 18624
rect 10140 18615 10192 18624
rect 10140 18581 10149 18615
rect 10149 18581 10183 18615
rect 10183 18581 10192 18615
rect 10140 18572 10192 18581
rect 14832 18572 14884 18624
rect 16856 18572 16908 18624
rect 17316 18572 17368 18624
rect 17592 18572 17644 18624
rect 22560 18572 22612 18624
rect 23664 18717 23673 18751
rect 23673 18717 23707 18751
rect 23707 18717 23716 18751
rect 23664 18708 23716 18717
rect 25228 18708 25280 18760
rect 26056 18708 26108 18760
rect 23848 18640 23900 18692
rect 27160 18640 27212 18692
rect 25872 18572 25924 18624
rect 30380 18819 30432 18828
rect 30380 18785 30389 18819
rect 30389 18785 30423 18819
rect 30423 18785 30432 18819
rect 30380 18776 30432 18785
rect 30932 18776 30984 18828
rect 33140 18776 33192 18828
rect 28448 18708 28500 18760
rect 31024 18708 31076 18760
rect 33784 18708 33836 18760
rect 35716 18751 35768 18760
rect 35716 18717 35725 18751
rect 35725 18717 35759 18751
rect 35759 18717 35768 18751
rect 35716 18708 35768 18717
rect 30840 18640 30892 18692
rect 30196 18572 30248 18624
rect 31024 18572 31076 18624
rect 35348 18640 35400 18692
rect 35992 18708 36044 18760
rect 36452 18751 36504 18760
rect 36452 18717 36461 18751
rect 36461 18717 36495 18751
rect 36495 18717 36504 18751
rect 36452 18708 36504 18717
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 2136 18343 2188 18352
rect 2136 18309 2145 18343
rect 2145 18309 2179 18343
rect 2179 18309 2188 18343
rect 2136 18300 2188 18309
rect 2780 18300 2832 18352
rect 3976 18368 4028 18420
rect 13360 18368 13412 18420
rect 15568 18368 15620 18420
rect 15936 18368 15988 18420
rect 26056 18411 26108 18420
rect 26056 18377 26065 18411
rect 26065 18377 26099 18411
rect 26099 18377 26108 18411
rect 26056 18368 26108 18377
rect 29644 18368 29696 18420
rect 32220 18368 32272 18420
rect 2688 18164 2740 18216
rect 4804 18232 4856 18284
rect 5448 18232 5500 18284
rect 4712 18164 4764 18216
rect 4436 18139 4488 18148
rect 4436 18105 4445 18139
rect 4445 18105 4479 18139
rect 4479 18105 4488 18139
rect 4436 18096 4488 18105
rect 9220 18232 9272 18284
rect 13820 18300 13872 18352
rect 17868 18300 17920 18352
rect 18880 18343 18932 18352
rect 18880 18309 18889 18343
rect 18889 18309 18923 18343
rect 18923 18309 18932 18343
rect 18880 18300 18932 18309
rect 22560 18343 22612 18352
rect 22560 18309 22569 18343
rect 22569 18309 22603 18343
rect 22603 18309 22612 18343
rect 22560 18300 22612 18309
rect 10600 18275 10652 18284
rect 10600 18241 10609 18275
rect 10609 18241 10643 18275
rect 10643 18241 10652 18275
rect 10600 18232 10652 18241
rect 12900 18275 12952 18284
rect 12900 18241 12909 18275
rect 12909 18241 12943 18275
rect 12943 18241 12952 18275
rect 12900 18232 12952 18241
rect 17224 18275 17276 18284
rect 17224 18241 17233 18275
rect 17233 18241 17267 18275
rect 17267 18241 17276 18275
rect 17224 18232 17276 18241
rect 17592 18275 17644 18284
rect 17592 18241 17601 18275
rect 17601 18241 17635 18275
rect 17635 18241 17644 18275
rect 17592 18232 17644 18241
rect 18512 18275 18564 18284
rect 18512 18241 18521 18275
rect 18521 18241 18555 18275
rect 18555 18241 18564 18275
rect 18512 18232 18564 18241
rect 18604 18232 18656 18284
rect 9404 18164 9456 18216
rect 26240 18232 26292 18284
rect 28632 18275 28684 18284
rect 28632 18241 28641 18275
rect 28641 18241 28675 18275
rect 28675 18241 28684 18275
rect 28632 18232 28684 18241
rect 30840 18275 30892 18284
rect 30840 18241 30849 18275
rect 30849 18241 30883 18275
rect 30883 18241 30892 18275
rect 30840 18232 30892 18241
rect 31024 18275 31076 18284
rect 31024 18241 31033 18275
rect 31033 18241 31067 18275
rect 31067 18241 31076 18275
rect 31024 18232 31076 18241
rect 32772 18275 32824 18284
rect 32772 18241 32781 18275
rect 32781 18241 32815 18275
rect 32815 18241 32824 18275
rect 32772 18232 32824 18241
rect 35992 18368 36044 18420
rect 36176 18411 36228 18420
rect 36176 18377 36185 18411
rect 36185 18377 36219 18411
rect 36219 18377 36228 18411
rect 36176 18368 36228 18377
rect 33324 18275 33376 18284
rect 33324 18241 33333 18275
rect 33333 18241 33367 18275
rect 33367 18241 33376 18275
rect 33324 18232 33376 18241
rect 35716 18300 35768 18352
rect 36452 18300 36504 18352
rect 27436 18164 27488 18216
rect 32864 18164 32916 18216
rect 33600 18164 33652 18216
rect 5448 18028 5500 18080
rect 10692 18028 10744 18080
rect 16488 18096 16540 18148
rect 32588 18096 32640 18148
rect 20812 18028 20864 18080
rect 29000 18028 29052 18080
rect 32772 18028 32824 18080
rect 34796 18207 34848 18216
rect 34796 18173 34805 18207
rect 34805 18173 34839 18207
rect 34839 18173 34848 18207
rect 34796 18164 34848 18173
rect 35716 18164 35768 18216
rect 35348 18096 35400 18148
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 2780 17867 2832 17876
rect 2780 17833 2789 17867
rect 2789 17833 2823 17867
rect 2823 17833 2832 17867
rect 2780 17824 2832 17833
rect 1400 17688 1452 17740
rect 2780 17663 2832 17672
rect 2780 17629 2789 17663
rect 2789 17629 2823 17663
rect 2823 17629 2832 17663
rect 2780 17620 2832 17629
rect 5080 17620 5132 17672
rect 8300 17552 8352 17604
rect 8484 17663 8536 17672
rect 8484 17629 8493 17663
rect 8493 17629 8527 17663
rect 8527 17629 8536 17663
rect 10600 17824 10652 17876
rect 22008 17824 22060 17876
rect 25044 17824 25096 17876
rect 25412 17824 25464 17876
rect 27804 17824 27856 17876
rect 33416 17867 33468 17876
rect 33416 17833 33425 17867
rect 33425 17833 33459 17867
rect 33459 17833 33468 17867
rect 33416 17824 33468 17833
rect 21548 17756 21600 17808
rect 23480 17756 23532 17808
rect 28448 17731 28500 17740
rect 8484 17620 8536 17629
rect 9128 17663 9180 17672
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 12164 17620 12216 17672
rect 17408 17620 17460 17672
rect 17868 17620 17920 17672
rect 18696 17663 18748 17672
rect 18696 17629 18705 17663
rect 18705 17629 18739 17663
rect 18739 17629 18748 17663
rect 18696 17620 18748 17629
rect 19248 17620 19300 17672
rect 9404 17595 9456 17604
rect 9404 17561 9413 17595
rect 9413 17561 9447 17595
rect 9447 17561 9456 17595
rect 9404 17552 9456 17561
rect 10784 17552 10836 17604
rect 13360 17552 13412 17604
rect 28448 17697 28457 17731
rect 28457 17697 28491 17731
rect 28491 17697 28500 17731
rect 28448 17688 28500 17697
rect 29000 17756 29052 17808
rect 20628 17620 20680 17672
rect 23480 17663 23532 17672
rect 23480 17629 23489 17663
rect 23489 17629 23523 17663
rect 23523 17629 23532 17663
rect 23480 17620 23532 17629
rect 30380 17688 30432 17740
rect 33600 17731 33652 17740
rect 33600 17697 33609 17731
rect 33609 17697 33643 17731
rect 33643 17697 33652 17731
rect 33600 17688 33652 17697
rect 29736 17663 29788 17672
rect 20812 17595 20864 17604
rect 6828 17484 6880 17536
rect 10140 17484 10192 17536
rect 10968 17484 11020 17536
rect 13728 17527 13780 17536
rect 13728 17493 13737 17527
rect 13737 17493 13771 17527
rect 13771 17493 13780 17527
rect 13728 17484 13780 17493
rect 16488 17484 16540 17536
rect 17316 17484 17368 17536
rect 18420 17484 18472 17536
rect 20812 17561 20821 17595
rect 20821 17561 20855 17595
rect 20855 17561 20864 17595
rect 20812 17552 20864 17561
rect 21916 17552 21968 17604
rect 24860 17595 24912 17604
rect 24860 17561 24869 17595
rect 24869 17561 24903 17595
rect 24903 17561 24912 17595
rect 24860 17552 24912 17561
rect 27252 17552 27304 17604
rect 29736 17629 29745 17663
rect 29745 17629 29779 17663
rect 29779 17629 29788 17663
rect 29736 17620 29788 17629
rect 32220 17620 32272 17672
rect 32588 17663 32640 17672
rect 32588 17629 32597 17663
rect 32597 17629 32631 17663
rect 32631 17629 32640 17663
rect 32588 17620 32640 17629
rect 33048 17620 33100 17672
rect 33784 17663 33836 17672
rect 33784 17629 33793 17663
rect 33793 17629 33827 17663
rect 33827 17629 33836 17663
rect 33784 17620 33836 17629
rect 32680 17595 32732 17604
rect 32680 17561 32689 17595
rect 32689 17561 32723 17595
rect 32723 17561 32732 17595
rect 34796 17620 34848 17672
rect 32680 17552 32732 17561
rect 23020 17527 23072 17536
rect 23020 17493 23029 17527
rect 23029 17493 23063 17527
rect 23063 17493 23072 17527
rect 23020 17484 23072 17493
rect 23388 17527 23440 17536
rect 23388 17493 23397 17527
rect 23397 17493 23431 17527
rect 23431 17493 23440 17527
rect 23388 17484 23440 17493
rect 25136 17484 25188 17536
rect 26240 17484 26292 17536
rect 28632 17484 28684 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 5356 17187 5408 17196
rect 5356 17153 5365 17187
rect 5365 17153 5399 17187
rect 5399 17153 5408 17187
rect 5356 17144 5408 17153
rect 5724 17280 5776 17332
rect 8484 17280 8536 17332
rect 10324 17280 10376 17332
rect 18144 17280 18196 17332
rect 22376 17280 22428 17332
rect 30196 17280 30248 17332
rect 33140 17323 33192 17332
rect 33140 17289 33149 17323
rect 33149 17289 33183 17323
rect 33183 17289 33192 17323
rect 33140 17280 33192 17289
rect 5908 17212 5960 17264
rect 7656 17144 7708 17196
rect 10692 17187 10744 17196
rect 10692 17153 10701 17187
rect 10701 17153 10735 17187
rect 10735 17153 10744 17187
rect 10692 17144 10744 17153
rect 10968 17212 11020 17264
rect 13268 17144 13320 17196
rect 14648 17187 14700 17196
rect 14648 17153 14657 17187
rect 14657 17153 14691 17187
rect 14691 17153 14700 17187
rect 14648 17144 14700 17153
rect 18052 17212 18104 17264
rect 21916 17212 21968 17264
rect 17316 17144 17368 17196
rect 5264 17119 5316 17128
rect 5264 17085 5273 17119
rect 5273 17085 5307 17119
rect 5307 17085 5316 17119
rect 5264 17076 5316 17085
rect 5356 17008 5408 17060
rect 10600 17076 10652 17128
rect 12164 17076 12216 17128
rect 15016 17119 15068 17128
rect 15016 17085 15025 17119
rect 15025 17085 15059 17119
rect 15059 17085 15068 17119
rect 15016 17076 15068 17085
rect 10232 17008 10284 17060
rect 10784 17051 10836 17060
rect 10784 17017 10793 17051
rect 10793 17017 10827 17051
rect 10827 17017 10836 17051
rect 10784 17008 10836 17017
rect 16856 17008 16908 17060
rect 18328 17187 18380 17196
rect 18328 17153 18338 17187
rect 18338 17153 18372 17187
rect 18372 17153 18380 17187
rect 18328 17144 18380 17153
rect 18696 17187 18748 17196
rect 18420 17076 18472 17128
rect 18696 17153 18710 17187
rect 18710 17153 18744 17187
rect 18744 17153 18748 17187
rect 18696 17144 18748 17153
rect 21180 17187 21232 17196
rect 21180 17153 21189 17187
rect 21189 17153 21223 17187
rect 21223 17153 21232 17187
rect 21180 17144 21232 17153
rect 21548 17144 21600 17196
rect 22008 17187 22060 17196
rect 22008 17153 22017 17187
rect 22017 17153 22051 17187
rect 22051 17153 22060 17187
rect 22008 17144 22060 17153
rect 23020 17144 23072 17196
rect 33416 17212 33468 17264
rect 23940 17144 23992 17196
rect 21824 17076 21876 17128
rect 22008 17008 22060 17060
rect 32680 17187 32732 17196
rect 32680 17153 32689 17187
rect 32689 17153 32723 17187
rect 32723 17153 32732 17187
rect 32680 17144 32732 17153
rect 33508 17144 33560 17196
rect 33232 17076 33284 17128
rect 34796 17144 34848 17196
rect 33508 17008 33560 17060
rect 6552 16940 6604 16992
rect 9496 16940 9548 16992
rect 14096 16983 14148 16992
rect 14096 16949 14105 16983
rect 14105 16949 14139 16983
rect 14139 16949 14148 16983
rect 14096 16940 14148 16949
rect 17408 16940 17460 16992
rect 21088 16940 21140 16992
rect 23388 16983 23440 16992
rect 23388 16949 23397 16983
rect 23397 16949 23431 16983
rect 23431 16949 23440 16983
rect 23388 16940 23440 16949
rect 25228 16983 25280 16992
rect 25228 16949 25237 16983
rect 25237 16949 25271 16983
rect 25271 16949 25280 16983
rect 25228 16940 25280 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2872 16736 2924 16788
rect 5080 16736 5132 16788
rect 13268 16779 13320 16788
rect 4620 16668 4672 16720
rect 5080 16643 5132 16652
rect 5080 16609 5089 16643
rect 5089 16609 5123 16643
rect 5123 16609 5132 16643
rect 5080 16600 5132 16609
rect 5356 16643 5408 16652
rect 5356 16609 5365 16643
rect 5365 16609 5399 16643
rect 5399 16609 5408 16643
rect 5356 16600 5408 16609
rect 13268 16745 13277 16779
rect 13277 16745 13311 16779
rect 13311 16745 13320 16779
rect 13268 16736 13320 16745
rect 21916 16736 21968 16788
rect 22008 16736 22060 16788
rect 23940 16736 23992 16788
rect 32864 16736 32916 16788
rect 33784 16736 33836 16788
rect 36728 16779 36780 16788
rect 36728 16745 36737 16779
rect 36737 16745 36771 16779
rect 36771 16745 36780 16779
rect 36728 16736 36780 16745
rect 28172 16668 28224 16720
rect 22008 16600 22060 16652
rect 26332 16600 26384 16652
rect 13452 16575 13504 16584
rect 13452 16541 13461 16575
rect 13461 16541 13495 16575
rect 13495 16541 13504 16575
rect 13452 16532 13504 16541
rect 13636 16532 13688 16584
rect 17408 16575 17460 16584
rect 2964 16464 3016 16516
rect 4712 16464 4764 16516
rect 6000 16464 6052 16516
rect 7656 16507 7708 16516
rect 7656 16473 7665 16507
rect 7665 16473 7699 16507
rect 7699 16473 7708 16507
rect 7656 16464 7708 16473
rect 6184 16396 6236 16448
rect 16856 16464 16908 16516
rect 17408 16541 17417 16575
rect 17417 16541 17451 16575
rect 17451 16541 17460 16575
rect 17408 16532 17460 16541
rect 17684 16575 17736 16584
rect 17684 16541 17693 16575
rect 17693 16541 17727 16575
rect 17727 16541 17736 16575
rect 17684 16532 17736 16541
rect 20720 16532 20772 16584
rect 20904 16532 20956 16584
rect 21088 16532 21140 16584
rect 21824 16532 21876 16584
rect 23572 16575 23624 16584
rect 23572 16541 23581 16575
rect 23581 16541 23615 16575
rect 23615 16541 23624 16575
rect 23572 16532 23624 16541
rect 23664 16532 23716 16584
rect 26148 16532 26200 16584
rect 17960 16464 18012 16516
rect 18604 16464 18656 16516
rect 24860 16464 24912 16516
rect 25228 16464 25280 16516
rect 26056 16464 26108 16516
rect 29460 16532 29512 16584
rect 33232 16575 33284 16584
rect 33232 16541 33241 16575
rect 33241 16541 33275 16575
rect 33275 16541 33284 16575
rect 33232 16532 33284 16541
rect 33508 16575 33560 16584
rect 33508 16541 33517 16575
rect 33517 16541 33551 16575
rect 33551 16541 33560 16575
rect 33508 16532 33560 16541
rect 34336 16532 34388 16584
rect 28540 16464 28592 16516
rect 35900 16507 35952 16516
rect 35900 16473 35909 16507
rect 35909 16473 35943 16507
rect 35943 16473 35952 16507
rect 35900 16464 35952 16473
rect 36912 16575 36964 16584
rect 36912 16541 36921 16575
rect 36921 16541 36955 16575
rect 36955 16541 36964 16575
rect 36912 16532 36964 16541
rect 37188 16575 37240 16584
rect 37188 16541 37197 16575
rect 37197 16541 37231 16575
rect 37231 16541 37240 16575
rect 37188 16532 37240 16541
rect 37832 16464 37884 16516
rect 14096 16396 14148 16448
rect 14648 16396 14700 16448
rect 22376 16439 22428 16448
rect 22376 16405 22385 16439
rect 22385 16405 22419 16439
rect 22419 16405 22428 16439
rect 22376 16396 22428 16405
rect 25780 16439 25832 16448
rect 25780 16405 25789 16439
rect 25789 16405 25823 16439
rect 25823 16405 25832 16439
rect 25780 16396 25832 16405
rect 26148 16439 26200 16448
rect 26148 16405 26157 16439
rect 26157 16405 26191 16439
rect 26191 16405 26200 16439
rect 26148 16396 26200 16405
rect 30932 16396 30984 16448
rect 33416 16439 33468 16448
rect 33416 16405 33425 16439
rect 33425 16405 33459 16439
rect 33459 16405 33468 16439
rect 33416 16396 33468 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 5080 16192 5132 16244
rect 3240 16124 3292 16176
rect 6000 16167 6052 16176
rect 5540 16056 5592 16108
rect 6000 16133 6009 16167
rect 6009 16133 6043 16167
rect 6043 16133 6052 16167
rect 6000 16124 6052 16133
rect 9128 16192 9180 16244
rect 13360 16235 13412 16244
rect 13360 16201 13369 16235
rect 13369 16201 13403 16235
rect 13403 16201 13412 16235
rect 13360 16192 13412 16201
rect 6828 16167 6880 16176
rect 5908 16099 5960 16108
rect 5908 16065 5917 16099
rect 5917 16065 5951 16099
rect 5951 16065 5960 16099
rect 5908 16056 5960 16065
rect 6828 16133 6837 16167
rect 6837 16133 6871 16167
rect 6871 16133 6880 16167
rect 6828 16124 6880 16133
rect 7288 16124 7340 16176
rect 9956 16124 10008 16176
rect 9128 16056 9180 16108
rect 15016 16192 15068 16244
rect 15200 16235 15252 16244
rect 15200 16201 15209 16235
rect 15209 16201 15243 16235
rect 15243 16201 15252 16235
rect 15200 16192 15252 16201
rect 21272 16192 21324 16244
rect 28540 16235 28592 16244
rect 28540 16201 28549 16235
rect 28549 16201 28583 16235
rect 28583 16201 28592 16235
rect 28540 16192 28592 16201
rect 35900 16235 35952 16244
rect 35900 16201 35909 16235
rect 35909 16201 35943 16235
rect 35943 16201 35952 16235
rect 35900 16192 35952 16201
rect 37188 16192 37240 16244
rect 37832 16235 37884 16244
rect 37832 16201 37841 16235
rect 37841 16201 37875 16235
rect 37875 16201 37884 16235
rect 37832 16192 37884 16201
rect 13636 16124 13688 16176
rect 14832 16167 14884 16176
rect 13728 16099 13780 16108
rect 13728 16065 13737 16099
rect 13737 16065 13771 16099
rect 13771 16065 13780 16099
rect 13728 16056 13780 16065
rect 14832 16133 14841 16167
rect 14841 16133 14875 16167
rect 14875 16133 14884 16167
rect 14832 16124 14884 16133
rect 16672 16124 16724 16176
rect 17684 16124 17736 16176
rect 5448 15988 5500 16040
rect 6828 15988 6880 16040
rect 9496 16031 9548 16040
rect 9496 15997 9505 16031
rect 9505 15997 9539 16031
rect 9539 15997 9548 16031
rect 9496 15988 9548 15997
rect 14648 16099 14700 16108
rect 14648 16065 14658 16099
rect 14658 16065 14692 16099
rect 14692 16065 14700 16099
rect 14648 16056 14700 16065
rect 14924 16099 14976 16108
rect 14924 16065 14933 16099
rect 14933 16065 14967 16099
rect 14967 16065 14976 16099
rect 14924 16056 14976 16065
rect 16028 16056 16080 16108
rect 16856 16099 16908 16108
rect 16856 16065 16865 16099
rect 16865 16065 16899 16099
rect 16899 16065 16908 16099
rect 16856 16056 16908 16065
rect 17224 16099 17276 16108
rect 17224 16065 17233 16099
rect 17233 16065 17267 16099
rect 17267 16065 17276 16099
rect 17224 16056 17276 16065
rect 17316 16056 17368 16108
rect 17868 16056 17920 16108
rect 18512 16056 18564 16108
rect 23388 16124 23440 16176
rect 25780 16124 25832 16176
rect 30932 16124 30984 16176
rect 21272 16099 21324 16108
rect 16396 15988 16448 16040
rect 21272 16065 21281 16099
rect 21281 16065 21315 16099
rect 21315 16065 21324 16099
rect 21272 16056 21324 16065
rect 21364 16099 21416 16108
rect 21364 16065 21373 16099
rect 21373 16065 21407 16099
rect 21407 16065 21416 16099
rect 21364 16056 21416 16065
rect 22192 15988 22244 16040
rect 24676 15988 24728 16040
rect 29000 16099 29052 16108
rect 29000 16065 29009 16099
rect 29009 16065 29043 16099
rect 29043 16065 29052 16099
rect 29000 16056 29052 16065
rect 30656 16056 30708 16108
rect 37372 16124 37424 16176
rect 36360 16056 36412 16108
rect 29092 15988 29144 16040
rect 29460 16031 29512 16040
rect 29460 15997 29469 16031
rect 29469 15997 29503 16031
rect 29503 15997 29512 16031
rect 29460 15988 29512 15997
rect 36452 16031 36504 16040
rect 36452 15997 36461 16031
rect 36461 15997 36495 16031
rect 36495 15997 36504 16031
rect 36452 15988 36504 15997
rect 36636 16099 36688 16108
rect 36636 16065 36645 16099
rect 36645 16065 36679 16099
rect 36679 16065 36688 16099
rect 36636 16056 36688 16065
rect 16856 15920 16908 15972
rect 35900 15920 35952 15972
rect 36636 15920 36688 15972
rect 8208 15852 8260 15904
rect 10508 15852 10560 15904
rect 25044 15852 25096 15904
rect 26148 15852 26200 15904
rect 31208 15852 31260 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 30656 15691 30708 15700
rect 30656 15657 30665 15691
rect 30665 15657 30699 15691
rect 30699 15657 30708 15691
rect 30656 15648 30708 15657
rect 33416 15648 33468 15700
rect 34336 15648 34388 15700
rect 37372 15691 37424 15700
rect 37372 15657 37381 15691
rect 37381 15657 37415 15691
rect 37415 15657 37424 15691
rect 37372 15648 37424 15657
rect 8208 15580 8260 15632
rect 7288 15512 7340 15564
rect 9956 15555 10008 15564
rect 5540 15444 5592 15496
rect 7656 15444 7708 15496
rect 9956 15521 9965 15555
rect 9965 15521 9999 15555
rect 9999 15521 10008 15555
rect 9956 15512 10008 15521
rect 12164 15555 12216 15564
rect 12164 15521 12173 15555
rect 12173 15521 12207 15555
rect 12207 15521 12216 15555
rect 12164 15512 12216 15521
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 14004 15444 14056 15496
rect 36912 15580 36964 15632
rect 16672 15555 16724 15564
rect 16672 15521 16681 15555
rect 16681 15521 16715 15555
rect 16715 15521 16724 15555
rect 16672 15512 16724 15521
rect 17592 15512 17644 15564
rect 10508 15376 10560 15428
rect 16856 15444 16908 15496
rect 18696 15512 18748 15564
rect 24676 15512 24728 15564
rect 29000 15512 29052 15564
rect 30196 15512 30248 15564
rect 19156 15444 19208 15496
rect 19248 15444 19300 15496
rect 16764 15376 16816 15428
rect 24860 15444 24912 15496
rect 25044 15487 25096 15496
rect 25044 15453 25053 15487
rect 25053 15453 25087 15487
rect 25087 15453 25096 15487
rect 25044 15444 25096 15453
rect 25136 15487 25188 15496
rect 25136 15453 25145 15487
rect 25145 15453 25179 15487
rect 25179 15453 25188 15487
rect 25136 15444 25188 15453
rect 29552 15444 29604 15496
rect 20260 15376 20312 15428
rect 22192 15376 22244 15428
rect 26148 15376 26200 15428
rect 33692 15444 33744 15496
rect 34888 15512 34940 15564
rect 36360 15555 36412 15564
rect 36360 15521 36369 15555
rect 36369 15521 36403 15555
rect 36403 15521 36412 15555
rect 36360 15512 36412 15521
rect 31392 15376 31444 15428
rect 13452 15308 13504 15360
rect 17040 15308 17092 15360
rect 25872 15308 25924 15360
rect 26516 15308 26568 15360
rect 31208 15308 31260 15360
rect 34704 15444 34756 15496
rect 36544 15487 36596 15496
rect 36544 15453 36553 15487
rect 36553 15453 36587 15487
rect 36587 15453 36596 15487
rect 36544 15444 36596 15453
rect 36912 15487 36964 15496
rect 36912 15453 36921 15487
rect 36921 15453 36955 15487
rect 36955 15453 36964 15487
rect 36912 15444 36964 15453
rect 37188 15444 37240 15496
rect 34796 15376 34848 15428
rect 35164 15308 35216 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 2136 15104 2188 15156
rect 7104 15104 7156 15156
rect 21364 15104 21416 15156
rect 26148 15147 26200 15156
rect 26148 15113 26157 15147
rect 26157 15113 26191 15147
rect 26191 15113 26200 15147
rect 26148 15104 26200 15113
rect 26516 15147 26568 15156
rect 26516 15113 26525 15147
rect 26525 15113 26559 15147
rect 26559 15113 26568 15147
rect 26516 15104 26568 15113
rect 28172 15147 28224 15156
rect 28172 15113 28181 15147
rect 28181 15113 28215 15147
rect 28215 15113 28224 15147
rect 28172 15104 28224 15113
rect 32772 15104 32824 15156
rect 13728 15036 13780 15088
rect 20904 15079 20956 15088
rect 13912 15011 13964 15020
rect 2688 14900 2740 14952
rect 3148 14900 3200 14952
rect 13912 14977 13921 15011
rect 13921 14977 13955 15011
rect 13955 14977 13964 15011
rect 13912 14968 13964 14977
rect 16856 15011 16908 15020
rect 16856 14977 16865 15011
rect 16865 14977 16899 15011
rect 16899 14977 16908 15011
rect 16856 14968 16908 14977
rect 4712 14900 4764 14952
rect 3792 14807 3844 14816
rect 3792 14773 3801 14807
rect 3801 14773 3835 14807
rect 3835 14773 3844 14807
rect 3792 14764 3844 14773
rect 14188 14943 14240 14952
rect 14188 14909 14197 14943
rect 14197 14909 14231 14943
rect 14231 14909 14240 14943
rect 14188 14900 14240 14909
rect 16764 14900 16816 14952
rect 17868 14968 17920 15020
rect 18512 14968 18564 15020
rect 19156 14968 19208 15020
rect 20904 15045 20913 15079
rect 20913 15045 20947 15079
rect 20947 15045 20956 15079
rect 20904 15036 20956 15045
rect 22284 15036 22336 15088
rect 25320 15036 25372 15088
rect 26056 15036 26108 15088
rect 19248 14832 19300 14884
rect 19340 14764 19392 14816
rect 21180 14968 21232 15020
rect 24124 14968 24176 15020
rect 26332 15011 26384 15020
rect 26332 14977 26341 15011
rect 26341 14977 26375 15011
rect 26375 14977 26384 15011
rect 26332 14968 26384 14977
rect 31852 15036 31904 15088
rect 28448 15011 28500 15020
rect 28448 14977 28457 15011
rect 28457 14977 28491 15011
rect 28491 14977 28500 15011
rect 28448 14968 28500 14977
rect 28724 14968 28776 15020
rect 30564 15011 30616 15020
rect 30564 14977 30573 15011
rect 30573 14977 30607 15011
rect 30607 14977 30616 15011
rect 30564 14968 30616 14977
rect 30932 15011 30984 15020
rect 30932 14977 30941 15011
rect 30941 14977 30975 15011
rect 30975 14977 30984 15011
rect 30932 14968 30984 14977
rect 21088 14832 21140 14884
rect 25136 14764 25188 14816
rect 26424 14764 26476 14816
rect 31208 14900 31260 14952
rect 33048 14968 33100 15020
rect 33508 14968 33560 15020
rect 34520 15104 34572 15156
rect 34612 15036 34664 15088
rect 36912 15104 36964 15156
rect 35164 15079 35216 15088
rect 35164 15045 35173 15079
rect 35173 15045 35207 15079
rect 35207 15045 35216 15079
rect 35164 15036 35216 15045
rect 34888 14968 34940 15020
rect 34704 14900 34756 14952
rect 34520 14832 34572 14884
rect 35900 14968 35952 15020
rect 35348 14900 35400 14952
rect 31208 14764 31260 14816
rect 33600 14764 33652 14816
rect 33692 14764 33744 14816
rect 34888 14764 34940 14816
rect 35808 14764 35860 14816
rect 36176 14764 36228 14816
rect 36544 14764 36596 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 1676 14560 1728 14612
rect 3056 14560 3108 14612
rect 3976 14560 4028 14612
rect 16396 14560 16448 14612
rect 28724 14560 28776 14612
rect 30564 14560 30616 14612
rect 33048 14560 33100 14612
rect 34796 14560 34848 14612
rect 37188 14560 37240 14612
rect 3056 14467 3108 14476
rect 3056 14433 3065 14467
rect 3065 14433 3099 14467
rect 3099 14433 3108 14467
rect 3056 14424 3108 14433
rect 3148 14467 3200 14476
rect 3148 14433 3157 14467
rect 3157 14433 3191 14467
rect 3191 14433 3200 14467
rect 3148 14424 3200 14433
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 2136 14356 2188 14365
rect 2780 14356 2832 14408
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 13452 14399 13504 14408
rect 3240 14356 3292 14365
rect 13452 14365 13461 14399
rect 13461 14365 13495 14399
rect 13495 14365 13504 14399
rect 13452 14356 13504 14365
rect 14188 14356 14240 14408
rect 15476 14356 15528 14408
rect 16672 14424 16724 14476
rect 17960 14424 18012 14476
rect 16212 14399 16264 14408
rect 16212 14365 16221 14399
rect 16221 14365 16255 14399
rect 16255 14365 16264 14399
rect 16212 14356 16264 14365
rect 16764 14399 16816 14408
rect 16764 14365 16773 14399
rect 16773 14365 16807 14399
rect 16807 14365 16816 14399
rect 16764 14356 16816 14365
rect 16856 14356 16908 14408
rect 18512 14424 18564 14476
rect 19064 14492 19116 14544
rect 21180 14492 21232 14544
rect 24124 14492 24176 14544
rect 18604 14399 18656 14408
rect 18604 14365 18613 14399
rect 18613 14365 18647 14399
rect 18647 14365 18656 14399
rect 18604 14356 18656 14365
rect 22376 14424 22428 14476
rect 23204 14467 23256 14476
rect 23204 14433 23213 14467
rect 23213 14433 23247 14467
rect 23247 14433 23256 14467
rect 23204 14424 23256 14433
rect 25320 14424 25372 14476
rect 20260 14399 20312 14408
rect 20260 14365 20269 14399
rect 20269 14365 20303 14399
rect 20303 14365 20312 14399
rect 20260 14356 20312 14365
rect 20444 14399 20496 14408
rect 20444 14365 20453 14399
rect 20453 14365 20487 14399
rect 20487 14365 20496 14399
rect 20444 14356 20496 14365
rect 22928 14399 22980 14408
rect 22928 14365 22937 14399
rect 22937 14365 22971 14399
rect 22971 14365 22980 14399
rect 22928 14356 22980 14365
rect 3792 14288 3844 14340
rect 20352 14331 20404 14340
rect 20352 14297 20361 14331
rect 20361 14297 20395 14331
rect 20395 14297 20404 14331
rect 20352 14288 20404 14297
rect 1860 14220 1912 14272
rect 2688 14220 2740 14272
rect 3056 14220 3108 14272
rect 3240 14220 3292 14272
rect 13268 14263 13320 14272
rect 13268 14229 13277 14263
rect 13277 14229 13311 14263
rect 13311 14229 13320 14263
rect 13268 14220 13320 14229
rect 14280 14220 14332 14272
rect 16028 14263 16080 14272
rect 16028 14229 16037 14263
rect 16037 14229 16071 14263
rect 16071 14229 16080 14263
rect 16028 14220 16080 14229
rect 26332 14399 26384 14408
rect 26332 14365 26342 14399
rect 26342 14365 26376 14399
rect 26376 14365 26384 14399
rect 30380 14492 30432 14544
rect 30932 14492 30984 14544
rect 26332 14356 26384 14365
rect 34520 14356 34572 14408
rect 26516 14331 26568 14340
rect 26516 14297 26525 14331
rect 26525 14297 26559 14331
rect 26559 14297 26568 14331
rect 26516 14288 26568 14297
rect 26792 14288 26844 14340
rect 31852 14288 31904 14340
rect 34612 14288 34664 14340
rect 35256 14399 35308 14408
rect 35256 14365 35270 14399
rect 35270 14365 35304 14399
rect 35304 14365 35308 14399
rect 35256 14356 35308 14365
rect 35808 14356 35860 14408
rect 36176 14399 36228 14408
rect 36176 14365 36185 14399
rect 36185 14365 36219 14399
rect 36219 14365 36228 14399
rect 36176 14356 36228 14365
rect 26700 14220 26752 14272
rect 33600 14220 33652 14272
rect 35900 14220 35952 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1676 14059 1728 14068
rect 1676 14025 1685 14059
rect 1685 14025 1719 14059
rect 1719 14025 1728 14059
rect 1676 14016 1728 14025
rect 2872 14016 2924 14068
rect 3424 14016 3476 14068
rect 14280 14059 14332 14068
rect 14280 14025 14289 14059
rect 14289 14025 14323 14059
rect 14323 14025 14332 14059
rect 14280 14016 14332 14025
rect 14924 14016 14976 14068
rect 16212 14016 16264 14068
rect 18604 14016 18656 14068
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 3976 13923 4028 13932
rect 3976 13889 3985 13923
rect 3985 13889 4019 13923
rect 4019 13889 4028 13923
rect 3976 13880 4028 13889
rect 13268 13948 13320 14000
rect 16948 13948 17000 14000
rect 26424 14016 26476 14068
rect 32680 14016 32732 14068
rect 35256 14016 35308 14068
rect 22284 13948 22336 14000
rect 23296 13948 23348 14000
rect 2780 13812 2832 13864
rect 3148 13812 3200 13864
rect 3792 13812 3844 13864
rect 3792 13676 3844 13728
rect 9496 13880 9548 13932
rect 15108 13923 15160 13932
rect 8760 13855 8812 13864
rect 8760 13821 8769 13855
rect 8769 13821 8803 13855
rect 8803 13821 8812 13855
rect 8760 13812 8812 13821
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 15108 13889 15117 13923
rect 15117 13889 15151 13923
rect 15151 13889 15160 13923
rect 15108 13880 15160 13889
rect 15476 13880 15528 13932
rect 17316 13880 17368 13932
rect 17960 13880 18012 13932
rect 18512 13880 18564 13932
rect 19156 13923 19208 13932
rect 19156 13889 19165 13923
rect 19165 13889 19199 13923
rect 19199 13889 19208 13923
rect 19156 13880 19208 13889
rect 15016 13812 15068 13864
rect 16304 13812 16356 13864
rect 22284 13812 22336 13864
rect 23204 13880 23256 13932
rect 24860 13880 24912 13932
rect 32404 13880 32456 13932
rect 25964 13812 26016 13864
rect 32312 13855 32364 13864
rect 32312 13821 32321 13855
rect 32321 13821 32355 13855
rect 32355 13821 32364 13855
rect 32312 13812 32364 13821
rect 29092 13744 29144 13796
rect 10140 13719 10192 13728
rect 10140 13685 10149 13719
rect 10149 13685 10183 13719
rect 10183 13685 10192 13719
rect 10140 13676 10192 13685
rect 14740 13719 14792 13728
rect 14740 13685 14749 13719
rect 14749 13685 14783 13719
rect 14783 13685 14792 13719
rect 14740 13676 14792 13685
rect 24584 13676 24636 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2780 13472 2832 13524
rect 3976 13472 4028 13524
rect 15752 13472 15804 13524
rect 19984 13404 20036 13456
rect 20444 13404 20496 13456
rect 3056 13336 3108 13388
rect 2780 13268 2832 13320
rect 3148 13311 3200 13320
rect 3148 13277 3157 13311
rect 3157 13277 3191 13311
rect 3191 13277 3200 13311
rect 3148 13268 3200 13277
rect 6644 13268 6696 13320
rect 9772 13336 9824 13388
rect 19156 13336 19208 13388
rect 21916 13472 21968 13524
rect 23388 13472 23440 13524
rect 28356 13472 28408 13524
rect 32312 13472 32364 13524
rect 24584 13379 24636 13388
rect 12900 13268 12952 13320
rect 16948 13268 17000 13320
rect 17316 13268 17368 13320
rect 18512 13311 18564 13320
rect 18512 13277 18521 13311
rect 18521 13277 18555 13311
rect 18555 13277 18564 13311
rect 18512 13268 18564 13277
rect 18604 13268 18656 13320
rect 2872 13243 2924 13252
rect 2872 13209 2890 13243
rect 2890 13209 2924 13243
rect 2872 13200 2924 13209
rect 3240 13200 3292 13252
rect 4160 13243 4212 13252
rect 4160 13209 4169 13243
rect 4169 13209 4203 13243
rect 4203 13209 4212 13243
rect 4160 13200 4212 13209
rect 4620 13200 4672 13252
rect 7472 13243 7524 13252
rect 7472 13209 7481 13243
rect 7481 13209 7515 13243
rect 7515 13209 7524 13243
rect 7472 13200 7524 13209
rect 7564 13243 7616 13252
rect 7564 13209 7573 13243
rect 7573 13209 7607 13243
rect 7607 13209 7616 13243
rect 7564 13200 7616 13209
rect 8208 13200 8260 13252
rect 8300 13243 8352 13252
rect 8300 13209 8309 13243
rect 8309 13209 8343 13243
rect 8343 13209 8352 13243
rect 8300 13200 8352 13209
rect 4344 13175 4396 13184
rect 4344 13141 4353 13175
rect 4353 13141 4387 13175
rect 4387 13141 4396 13175
rect 4344 13132 4396 13141
rect 6000 13132 6052 13184
rect 8484 13175 8536 13184
rect 8484 13141 8493 13175
rect 8493 13141 8527 13175
rect 8527 13141 8536 13175
rect 8484 13132 8536 13141
rect 12808 13200 12860 13252
rect 19248 13268 19300 13320
rect 20812 13311 20864 13320
rect 20812 13277 20821 13311
rect 20821 13277 20855 13311
rect 20855 13277 20864 13311
rect 20812 13268 20864 13277
rect 24584 13345 24593 13379
rect 24593 13345 24627 13379
rect 24627 13345 24636 13379
rect 24584 13336 24636 13345
rect 29092 13268 29144 13320
rect 30196 13311 30248 13320
rect 20444 13200 20496 13252
rect 27160 13200 27212 13252
rect 30196 13277 30205 13311
rect 30205 13277 30239 13311
rect 30239 13277 30248 13311
rect 30196 13268 30248 13277
rect 30472 13200 30524 13252
rect 32128 13200 32180 13252
rect 12992 13132 13044 13184
rect 19064 13132 19116 13184
rect 19432 13132 19484 13184
rect 26332 13132 26384 13184
rect 26608 13175 26660 13184
rect 26608 13141 26617 13175
rect 26617 13141 26651 13175
rect 26651 13141 26660 13175
rect 26608 13132 26660 13141
rect 29736 13175 29788 13184
rect 29736 13141 29745 13175
rect 29745 13141 29779 13175
rect 29779 13141 29788 13175
rect 29736 13132 29788 13141
rect 30564 13132 30616 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 4160 12928 4212 12980
rect 6000 12971 6052 12980
rect 6000 12937 6009 12971
rect 6009 12937 6043 12971
rect 6043 12937 6052 12971
rect 6000 12928 6052 12937
rect 10140 12928 10192 12980
rect 10232 12928 10284 12980
rect 3240 12903 3292 12912
rect 3240 12869 3249 12903
rect 3249 12869 3283 12903
rect 3283 12869 3292 12903
rect 3240 12860 3292 12869
rect 3976 12860 4028 12912
rect 4344 12860 4396 12912
rect 3148 12792 3200 12844
rect 4068 12792 4120 12844
rect 8760 12860 8812 12912
rect 10508 12903 10560 12912
rect 5448 12792 5500 12844
rect 7564 12792 7616 12844
rect 10048 12835 10100 12844
rect 10048 12801 10057 12835
rect 10057 12801 10091 12835
rect 10091 12801 10100 12835
rect 10048 12792 10100 12801
rect 10508 12869 10517 12903
rect 10517 12869 10551 12903
rect 10551 12869 10560 12903
rect 10508 12860 10560 12869
rect 15108 12928 15160 12980
rect 16948 12928 17000 12980
rect 17132 12928 17184 12980
rect 10416 12792 10468 12844
rect 10232 12724 10284 12776
rect 14188 12860 14240 12912
rect 15476 12860 15528 12912
rect 21272 12928 21324 12980
rect 24676 12971 24728 12980
rect 24676 12937 24685 12971
rect 24685 12937 24719 12971
rect 24719 12937 24728 12971
rect 24676 12928 24728 12937
rect 27160 12971 27212 12980
rect 27160 12937 27169 12971
rect 27169 12937 27203 12971
rect 27203 12937 27212 12971
rect 27160 12928 27212 12937
rect 29460 12928 29512 12980
rect 36176 12928 36228 12980
rect 12900 12792 12952 12844
rect 14740 12792 14792 12844
rect 15384 12835 15436 12844
rect 15384 12801 15393 12835
rect 15393 12801 15427 12835
rect 15427 12801 15436 12835
rect 15384 12792 15436 12801
rect 15568 12835 15620 12844
rect 15568 12801 15577 12835
rect 15577 12801 15611 12835
rect 15611 12801 15620 12835
rect 15568 12792 15620 12801
rect 18880 12860 18932 12912
rect 16948 12835 17000 12844
rect 16948 12801 16958 12835
rect 16958 12801 16992 12835
rect 16992 12801 17000 12835
rect 17132 12835 17184 12844
rect 16948 12792 17000 12801
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 17224 12835 17276 12844
rect 17224 12801 17233 12835
rect 17233 12801 17267 12835
rect 17267 12801 17276 12835
rect 17224 12792 17276 12801
rect 18696 12792 18748 12844
rect 18972 12835 19024 12844
rect 18972 12801 18981 12835
rect 18981 12801 19015 12835
rect 19015 12801 19024 12835
rect 18972 12792 19024 12801
rect 19156 12835 19208 12844
rect 19156 12801 19163 12835
rect 19163 12801 19208 12835
rect 19156 12792 19208 12801
rect 19432 12835 19484 12844
rect 19432 12801 19446 12835
rect 19446 12801 19480 12835
rect 19480 12801 19484 12835
rect 26240 12860 26292 12912
rect 26332 12860 26384 12912
rect 26792 12860 26844 12912
rect 28632 12903 28684 12912
rect 28632 12869 28641 12903
rect 28641 12869 28675 12903
rect 28675 12869 28684 12903
rect 28632 12860 28684 12869
rect 30196 12860 30248 12912
rect 25780 12835 25832 12844
rect 19432 12792 19484 12801
rect 25780 12801 25789 12835
rect 25789 12801 25823 12835
rect 25823 12801 25832 12835
rect 25780 12792 25832 12801
rect 3424 12631 3476 12640
rect 3424 12597 3433 12631
rect 3433 12597 3467 12631
rect 3467 12597 3476 12631
rect 3424 12588 3476 12597
rect 4620 12588 4672 12640
rect 11060 12631 11112 12640
rect 11060 12597 11069 12631
rect 11069 12597 11103 12631
rect 11103 12597 11112 12631
rect 11060 12588 11112 12597
rect 12624 12631 12676 12640
rect 12624 12597 12633 12631
rect 12633 12597 12667 12631
rect 12667 12597 12676 12631
rect 12624 12588 12676 12597
rect 12808 12631 12860 12640
rect 12808 12597 12817 12631
rect 12817 12597 12851 12631
rect 12851 12597 12860 12631
rect 12808 12588 12860 12597
rect 15200 12631 15252 12640
rect 15200 12597 15209 12631
rect 15209 12597 15243 12631
rect 15243 12597 15252 12631
rect 15200 12588 15252 12597
rect 23388 12656 23440 12708
rect 23572 12724 23624 12776
rect 26608 12792 26660 12844
rect 27344 12835 27396 12844
rect 27344 12801 27353 12835
rect 27353 12801 27387 12835
rect 27387 12801 27396 12835
rect 27344 12792 27396 12801
rect 26148 12724 26200 12776
rect 31116 12792 31168 12844
rect 32312 12835 32364 12844
rect 32312 12801 32321 12835
rect 32321 12801 32355 12835
rect 32355 12801 32364 12835
rect 32312 12792 32364 12801
rect 28080 12656 28132 12708
rect 16028 12588 16080 12640
rect 17132 12588 17184 12640
rect 18880 12588 18932 12640
rect 19248 12588 19300 12640
rect 23480 12588 23532 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 7472 12384 7524 12436
rect 10048 12384 10100 12436
rect 5448 12316 5500 12368
rect 4620 12248 4672 12300
rect 4068 12223 4120 12232
rect 4068 12189 4077 12223
rect 4077 12189 4111 12223
rect 4111 12189 4120 12223
rect 4068 12180 4120 12189
rect 4712 12180 4764 12232
rect 5264 12180 5316 12232
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 15476 12384 15528 12436
rect 15568 12384 15620 12436
rect 19156 12384 19208 12436
rect 23296 12427 23348 12436
rect 14280 12223 14332 12232
rect 9496 12112 9548 12164
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 14832 12180 14884 12232
rect 15292 12180 15344 12232
rect 21364 12316 21416 12368
rect 23296 12393 23305 12427
rect 23305 12393 23339 12427
rect 23339 12393 23348 12427
rect 23296 12384 23348 12393
rect 23848 12384 23900 12436
rect 25320 12384 25372 12436
rect 26056 12384 26108 12436
rect 26792 12427 26844 12436
rect 26792 12393 26801 12427
rect 26801 12393 26835 12427
rect 26835 12393 26844 12427
rect 26792 12384 26844 12393
rect 27252 12384 27304 12436
rect 28080 12427 28132 12436
rect 28080 12393 28089 12427
rect 28089 12393 28123 12427
rect 28123 12393 28132 12427
rect 28080 12384 28132 12393
rect 19064 12248 19116 12300
rect 20536 12248 20588 12300
rect 18512 12223 18564 12232
rect 18512 12189 18521 12223
rect 18521 12189 18555 12223
rect 18555 12189 18564 12223
rect 18512 12180 18564 12189
rect 15200 12112 15252 12164
rect 15568 12112 15620 12164
rect 4620 12044 4672 12096
rect 13268 12087 13320 12096
rect 13268 12053 13277 12087
rect 13277 12053 13311 12087
rect 13311 12053 13320 12087
rect 13268 12044 13320 12053
rect 13636 12087 13688 12096
rect 13636 12053 13645 12087
rect 13645 12053 13679 12087
rect 13679 12053 13688 12087
rect 13636 12044 13688 12053
rect 19524 12223 19576 12232
rect 19524 12189 19534 12223
rect 19534 12189 19568 12223
rect 19568 12189 19576 12223
rect 19524 12180 19576 12189
rect 19984 12180 20036 12232
rect 20904 12180 20956 12232
rect 21180 12223 21232 12232
rect 21180 12189 21189 12223
rect 21189 12189 21223 12223
rect 21223 12189 21232 12223
rect 21456 12223 21508 12232
rect 21180 12180 21232 12189
rect 21456 12189 21465 12223
rect 21465 12189 21499 12223
rect 21499 12189 21508 12223
rect 21456 12180 21508 12189
rect 19248 12112 19300 12164
rect 20168 12112 20220 12164
rect 24584 12248 24636 12300
rect 28448 12248 28500 12300
rect 30380 12248 30432 12300
rect 20996 12087 21048 12096
rect 20996 12053 21005 12087
rect 21005 12053 21039 12087
rect 21039 12053 21048 12087
rect 20996 12044 21048 12053
rect 21364 12087 21416 12096
rect 21364 12053 21373 12087
rect 21373 12053 21407 12087
rect 21407 12053 21416 12087
rect 21364 12044 21416 12053
rect 22284 12112 22336 12164
rect 24308 12112 24360 12164
rect 30288 12180 30340 12232
rect 24860 12044 24912 12096
rect 28540 12155 28592 12164
rect 28540 12121 28575 12155
rect 28575 12121 28592 12155
rect 30840 12155 30892 12164
rect 28540 12112 28592 12121
rect 30840 12121 30849 12155
rect 30849 12121 30883 12155
rect 30883 12121 30892 12155
rect 30840 12112 30892 12121
rect 30564 12044 30616 12096
rect 32128 12087 32180 12096
rect 32128 12053 32137 12087
rect 32137 12053 32171 12087
rect 32171 12053 32180 12087
rect 32128 12044 32180 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 23572 11840 23624 11892
rect 24124 11883 24176 11892
rect 24124 11849 24133 11883
rect 24133 11849 24167 11883
rect 24167 11849 24176 11883
rect 24124 11840 24176 11849
rect 24308 11883 24360 11892
rect 24308 11849 24317 11883
rect 24317 11849 24351 11883
rect 24351 11849 24360 11883
rect 24308 11840 24360 11849
rect 26792 11840 26844 11892
rect 28448 11883 28500 11892
rect 28448 11849 28457 11883
rect 28457 11849 28491 11883
rect 28491 11849 28500 11883
rect 28448 11840 28500 11849
rect 30840 11840 30892 11892
rect 32404 11840 32456 11892
rect 32680 11883 32732 11892
rect 32680 11849 32689 11883
rect 32689 11849 32723 11883
rect 32723 11849 32732 11883
rect 32680 11840 32732 11849
rect 16488 11704 16540 11756
rect 21456 11704 21508 11756
rect 23848 11772 23900 11824
rect 28264 11815 28316 11824
rect 14188 11636 14240 11688
rect 15108 11636 15160 11688
rect 22008 11636 22060 11688
rect 23480 11636 23532 11688
rect 16488 11568 16540 11620
rect 18236 11568 18288 11620
rect 23388 11568 23440 11620
rect 28264 11781 28273 11815
rect 28273 11781 28307 11815
rect 28307 11781 28316 11815
rect 28264 11772 28316 11781
rect 30196 11772 30248 11824
rect 25872 11747 25924 11756
rect 25872 11713 25881 11747
rect 25881 11713 25915 11747
rect 25915 11713 25924 11747
rect 25872 11704 25924 11713
rect 25228 11636 25280 11688
rect 26056 11704 26108 11756
rect 26424 11704 26476 11756
rect 28540 11704 28592 11756
rect 29736 11704 29788 11756
rect 31392 11704 31444 11756
rect 31852 11772 31904 11824
rect 32588 11772 32640 11824
rect 32496 11747 32548 11756
rect 29184 11679 29236 11688
rect 29184 11645 29193 11679
rect 29193 11645 29227 11679
rect 29227 11645 29236 11679
rect 29184 11636 29236 11645
rect 30564 11679 30616 11688
rect 30564 11645 30573 11679
rect 30573 11645 30607 11679
rect 30607 11645 30616 11679
rect 30564 11636 30616 11645
rect 32496 11713 32505 11747
rect 32505 11713 32539 11747
rect 32539 11713 32548 11747
rect 32496 11704 32548 11713
rect 29092 11568 29144 11620
rect 23572 11500 23624 11552
rect 25412 11500 25464 11552
rect 27988 11500 28040 11552
rect 31484 11500 31536 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 13636 11296 13688 11348
rect 19432 11296 19484 11348
rect 21364 11296 21416 11348
rect 32588 11339 32640 11348
rect 32588 11305 32597 11339
rect 32597 11305 32631 11339
rect 32631 11305 32640 11339
rect 32588 11296 32640 11305
rect 16396 11228 16448 11280
rect 17224 11228 17276 11280
rect 6644 11160 6696 11212
rect 8760 11160 8812 11212
rect 13268 11160 13320 11212
rect 6184 11135 6236 11144
rect 6184 11101 6193 11135
rect 6193 11101 6227 11135
rect 6227 11101 6236 11135
rect 6184 11092 6236 11101
rect 5724 11067 5776 11076
rect 5724 11033 5733 11067
rect 5733 11033 5767 11067
rect 5767 11033 5776 11067
rect 5724 11024 5776 11033
rect 7564 11092 7616 11144
rect 9404 11135 9456 11144
rect 9404 11101 9438 11135
rect 9438 11101 9456 11135
rect 9404 11092 9456 11101
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 20996 11160 21048 11212
rect 31484 11203 31536 11212
rect 22008 11135 22060 11144
rect 22008 11101 22017 11135
rect 22017 11101 22051 11135
rect 22051 11101 22060 11135
rect 22008 11092 22060 11101
rect 31484 11169 31493 11203
rect 31493 11169 31527 11203
rect 31527 11169 31536 11203
rect 31484 11160 31536 11169
rect 29920 11092 29972 11144
rect 6552 11067 6604 11076
rect 6552 11033 6561 11067
rect 6561 11033 6595 11067
rect 6595 11033 6604 11067
rect 6552 11024 6604 11033
rect 5448 10999 5500 11008
rect 5448 10965 5457 10999
rect 5457 10965 5491 10999
rect 5491 10965 5500 10999
rect 5448 10956 5500 10965
rect 6460 10956 6512 11008
rect 10508 10999 10560 11008
rect 10508 10965 10517 10999
rect 10517 10965 10551 10999
rect 10551 10965 10560 10999
rect 10508 10956 10560 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 5724 10752 5776 10804
rect 10508 10752 10560 10804
rect 14280 10795 14332 10804
rect 14280 10761 14289 10795
rect 14289 10761 14323 10795
rect 14323 10761 14332 10795
rect 14280 10752 14332 10761
rect 29184 10752 29236 10804
rect 29920 10795 29972 10804
rect 29920 10761 29929 10795
rect 29929 10761 29963 10795
rect 29963 10761 29972 10795
rect 29920 10752 29972 10761
rect 9220 10684 9272 10736
rect 12992 10727 13044 10736
rect 12992 10693 13001 10727
rect 13001 10693 13035 10727
rect 13035 10693 13044 10727
rect 12992 10684 13044 10693
rect 18236 10727 18288 10736
rect 18236 10693 18245 10727
rect 18245 10693 18279 10727
rect 18279 10693 18288 10727
rect 18236 10684 18288 10693
rect 32128 10684 32180 10736
rect 4712 10616 4764 10668
rect 5172 10616 5224 10668
rect 5264 10616 5316 10668
rect 9128 10616 9180 10668
rect 10048 10659 10100 10668
rect 10048 10625 10057 10659
rect 10057 10625 10091 10659
rect 10091 10625 10100 10659
rect 10048 10616 10100 10625
rect 10416 10616 10468 10668
rect 10968 10616 11020 10668
rect 9772 10548 9824 10600
rect 19984 10591 20036 10600
rect 19984 10557 19993 10591
rect 19993 10557 20027 10591
rect 20027 10557 20036 10591
rect 19984 10548 20036 10557
rect 11152 10412 11204 10464
rect 26424 10412 26476 10464
rect 31116 10412 31168 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 5448 10208 5500 10260
rect 10048 10208 10100 10260
rect 22008 10208 22060 10260
rect 26700 10251 26752 10260
rect 3976 10115 4028 10124
rect 3976 10081 3985 10115
rect 3985 10081 4019 10115
rect 4019 10081 4028 10115
rect 3976 10072 4028 10081
rect 9128 10115 9180 10124
rect 9128 10081 9137 10115
rect 9137 10081 9171 10115
rect 9171 10081 9180 10115
rect 9128 10072 9180 10081
rect 19340 10072 19392 10124
rect 19248 10004 19300 10056
rect 21180 10072 21232 10124
rect 26700 10217 26709 10251
rect 26709 10217 26743 10251
rect 26743 10217 26752 10251
rect 26700 10208 26752 10217
rect 27988 10251 28040 10260
rect 27988 10217 27997 10251
rect 27997 10217 28031 10251
rect 28031 10217 28040 10251
rect 27988 10208 28040 10217
rect 4712 9936 4764 9988
rect 9220 9936 9272 9988
rect 9404 9979 9456 9988
rect 9404 9945 9416 9979
rect 9416 9945 9456 9979
rect 9404 9936 9456 9945
rect 19432 9911 19484 9920
rect 19432 9877 19441 9911
rect 19441 9877 19475 9911
rect 19475 9877 19484 9911
rect 19432 9868 19484 9877
rect 24860 10004 24912 10056
rect 25228 10047 25280 10056
rect 25228 10013 25237 10047
rect 25237 10013 25271 10047
rect 25271 10013 25280 10047
rect 25228 10004 25280 10013
rect 25320 10047 25372 10056
rect 25320 10013 25329 10047
rect 25329 10013 25363 10047
rect 25363 10013 25372 10047
rect 25320 10004 25372 10013
rect 25964 10004 26016 10056
rect 26424 10047 26476 10056
rect 26424 10013 26433 10047
rect 26433 10013 26467 10047
rect 26467 10013 26476 10047
rect 26424 10004 26476 10013
rect 26516 10047 26568 10056
rect 26516 10013 26525 10047
rect 26525 10013 26559 10047
rect 26559 10013 26568 10047
rect 26516 10004 26568 10013
rect 29092 10004 29144 10056
rect 20168 9936 20220 9988
rect 25412 9936 25464 9988
rect 26056 9936 26108 9988
rect 21180 9868 21232 9920
rect 24860 9911 24912 9920
rect 24860 9877 24869 9911
rect 24869 9877 24903 9911
rect 24903 9877 24912 9911
rect 24860 9868 24912 9877
rect 27620 9936 27672 9988
rect 28264 9936 28316 9988
rect 29000 9936 29052 9988
rect 30196 10047 30248 10056
rect 30196 10013 30205 10047
rect 30205 10013 30239 10047
rect 30239 10013 30248 10047
rect 30196 10004 30248 10013
rect 30472 10004 30524 10056
rect 30288 9936 30340 9988
rect 29644 9868 29696 9920
rect 30656 9911 30708 9920
rect 30656 9877 30665 9911
rect 30665 9877 30699 9911
rect 30699 9877 30708 9911
rect 30656 9868 30708 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 11152 9664 11204 9716
rect 17224 9664 17276 9716
rect 20168 9664 20220 9716
rect 20536 9664 20588 9716
rect 15568 9639 15620 9648
rect 15568 9605 15577 9639
rect 15577 9605 15611 9639
rect 15611 9605 15620 9639
rect 15568 9596 15620 9605
rect 19432 9596 19484 9648
rect 20444 9596 20496 9648
rect 29092 9664 29144 9716
rect 25412 9639 25464 9648
rect 25412 9605 25421 9639
rect 25421 9605 25455 9639
rect 25455 9605 25464 9639
rect 25412 9596 25464 9605
rect 27712 9596 27764 9648
rect 2964 9528 3016 9580
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 15292 9528 15344 9580
rect 15476 9528 15528 9580
rect 16488 9528 16540 9580
rect 19248 9528 19300 9580
rect 20536 9571 20588 9580
rect 20536 9537 20545 9571
rect 20545 9537 20579 9571
rect 20579 9537 20588 9571
rect 20536 9528 20588 9537
rect 1860 9324 1912 9376
rect 14280 9367 14332 9376
rect 14280 9333 14289 9367
rect 14289 9333 14323 9367
rect 14323 9333 14332 9367
rect 14280 9324 14332 9333
rect 15200 9367 15252 9376
rect 15200 9333 15209 9367
rect 15209 9333 15243 9367
rect 15243 9333 15252 9367
rect 15200 9324 15252 9333
rect 20904 9571 20956 9580
rect 20904 9537 20913 9571
rect 20913 9537 20947 9571
rect 20947 9537 20956 9571
rect 20904 9528 20956 9537
rect 26516 9528 26568 9580
rect 29000 9596 29052 9648
rect 29644 9639 29696 9648
rect 29644 9605 29653 9639
rect 29653 9605 29687 9639
rect 29687 9605 29696 9639
rect 29644 9596 29696 9605
rect 26148 9460 26200 9512
rect 20812 9392 20864 9444
rect 21088 9435 21140 9444
rect 21088 9401 21097 9435
rect 21097 9401 21131 9435
rect 21131 9401 21140 9435
rect 21088 9392 21140 9401
rect 19340 9324 19392 9376
rect 20260 9324 20312 9376
rect 28816 9392 28868 9444
rect 29736 9324 29788 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2964 9120 3016 9172
rect 4068 9120 4120 9172
rect 16396 9120 16448 9172
rect 16488 9052 16540 9104
rect 18604 9120 18656 9172
rect 18972 9120 19024 9172
rect 20444 9120 20496 9172
rect 23572 9163 23624 9172
rect 23572 9129 23581 9163
rect 23581 9129 23615 9163
rect 23615 9129 23624 9163
rect 23572 9120 23624 9129
rect 25228 9120 25280 9172
rect 27712 9120 27764 9172
rect 30932 9120 30984 9172
rect 31116 9163 31168 9172
rect 31116 9129 31125 9163
rect 31125 9129 31159 9163
rect 31159 9129 31168 9163
rect 31116 9120 31168 9129
rect 1860 9027 1912 9036
rect 1860 8993 1869 9027
rect 1869 8993 1903 9027
rect 1903 8993 1912 9027
rect 1860 8984 1912 8993
rect 14280 9027 14332 9036
rect 14280 8993 14289 9027
rect 14289 8993 14323 9027
rect 14323 8993 14332 9027
rect 14280 8984 14332 8993
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 2964 8916 3016 8968
rect 16304 8959 16356 8968
rect 16304 8925 16313 8959
rect 16313 8925 16347 8959
rect 16347 8925 16356 8959
rect 16304 8916 16356 8925
rect 16396 8916 16448 8968
rect 18880 8984 18932 9036
rect 18236 8916 18288 8968
rect 18512 8959 18564 8968
rect 18512 8925 18521 8959
rect 18521 8925 18555 8959
rect 18555 8925 18564 8959
rect 18512 8916 18564 8925
rect 18604 8916 18656 8968
rect 21916 8916 21968 8968
rect 18328 8891 18380 8900
rect 18328 8857 18337 8891
rect 18337 8857 18371 8891
rect 18371 8857 18380 8891
rect 18328 8848 18380 8857
rect 19432 8891 19484 8900
rect 2780 8780 2832 8832
rect 5632 8780 5684 8832
rect 6736 8780 6788 8832
rect 16672 8780 16724 8832
rect 19432 8857 19441 8891
rect 19441 8857 19475 8891
rect 19475 8857 19484 8891
rect 19432 8848 19484 8857
rect 19984 8848 20036 8900
rect 22192 8848 22244 8900
rect 23388 8891 23440 8900
rect 23388 8857 23397 8891
rect 23397 8857 23431 8891
rect 23431 8857 23440 8891
rect 23388 8848 23440 8857
rect 24584 8959 24636 8968
rect 24584 8925 24593 8959
rect 24593 8925 24627 8959
rect 24627 8925 24636 8959
rect 24584 8916 24636 8925
rect 24860 8959 24912 8968
rect 24860 8925 24894 8959
rect 24894 8925 24912 8959
rect 24860 8916 24912 8925
rect 29092 8916 29144 8968
rect 29736 8959 29788 8968
rect 29736 8925 29745 8959
rect 29745 8925 29779 8959
rect 29779 8925 29788 8959
rect 29736 8916 29788 8925
rect 25412 8848 25464 8900
rect 29644 8848 29696 8900
rect 29828 8848 29880 8900
rect 20076 8780 20128 8832
rect 21640 8823 21692 8832
rect 21640 8789 21649 8823
rect 21649 8789 21683 8823
rect 21683 8789 21692 8823
rect 21640 8780 21692 8789
rect 22008 8823 22060 8832
rect 22008 8789 22017 8823
rect 22017 8789 22051 8823
rect 22051 8789 22060 8823
rect 22008 8780 22060 8789
rect 24676 8780 24728 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1584 8576 1636 8628
rect 5540 8576 5592 8628
rect 2964 8551 3016 8560
rect 2964 8517 2973 8551
rect 2973 8517 3007 8551
rect 3007 8517 3016 8551
rect 2964 8508 3016 8517
rect 5356 8508 5408 8560
rect 2780 8483 2832 8492
rect 2780 8449 2789 8483
rect 2789 8449 2823 8483
rect 2823 8449 2832 8483
rect 4620 8483 4672 8492
rect 2780 8440 2832 8449
rect 4620 8449 4629 8483
rect 4629 8449 4663 8483
rect 4663 8449 4672 8483
rect 4620 8440 4672 8449
rect 5448 8440 5500 8492
rect 15752 8576 15804 8628
rect 18236 8576 18288 8628
rect 19432 8576 19484 8628
rect 20352 8576 20404 8628
rect 22008 8576 22060 8628
rect 23388 8576 23440 8628
rect 29644 8576 29696 8628
rect 30932 8619 30984 8628
rect 30932 8585 30941 8619
rect 30941 8585 30975 8619
rect 30975 8585 30984 8619
rect 30932 8576 30984 8585
rect 12716 8508 12768 8560
rect 6736 8483 6788 8492
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 10876 8440 10928 8492
rect 13452 8440 13504 8492
rect 14740 8440 14792 8492
rect 8300 8372 8352 8424
rect 10232 8372 10284 8424
rect 10600 8415 10652 8424
rect 10600 8381 10609 8415
rect 10609 8381 10643 8415
rect 10643 8381 10652 8415
rect 10600 8372 10652 8381
rect 14648 8372 14700 8424
rect 15108 8508 15160 8560
rect 17868 8508 17920 8560
rect 18420 8508 18472 8560
rect 14924 8440 14976 8492
rect 19340 8440 19392 8492
rect 21640 8508 21692 8560
rect 20904 8440 20956 8492
rect 24492 8508 24544 8560
rect 24676 8551 24728 8560
rect 24676 8517 24685 8551
rect 24685 8517 24719 8551
rect 24719 8517 24728 8551
rect 24676 8508 24728 8517
rect 22928 8440 22980 8492
rect 29092 8508 29144 8560
rect 29920 8508 29972 8560
rect 30196 8508 30248 8560
rect 30656 8440 30708 8492
rect 30748 8483 30800 8492
rect 30748 8449 30757 8483
rect 30757 8449 30791 8483
rect 30791 8449 30800 8483
rect 30748 8440 30800 8449
rect 15292 8372 15344 8424
rect 16488 8372 16540 8424
rect 32496 8372 32548 8424
rect 7012 8304 7064 8356
rect 10140 8304 10192 8356
rect 12992 8304 13044 8356
rect 16304 8304 16356 8356
rect 6552 8236 6604 8288
rect 12624 8236 12676 8288
rect 18512 8279 18564 8288
rect 18512 8245 18521 8279
rect 18521 8245 18555 8279
rect 18555 8245 18564 8279
rect 18512 8236 18564 8245
rect 30288 8304 30340 8356
rect 20628 8236 20680 8288
rect 20720 8236 20772 8288
rect 23112 8236 23164 8288
rect 23204 8236 23256 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 6920 8075 6972 8084
rect 6920 8041 6929 8075
rect 6929 8041 6963 8075
rect 6963 8041 6972 8075
rect 6920 8032 6972 8041
rect 8300 8032 8352 8084
rect 10876 8075 10928 8084
rect 10876 8041 10885 8075
rect 10885 8041 10919 8075
rect 10919 8041 10928 8075
rect 10876 8032 10928 8041
rect 8944 7896 8996 7948
rect 9496 7896 9548 7948
rect 12716 8032 12768 8084
rect 15108 8032 15160 8084
rect 15568 8032 15620 8084
rect 18512 8032 18564 8084
rect 20812 8075 20864 8084
rect 16488 7964 16540 8016
rect 20812 8041 20821 8075
rect 20821 8041 20855 8075
rect 20855 8041 20864 8075
rect 20812 8032 20864 8041
rect 22928 8032 22980 8084
rect 23112 8032 23164 8084
rect 23572 8032 23624 8084
rect 26148 8032 26200 8084
rect 29828 8032 29880 8084
rect 20720 7964 20772 8016
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 6552 7828 6604 7880
rect 14280 7896 14332 7948
rect 4620 7760 4672 7812
rect 5356 7760 5408 7812
rect 6736 7692 6788 7744
rect 15200 7828 15252 7880
rect 15476 7828 15528 7880
rect 16672 7871 16724 7880
rect 16672 7837 16681 7871
rect 16681 7837 16715 7871
rect 16715 7837 16724 7871
rect 16672 7828 16724 7837
rect 19248 7828 19300 7880
rect 19432 7871 19484 7880
rect 19432 7837 19441 7871
rect 19441 7837 19475 7871
rect 19475 7837 19484 7871
rect 19432 7828 19484 7837
rect 20628 7828 20680 7880
rect 16304 7735 16356 7744
rect 16304 7701 16313 7735
rect 16313 7701 16347 7735
rect 16347 7701 16356 7735
rect 16304 7692 16356 7701
rect 18420 7735 18472 7744
rect 18420 7701 18429 7735
rect 18429 7701 18463 7735
rect 18463 7701 18472 7735
rect 18420 7692 18472 7701
rect 18880 7692 18932 7744
rect 20444 7760 20496 7812
rect 20536 7760 20588 7812
rect 23204 7803 23256 7812
rect 23204 7769 23213 7803
rect 23213 7769 23247 7803
rect 23247 7769 23256 7803
rect 23204 7760 23256 7769
rect 20904 7692 20956 7744
rect 24676 7828 24728 7880
rect 27436 7828 27488 7880
rect 31392 7896 31444 7948
rect 30196 7871 30248 7880
rect 30196 7837 30205 7871
rect 30205 7837 30239 7871
rect 30239 7837 30248 7871
rect 30196 7828 30248 7837
rect 25596 7760 25648 7812
rect 31116 7760 31168 7812
rect 25320 7692 25372 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 7012 7531 7064 7540
rect 7012 7497 7021 7531
rect 7021 7497 7055 7531
rect 7055 7497 7064 7531
rect 7012 7488 7064 7497
rect 6920 7463 6972 7472
rect 6920 7429 6929 7463
rect 6929 7429 6963 7463
rect 6963 7429 6972 7463
rect 6920 7420 6972 7429
rect 10416 7488 10468 7540
rect 9588 7395 9640 7404
rect 9588 7361 9611 7395
rect 9611 7361 9640 7395
rect 9588 7352 9640 7361
rect 15292 7488 15344 7540
rect 15752 7531 15804 7540
rect 15752 7497 15761 7531
rect 15761 7497 15795 7531
rect 15795 7497 15804 7531
rect 15752 7488 15804 7497
rect 18052 7488 18104 7540
rect 19340 7488 19392 7540
rect 20444 7531 20496 7540
rect 20444 7497 20453 7531
rect 20453 7497 20487 7531
rect 20487 7497 20496 7531
rect 20444 7488 20496 7497
rect 20812 7531 20864 7540
rect 20812 7497 20821 7531
rect 20821 7497 20855 7531
rect 20855 7497 20864 7531
rect 20812 7488 20864 7497
rect 24584 7488 24636 7540
rect 25596 7531 25648 7540
rect 25596 7497 25605 7531
rect 25605 7497 25639 7531
rect 25639 7497 25648 7531
rect 25596 7488 25648 7497
rect 26148 7488 26200 7540
rect 29736 7488 29788 7540
rect 14648 7463 14700 7472
rect 14648 7429 14682 7463
rect 14682 7429 14700 7463
rect 14648 7420 14700 7429
rect 20076 7420 20128 7472
rect 23388 7463 23440 7472
rect 23388 7429 23397 7463
rect 23397 7429 23431 7463
rect 23431 7429 23440 7463
rect 23388 7420 23440 7429
rect 25320 7420 25372 7472
rect 25688 7420 25740 7472
rect 12624 7352 12676 7404
rect 14464 7352 14516 7404
rect 19340 7352 19392 7404
rect 20628 7395 20680 7404
rect 20628 7361 20637 7395
rect 20637 7361 20671 7395
rect 20671 7361 20680 7395
rect 20628 7352 20680 7361
rect 20904 7395 20956 7404
rect 20904 7361 20913 7395
rect 20913 7361 20947 7395
rect 20947 7361 20956 7395
rect 20904 7352 20956 7361
rect 28816 7420 28868 7472
rect 5448 7216 5500 7268
rect 8300 7216 8352 7268
rect 30748 7284 30800 7336
rect 6552 7191 6604 7200
rect 6552 7157 6561 7191
rect 6561 7157 6595 7191
rect 6595 7157 6604 7191
rect 6552 7148 6604 7157
rect 10692 7191 10744 7200
rect 10692 7157 10701 7191
rect 10701 7157 10735 7191
rect 10735 7157 10744 7191
rect 10692 7148 10744 7157
rect 12164 7191 12216 7200
rect 12164 7157 12173 7191
rect 12173 7157 12207 7191
rect 12207 7157 12216 7191
rect 12164 7148 12216 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 10416 6876 10468 6928
rect 6092 6808 6144 6860
rect 7012 6851 7064 6860
rect 7012 6817 7021 6851
rect 7021 6817 7055 6851
rect 7055 6817 7064 6851
rect 7012 6808 7064 6817
rect 10692 6808 10744 6860
rect 6552 6740 6604 6792
rect 10876 6783 10928 6792
rect 10876 6749 10885 6783
rect 10885 6749 10919 6783
rect 10919 6749 10928 6783
rect 10876 6740 10928 6749
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 16304 6740 16356 6792
rect 24676 6740 24728 6792
rect 25320 6672 25372 6724
rect 6644 6604 6696 6656
rect 10508 6647 10560 6656
rect 10508 6613 10517 6647
rect 10517 6613 10551 6647
rect 10551 6613 10560 6647
rect 10508 6604 10560 6613
rect 16672 6604 16724 6656
rect 25964 6647 26016 6656
rect 25964 6613 25973 6647
rect 25973 6613 26007 6647
rect 26007 6613 26016 6647
rect 25964 6604 26016 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 12164 6443 12216 6452
rect 12164 6409 12173 6443
rect 12173 6409 12207 6443
rect 12207 6409 12216 6443
rect 12164 6400 12216 6409
rect 18880 6400 18932 6452
rect 25320 6443 25372 6452
rect 25320 6409 25329 6443
rect 25329 6409 25363 6443
rect 25363 6409 25372 6443
rect 25320 6400 25372 6409
rect 25964 6400 26016 6452
rect 10508 6332 10560 6384
rect 18420 6332 18472 6384
rect 27436 6332 27488 6384
rect 25688 6264 25740 6316
rect 12256 6239 12308 6248
rect 12256 6205 12265 6239
rect 12265 6205 12299 6239
rect 12299 6205 12308 6239
rect 12256 6196 12308 6205
rect 11704 6103 11756 6112
rect 11704 6069 11713 6103
rect 11713 6069 11747 6103
rect 11747 6069 11756 6103
rect 11704 6060 11756 6069
rect 19432 6060 19484 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 7012 5856 7064 5908
rect 11704 5856 11756 5908
rect 21916 5856 21968 5908
rect 4620 5763 4672 5772
rect 4620 5729 4629 5763
rect 4629 5729 4663 5763
rect 4663 5729 4672 5763
rect 4620 5720 4672 5729
rect 5724 5584 5776 5636
rect 27528 5720 27580 5772
rect 10324 5652 10376 5704
rect 12256 5652 12308 5704
rect 28080 5627 28132 5636
rect 28080 5593 28114 5627
rect 28114 5593 28132 5627
rect 28080 5584 28132 5593
rect 9772 5516 9824 5568
rect 28632 5516 28684 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 10140 5355 10192 5364
rect 10140 5321 10149 5355
rect 10149 5321 10183 5355
rect 10183 5321 10192 5355
rect 10140 5312 10192 5321
rect 14464 5355 14516 5364
rect 14464 5321 14473 5355
rect 14473 5321 14507 5355
rect 14507 5321 14516 5355
rect 14464 5312 14516 5321
rect 19432 5312 19484 5364
rect 24676 5355 24728 5364
rect 24676 5321 24685 5355
rect 24685 5321 24719 5355
rect 24719 5321 24728 5355
rect 24676 5312 24728 5321
rect 29920 5355 29972 5364
rect 29920 5321 29929 5355
rect 29929 5321 29963 5355
rect 29963 5321 29972 5355
rect 29920 5312 29972 5321
rect 5540 5244 5592 5296
rect 5724 5287 5776 5296
rect 5724 5253 5733 5287
rect 5733 5253 5767 5287
rect 5767 5253 5776 5287
rect 5724 5244 5776 5253
rect 12992 5287 13044 5296
rect 12992 5253 13001 5287
rect 13001 5253 13035 5287
rect 13035 5253 13044 5287
rect 12992 5244 13044 5253
rect 19340 5244 19392 5296
rect 23388 5287 23440 5296
rect 23388 5253 23397 5287
rect 23397 5253 23431 5287
rect 23431 5253 23440 5287
rect 23388 5244 23440 5253
rect 28816 5244 28868 5296
rect 5632 5219 5684 5228
rect 5632 5185 5641 5219
rect 5641 5185 5675 5219
rect 5675 5185 5684 5219
rect 5632 5176 5684 5185
rect 9956 5219 10008 5228
rect 9956 5185 9965 5219
rect 9965 5185 9999 5219
rect 9999 5185 10008 5219
rect 9956 5176 10008 5185
rect 8208 5108 8260 5160
rect 17868 5176 17920 5228
rect 22192 5176 22244 5228
rect 22100 4972 22152 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 10416 4768 10468 4820
rect 12716 4768 12768 4820
rect 5632 4632 5684 4684
rect 9772 4700 9824 4752
rect 5540 4564 5592 4616
rect 6368 4607 6420 4616
rect 6368 4573 6377 4607
rect 6377 4573 6411 4607
rect 6411 4573 6420 4607
rect 6368 4564 6420 4573
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 8208 4607 8260 4616
rect 6552 4564 6604 4573
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 10324 4607 10376 4616
rect 10324 4573 10333 4607
rect 10333 4573 10367 4607
rect 10367 4573 10376 4607
rect 10324 4564 10376 4573
rect 10508 4564 10560 4616
rect 10692 4564 10744 4616
rect 12716 4607 12768 4616
rect 6920 4496 6972 4548
rect 7932 4496 7984 4548
rect 10232 4496 10284 4548
rect 12716 4573 12725 4607
rect 12725 4573 12759 4607
rect 12759 4573 12768 4607
rect 12716 4564 12768 4573
rect 17500 4768 17552 4820
rect 22284 4700 22336 4752
rect 28632 4743 28684 4752
rect 28632 4709 28641 4743
rect 28641 4709 28675 4743
rect 28675 4709 28684 4743
rect 28632 4700 28684 4709
rect 28724 4743 28776 4752
rect 28724 4709 28733 4743
rect 28733 4709 28767 4743
rect 28767 4709 28776 4743
rect 28724 4700 28776 4709
rect 15108 4564 15160 4616
rect 17868 4564 17920 4616
rect 21916 4607 21968 4616
rect 21916 4573 21925 4607
rect 21925 4573 21959 4607
rect 21959 4573 21968 4607
rect 21916 4564 21968 4573
rect 28816 4675 28868 4684
rect 28816 4641 28825 4675
rect 28825 4641 28859 4675
rect 28859 4641 28868 4675
rect 28816 4632 28868 4641
rect 23204 4607 23256 4616
rect 23204 4573 23213 4607
rect 23213 4573 23247 4607
rect 23247 4573 23256 4607
rect 23204 4564 23256 4573
rect 27160 4564 27212 4616
rect 27528 4564 27580 4616
rect 9128 4471 9180 4480
rect 9128 4437 9137 4471
rect 9137 4437 9171 4471
rect 9171 4437 9180 4471
rect 9128 4428 9180 4437
rect 12624 4428 12676 4480
rect 26792 4496 26844 4548
rect 14556 4428 14608 4480
rect 17684 4428 17736 4480
rect 19432 4428 19484 4480
rect 22652 4428 22704 4480
rect 22836 4428 22888 4480
rect 23572 4428 23624 4480
rect 23848 4428 23900 4480
rect 27804 4471 27856 4480
rect 27804 4437 27813 4471
rect 27813 4437 27847 4471
rect 27847 4437 27856 4471
rect 27804 4428 27856 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 7932 4267 7984 4276
rect 7932 4233 7941 4267
rect 7941 4233 7975 4267
rect 7975 4233 7984 4267
rect 7932 4224 7984 4233
rect 9956 4224 10008 4276
rect 10692 4267 10744 4276
rect 10692 4233 10701 4267
rect 10701 4233 10735 4267
rect 10735 4233 10744 4267
rect 10692 4224 10744 4233
rect 17868 4224 17920 4276
rect 22652 4224 22704 4276
rect 23020 4224 23072 4276
rect 28816 4224 28868 4276
rect 10232 4156 10284 4208
rect 4712 4088 4764 4140
rect 5908 4088 5960 4140
rect 8944 4131 8996 4140
rect 8944 4097 8953 4131
rect 8953 4097 8987 4131
rect 8987 4097 8996 4131
rect 8944 4088 8996 4097
rect 12624 4131 12676 4140
rect 12624 4097 12633 4131
rect 12633 4097 12667 4131
rect 12667 4097 12676 4131
rect 12624 4088 12676 4097
rect 14096 4088 14148 4140
rect 14556 4088 14608 4140
rect 14740 4131 14792 4140
rect 14740 4097 14774 4131
rect 14774 4097 14792 4131
rect 22284 4199 22336 4208
rect 22284 4165 22318 4199
rect 22318 4165 22336 4199
rect 22284 4156 22336 4165
rect 14740 4088 14792 4097
rect 17684 4131 17736 4140
rect 17684 4097 17693 4131
rect 17693 4097 17727 4131
rect 17727 4097 17736 4131
rect 17684 4088 17736 4097
rect 18420 4088 18472 4140
rect 19432 4088 19484 4140
rect 19800 4131 19852 4140
rect 19800 4097 19834 4131
rect 19834 4097 19852 4131
rect 19800 4088 19852 4097
rect 22100 4088 22152 4140
rect 23848 4131 23900 4140
rect 23848 4097 23857 4131
rect 23857 4097 23891 4131
rect 23891 4097 23900 4131
rect 23848 4088 23900 4097
rect 24584 4088 24636 4140
rect 27160 4131 27212 4140
rect 27160 4097 27169 4131
rect 27169 4097 27203 4131
rect 27203 4097 27212 4131
rect 27160 4088 27212 4097
rect 9220 4063 9272 4072
rect 9220 4029 9229 4063
rect 9229 4029 9263 4063
rect 9263 4029 9272 4063
rect 9220 4020 9272 4029
rect 26424 4020 26476 4072
rect 29092 4088 29144 4140
rect 17132 3952 17184 4004
rect 8300 3884 8352 3936
rect 14464 3884 14516 3936
rect 16580 3884 16632 3936
rect 19340 3884 19392 3936
rect 20904 3927 20956 3936
rect 20904 3893 20913 3927
rect 20913 3893 20947 3927
rect 20947 3893 20956 3927
rect 20904 3884 20956 3893
rect 25044 3884 25096 3936
rect 27436 3884 27488 3936
rect 28724 3884 28776 3936
rect 32312 3884 32364 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 6644 3680 6696 3732
rect 8208 3680 8260 3732
rect 10508 3680 10560 3732
rect 14740 3680 14792 3732
rect 19800 3723 19852 3732
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 9128 3544 9180 3596
rect 8300 3476 8352 3528
rect 15108 3544 15160 3596
rect 16580 3587 16632 3596
rect 16580 3553 16589 3587
rect 16589 3553 16623 3587
rect 16623 3553 16632 3587
rect 16580 3544 16632 3553
rect 19800 3689 19809 3723
rect 19809 3689 19843 3723
rect 19843 3689 19852 3723
rect 19800 3680 19852 3689
rect 19064 3544 19116 3596
rect 23204 3680 23256 3732
rect 23572 3680 23624 3732
rect 23756 3680 23808 3732
rect 24584 3723 24636 3732
rect 24584 3689 24593 3723
rect 24593 3689 24627 3723
rect 24627 3689 24636 3723
rect 24584 3680 24636 3689
rect 26792 3723 26844 3732
rect 26792 3689 26801 3723
rect 26801 3689 26835 3723
rect 26835 3689 26844 3723
rect 26792 3680 26844 3689
rect 27436 3680 27488 3732
rect 27804 3680 27856 3732
rect 28632 3680 28684 3732
rect 29092 3723 29144 3732
rect 29092 3689 29101 3723
rect 29101 3689 29135 3723
rect 29135 3689 29144 3723
rect 29092 3680 29144 3689
rect 25044 3587 25096 3596
rect 25044 3553 25053 3587
rect 25053 3553 25087 3587
rect 25087 3553 25096 3587
rect 25044 3544 25096 3553
rect 6920 3408 6972 3460
rect 9220 3408 9272 3460
rect 11060 3408 11112 3460
rect 16856 3451 16908 3460
rect 16856 3417 16890 3451
rect 16890 3417 16908 3451
rect 20904 3476 20956 3528
rect 22560 3519 22612 3528
rect 22560 3485 22569 3519
rect 22569 3485 22603 3519
rect 22603 3485 22612 3519
rect 22560 3476 22612 3485
rect 22836 3519 22888 3528
rect 22836 3485 22870 3519
rect 22870 3485 22888 3519
rect 22836 3476 22888 3485
rect 23204 3476 23256 3528
rect 16856 3408 16908 3417
rect 8944 3340 8996 3392
rect 17132 3340 17184 3392
rect 17960 3383 18012 3392
rect 17960 3349 17969 3383
rect 17969 3349 18003 3383
rect 18003 3349 18012 3383
rect 17960 3340 18012 3349
rect 28724 3612 28776 3664
rect 28908 3655 28960 3664
rect 28908 3621 28917 3655
rect 28917 3621 28951 3655
rect 28951 3621 28960 3655
rect 28908 3612 28960 3621
rect 27896 3544 27948 3596
rect 28816 3544 28868 3596
rect 28908 3476 28960 3528
rect 26424 3451 26476 3460
rect 26424 3417 26433 3451
rect 26433 3417 26467 3451
rect 26467 3417 26476 3451
rect 26424 3408 26476 3417
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 10140 3136 10192 3188
rect 12716 3136 12768 3188
rect 14096 3179 14148 3188
rect 14096 3145 14105 3179
rect 14105 3145 14139 3179
rect 14139 3145 14148 3179
rect 14096 3136 14148 3145
rect 14464 3136 14516 3188
rect 15660 3136 15712 3188
rect 16856 3179 16908 3188
rect 16856 3145 16865 3179
rect 16865 3145 16899 3179
rect 16899 3145 16908 3179
rect 16856 3136 16908 3145
rect 17224 3179 17276 3188
rect 17224 3145 17233 3179
rect 17233 3145 17267 3179
rect 17267 3145 17276 3179
rect 17224 3136 17276 3145
rect 17960 3136 18012 3188
rect 18420 3179 18472 3188
rect 18420 3145 18429 3179
rect 18429 3145 18463 3179
rect 18463 3145 18472 3179
rect 18420 3136 18472 3145
rect 22560 3136 22612 3188
rect 28080 3136 28132 3188
rect 8484 3068 8536 3120
rect 6368 3000 6420 3052
rect 9956 3000 10008 3052
rect 18788 3043 18840 3052
rect 848 2932 900 2984
rect 6552 2932 6604 2984
rect 18788 3009 18797 3043
rect 18797 3009 18831 3043
rect 18831 3009 18840 3043
rect 18788 3000 18840 3009
rect 19340 3000 19392 3052
rect 20076 3000 20128 3052
rect 22192 3000 22244 3052
rect 10232 2975 10284 2984
rect 10232 2941 10241 2975
rect 10241 2941 10275 2975
rect 10275 2941 10284 2975
rect 10232 2932 10284 2941
rect 15108 2932 15160 2984
rect 19064 2975 19116 2984
rect 19064 2941 19073 2975
rect 19073 2941 19107 2975
rect 19107 2941 19116 2975
rect 19064 2932 19116 2941
rect 9680 2864 9732 2916
rect 26424 2864 26476 2916
rect 39120 2932 39172 2984
rect 27896 2907 27948 2916
rect 27896 2873 27905 2907
rect 27905 2873 27939 2907
rect 27939 2873 27948 2907
rect 27896 2864 27948 2873
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 6368 2592 6420 2644
rect 18788 2592 18840 2644
rect 11060 2524 11112 2576
rect 11152 2524 11204 2576
rect 28908 2456 28960 2508
rect 6368 2388 6420 2440
rect 6736 2388 6788 2440
rect 8208 2388 8260 2440
rect 9680 2388 9732 2440
rect 11152 2388 11204 2440
rect 12624 2388 12676 2440
rect 14096 2388 14148 2440
rect 15660 2431 15712 2440
rect 15660 2397 15669 2431
rect 15669 2397 15703 2431
rect 15703 2397 15712 2431
rect 15660 2388 15712 2397
rect 17132 2431 17184 2440
rect 17132 2397 17141 2431
rect 17141 2397 17175 2431
rect 17175 2397 17184 2431
rect 17132 2388 17184 2397
rect 17960 2388 18012 2440
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 20904 2388 20956 2440
rect 23020 2431 23072 2440
rect 23020 2397 23029 2431
rect 23029 2397 23063 2431
rect 23063 2397 23072 2431
rect 23020 2388 23072 2397
rect 23756 2388 23808 2440
rect 25044 2388 25096 2440
rect 27436 2431 27488 2440
rect 27436 2397 27445 2431
rect 27445 2397 27479 2431
rect 27479 2397 27488 2431
rect 27436 2388 27488 2397
rect 27896 2388 27948 2440
rect 32312 2431 32364 2440
rect 32312 2397 32321 2431
rect 32321 2397 32355 2431
rect 32355 2397 32364 2431
rect 32312 2388 32364 2397
rect 33232 2388 33284 2440
rect 34704 2388 34756 2440
rect 36176 2388 36228 2440
rect 37648 2388 37700 2440
rect 2320 2320 2372 2372
rect 3792 2320 3844 2372
rect 5264 2320 5316 2372
rect 15568 2320 15620 2372
rect 17040 2320 17092 2372
rect 18512 2320 18564 2372
rect 19984 2320 20036 2372
rect 21456 2320 21508 2372
rect 22928 2320 22980 2372
rect 24400 2320 24452 2372
rect 25872 2320 25924 2372
rect 27344 2320 27396 2372
rect 28816 2320 28868 2372
rect 30288 2320 30340 2372
rect 31760 2320 31812 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 1412 39222 1716 39250
rect 1412 17746 1440 39222
rect 1688 39114 1716 39222
rect 1766 39200 1822 40000
rect 5078 39200 5134 40000
rect 8390 39200 8446 40000
rect 11702 39200 11758 40000
rect 15014 39200 15070 40000
rect 18326 39200 18382 40000
rect 21638 39200 21694 40000
rect 21744 39222 22048 39250
rect 1780 39114 1808 39200
rect 1688 39086 1808 39114
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 5092 37262 5120 39200
rect 5448 37324 5500 37330
rect 5448 37266 5500 37272
rect 5080 37256 5132 37262
rect 5080 37198 5132 37204
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 5460 31822 5488 37266
rect 8404 37262 8432 39200
rect 11716 37262 11744 39200
rect 14280 37392 14332 37398
rect 14280 37334 14332 37340
rect 14924 37392 14976 37398
rect 14924 37334 14976 37340
rect 13452 37324 13504 37330
rect 13452 37266 13504 37272
rect 8392 37256 8444 37262
rect 8392 37198 8444 37204
rect 11704 37256 11756 37262
rect 11704 37198 11756 37204
rect 13464 36922 13492 37266
rect 13452 36916 13504 36922
rect 13452 36858 13504 36864
rect 13820 36576 13872 36582
rect 13820 36518 13872 36524
rect 5448 31816 5500 31822
rect 5448 31758 5500 31764
rect 13832 31482 13860 36518
rect 14188 36304 14240 36310
rect 14188 36246 14240 36252
rect 14096 35488 14148 35494
rect 14096 35430 14148 35436
rect 13820 31476 13872 31482
rect 13820 31418 13872 31424
rect 6736 31340 6788 31346
rect 6736 31282 6788 31288
rect 12624 31340 12676 31346
rect 12676 31300 12756 31328
rect 12624 31282 12676 31288
rect 5540 31272 5592 31278
rect 5540 31214 5592 31220
rect 5448 31136 5500 31142
rect 5448 31078 5500 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 5264 30796 5316 30802
rect 5264 30738 5316 30744
rect 4620 30728 4672 30734
rect 4620 30670 4672 30676
rect 4632 30394 4660 30670
rect 4620 30388 4672 30394
rect 4620 30330 4672 30336
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4988 29640 5040 29646
rect 5040 29588 5120 29594
rect 4988 29582 5120 29588
rect 5000 29566 5120 29582
rect 5092 29306 5120 29566
rect 5172 29504 5224 29510
rect 5172 29446 5224 29452
rect 5080 29300 5132 29306
rect 5080 29242 5132 29248
rect 4988 29164 5040 29170
rect 4988 29106 5040 29112
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4528 27532 4580 27538
rect 4528 27474 4580 27480
rect 4540 26926 4568 27474
rect 4620 27396 4672 27402
rect 4620 27338 4672 27344
rect 4632 26994 4660 27338
rect 4712 27328 4764 27334
rect 4712 27270 4764 27276
rect 4620 26988 4672 26994
rect 4620 26930 4672 26936
rect 4528 26920 4580 26926
rect 4528 26862 4580 26868
rect 3148 26852 3200 26858
rect 3148 26794 3200 26800
rect 3160 26314 3188 26794
rect 4620 26784 4672 26790
rect 4620 26726 4672 26732
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4632 26450 4660 26726
rect 4620 26444 4672 26450
rect 4620 26386 4672 26392
rect 4724 26382 4752 27270
rect 5000 26382 5028 29106
rect 5092 28150 5120 29242
rect 5184 29238 5212 29446
rect 5172 29232 5224 29238
rect 5172 29174 5224 29180
rect 5080 28144 5132 28150
rect 5080 28086 5132 28092
rect 5184 27878 5212 29174
rect 5276 28966 5304 30738
rect 5460 30326 5488 31078
rect 5448 30320 5500 30326
rect 5448 30262 5500 30268
rect 5356 29708 5408 29714
rect 5356 29650 5408 29656
rect 5368 29034 5396 29650
rect 5552 29646 5580 31214
rect 6000 30660 6052 30666
rect 6000 30602 6052 30608
rect 6012 30190 6040 30602
rect 6748 30326 6776 31282
rect 6828 31204 6880 31210
rect 6828 31146 6880 31152
rect 6736 30320 6788 30326
rect 6736 30262 6788 30268
rect 6840 30258 6868 31146
rect 12072 31136 12124 31142
rect 12072 31078 12124 31084
rect 10324 30796 10376 30802
rect 10324 30738 10376 30744
rect 8484 30728 8536 30734
rect 8484 30670 8536 30676
rect 7104 30320 7156 30326
rect 7104 30262 7156 30268
rect 6368 30252 6420 30258
rect 6368 30194 6420 30200
rect 6460 30252 6512 30258
rect 6460 30194 6512 30200
rect 6828 30252 6880 30258
rect 6828 30194 6880 30200
rect 6000 30184 6052 30190
rect 6000 30126 6052 30132
rect 5724 30048 5776 30054
rect 5724 29990 5776 29996
rect 5540 29640 5592 29646
rect 5540 29582 5592 29588
rect 5448 29504 5500 29510
rect 5448 29446 5500 29452
rect 5460 29170 5488 29446
rect 5448 29164 5500 29170
rect 5448 29106 5500 29112
rect 5540 29164 5592 29170
rect 5540 29106 5592 29112
rect 5356 29028 5408 29034
rect 5356 28970 5408 28976
rect 5264 28960 5316 28966
rect 5264 28902 5316 28908
rect 5368 28234 5396 28970
rect 5552 28626 5580 29106
rect 5540 28620 5592 28626
rect 5540 28562 5592 28568
rect 5736 28422 5764 29990
rect 6012 29306 6040 30126
rect 6092 29572 6144 29578
rect 6092 29514 6144 29520
rect 6000 29300 6052 29306
rect 6000 29242 6052 29248
rect 6104 29102 6132 29514
rect 6380 29306 6408 30194
rect 6472 29850 6500 30194
rect 6644 30184 6696 30190
rect 6644 30126 6696 30132
rect 6656 29850 6684 30126
rect 6840 29850 6868 30194
rect 6920 30048 6972 30054
rect 6920 29990 6972 29996
rect 6460 29844 6512 29850
rect 6460 29786 6512 29792
rect 6644 29844 6696 29850
rect 6644 29786 6696 29792
rect 6736 29844 6788 29850
rect 6736 29786 6788 29792
rect 6828 29844 6880 29850
rect 6828 29786 6880 29792
rect 6748 29730 6776 29786
rect 6748 29702 6868 29730
rect 6368 29300 6420 29306
rect 6368 29242 6420 29248
rect 6092 29096 6144 29102
rect 6092 29038 6144 29044
rect 6104 28626 6132 29038
rect 6092 28620 6144 28626
rect 6092 28562 6144 28568
rect 6840 28490 6868 29702
rect 6932 29170 6960 29990
rect 7116 29782 7144 30262
rect 8392 30252 8444 30258
rect 8392 30194 8444 30200
rect 7104 29776 7156 29782
rect 7104 29718 7156 29724
rect 8024 29776 8076 29782
rect 8024 29718 8076 29724
rect 8300 29776 8352 29782
rect 8300 29718 8352 29724
rect 6920 29164 6972 29170
rect 6920 29106 6972 29112
rect 6932 28558 6960 29106
rect 6920 28552 6972 28558
rect 6920 28494 6972 28500
rect 6828 28484 6880 28490
rect 6828 28426 6880 28432
rect 5724 28416 5776 28422
rect 5724 28358 5776 28364
rect 5276 28218 5396 28234
rect 5264 28212 5396 28218
rect 5316 28206 5396 28212
rect 5264 28154 5316 28160
rect 5632 28076 5684 28082
rect 5632 28018 5684 28024
rect 5172 27872 5224 27878
rect 5172 27814 5224 27820
rect 5448 27872 5500 27878
rect 5448 27814 5500 27820
rect 5080 27056 5132 27062
rect 5080 26998 5132 27004
rect 4252 26376 4304 26382
rect 4252 26318 4304 26324
rect 4712 26376 4764 26382
rect 4712 26318 4764 26324
rect 4988 26376 5040 26382
rect 4988 26318 5040 26324
rect 3148 26308 3200 26314
rect 3148 26250 3200 26256
rect 3160 25974 3188 26250
rect 3976 26240 4028 26246
rect 3976 26182 4028 26188
rect 3148 25968 3200 25974
rect 3148 25910 3200 25916
rect 3988 25906 4016 26182
rect 4264 26042 4292 26318
rect 4620 26308 4672 26314
rect 4620 26250 4672 26256
rect 4252 26036 4304 26042
rect 4252 25978 4304 25984
rect 3976 25900 4028 25906
rect 3976 25842 4028 25848
rect 3056 25832 3108 25838
rect 3056 25774 3108 25780
rect 3068 24886 3096 25774
rect 4068 25696 4120 25702
rect 4068 25638 4120 25644
rect 3516 25424 3568 25430
rect 3516 25366 3568 25372
rect 3056 24880 3108 24886
rect 3056 24822 3108 24828
rect 3240 23112 3292 23118
rect 3240 23054 3292 23060
rect 2964 22772 3016 22778
rect 2964 22714 3016 22720
rect 2976 21962 3004 22714
rect 3252 22234 3280 23054
rect 3528 22710 3556 25366
rect 4080 25294 4108 25638
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4632 25498 4660 26250
rect 4620 25492 4672 25498
rect 4620 25434 4672 25440
rect 4160 25424 4212 25430
rect 4160 25366 4212 25372
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 4172 25158 4200 25366
rect 4724 25294 4752 26318
rect 5000 26246 5028 26318
rect 5092 26314 5120 26998
rect 5080 26308 5132 26314
rect 5080 26250 5132 26256
rect 4988 26240 5040 26246
rect 4988 26182 5040 26188
rect 5000 25430 5028 26182
rect 5092 25838 5120 26250
rect 5080 25832 5132 25838
rect 5080 25774 5132 25780
rect 5092 25498 5120 25774
rect 5080 25492 5132 25498
rect 5080 25434 5132 25440
rect 4988 25424 5040 25430
rect 4988 25366 5040 25372
rect 5184 25294 5212 27814
rect 5460 27402 5488 27814
rect 5448 27396 5500 27402
rect 5448 27338 5500 27344
rect 5644 26994 5672 28018
rect 5736 27606 5764 28358
rect 6840 28082 6868 28426
rect 6920 28144 6972 28150
rect 6920 28086 6972 28092
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6932 27606 6960 28086
rect 5724 27600 5776 27606
rect 5724 27542 5776 27548
rect 6920 27600 6972 27606
rect 6920 27542 6972 27548
rect 5632 26988 5684 26994
rect 5632 26930 5684 26936
rect 5644 26738 5672 26930
rect 5736 26858 5764 27542
rect 5724 26852 5776 26858
rect 5724 26794 5776 26800
rect 5644 26710 5764 26738
rect 5356 26376 5408 26382
rect 5356 26318 5408 26324
rect 5264 25968 5316 25974
rect 5264 25910 5316 25916
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 5172 25288 5224 25294
rect 5172 25230 5224 25236
rect 4620 25220 4672 25226
rect 4620 25162 4672 25168
rect 4160 25152 4212 25158
rect 4160 25094 4212 25100
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23322 4660 25162
rect 4712 24812 4764 24818
rect 4712 24754 4764 24760
rect 4160 23316 4212 23322
rect 4160 23258 4212 23264
rect 4620 23316 4672 23322
rect 4620 23258 4672 23264
rect 3608 23180 3660 23186
rect 3608 23122 3660 23128
rect 3516 22704 3568 22710
rect 3516 22646 3568 22652
rect 3620 22574 3648 23122
rect 4172 23050 4200 23258
rect 4724 23254 4752 24754
rect 5184 24614 5212 25230
rect 5276 25226 5304 25910
rect 5368 25906 5396 26318
rect 5736 25906 5764 26710
rect 5816 26512 5868 26518
rect 5816 26454 5868 26460
rect 5828 25906 5856 26454
rect 6932 26314 6960 27542
rect 7116 27470 7144 29718
rect 8036 29578 8064 29718
rect 8024 29572 8076 29578
rect 8024 29514 8076 29520
rect 8116 29232 8168 29238
rect 8312 29186 8340 29718
rect 8404 29306 8432 30194
rect 8496 29646 8524 30670
rect 9772 30660 9824 30666
rect 9772 30602 9824 30608
rect 9404 30592 9456 30598
rect 9404 30534 9456 30540
rect 8852 30184 8904 30190
rect 8852 30126 8904 30132
rect 8484 29640 8536 29646
rect 8484 29582 8536 29588
rect 8392 29300 8444 29306
rect 8392 29242 8444 29248
rect 8168 29180 8340 29186
rect 8116 29174 8340 29180
rect 8128 29158 8340 29174
rect 7748 29096 7800 29102
rect 7748 29038 7800 29044
rect 7760 27878 7788 29038
rect 7932 29028 7984 29034
rect 7932 28970 7984 28976
rect 7748 27872 7800 27878
rect 7748 27814 7800 27820
rect 7104 27464 7156 27470
rect 7104 27406 7156 27412
rect 6920 26308 6972 26314
rect 6920 26250 6972 26256
rect 5356 25900 5408 25906
rect 5356 25842 5408 25848
rect 5724 25900 5776 25906
rect 5724 25842 5776 25848
rect 5816 25900 5868 25906
rect 5816 25842 5868 25848
rect 5368 25362 5396 25842
rect 5356 25356 5408 25362
rect 5356 25298 5408 25304
rect 5264 25220 5316 25226
rect 5264 25162 5316 25168
rect 5172 24608 5224 24614
rect 5172 24550 5224 24556
rect 4712 23248 4764 23254
rect 4712 23190 4764 23196
rect 4804 23248 4856 23254
rect 4804 23190 4856 23196
rect 4160 23044 4212 23050
rect 4160 22986 4212 22992
rect 4344 22976 4396 22982
rect 4344 22918 4396 22924
rect 4356 22778 4384 22918
rect 4344 22772 4396 22778
rect 4344 22714 4396 22720
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 3608 22568 3660 22574
rect 3608 22510 3660 22516
rect 3620 22234 3648 22510
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 3608 22228 3660 22234
rect 3608 22170 3660 22176
rect 3252 22094 3280 22170
rect 4632 22098 4660 22578
rect 3160 22066 3280 22094
rect 4620 22092 4672 22098
rect 2964 21956 3016 21962
rect 2964 21898 3016 21904
rect 1860 21888 1912 21894
rect 1860 21830 1912 21836
rect 1872 21554 1900 21830
rect 1860 21548 1912 21554
rect 1860 21490 1912 21496
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 2792 20942 2820 21422
rect 2872 21344 2924 21350
rect 2872 21286 2924 21292
rect 2780 20936 2832 20942
rect 2780 20878 2832 20884
rect 2792 20602 2820 20878
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2884 20466 2912 21286
rect 2976 20874 3004 21898
rect 3160 21350 3188 22066
rect 4620 22034 4672 22040
rect 4816 22030 4844 23190
rect 4436 22024 4488 22030
rect 4436 21966 4488 21972
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 4252 21956 4304 21962
rect 4252 21898 4304 21904
rect 4264 21554 4292 21898
rect 4448 21554 4476 21966
rect 4252 21548 4304 21554
rect 4252 21490 4304 21496
rect 4436 21548 4488 21554
rect 4436 21490 4488 21496
rect 5080 21548 5132 21554
rect 5080 21490 5132 21496
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 3148 21344 3200 21350
rect 3148 21286 3200 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4620 21072 4672 21078
rect 4620 21014 4672 21020
rect 2964 20868 3016 20874
rect 2964 20810 3016 20816
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 2884 18766 2912 20402
rect 2976 18766 3004 20810
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4632 18834 4660 21014
rect 4712 20460 4764 20466
rect 4712 20402 4764 20408
rect 4724 18970 4752 20402
rect 4816 19378 4844 21422
rect 5092 19378 5120 21490
rect 5276 20806 5304 25162
rect 5368 23118 5396 25298
rect 5356 23112 5408 23118
rect 5356 23054 5408 23060
rect 5264 20800 5316 20806
rect 5264 20742 5316 20748
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2964 18760 3016 18766
rect 2964 18702 3016 18708
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 2136 18624 2188 18630
rect 2136 18566 2188 18572
rect 2148 18358 2176 18566
rect 2136 18352 2188 18358
rect 2136 18294 2188 18300
rect 2780 18352 2832 18358
rect 2780 18294 2832 18300
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 2700 17762 2728 18158
rect 2792 17882 2820 18294
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 1400 17740 1452 17746
rect 2700 17734 2820 17762
rect 1400 17682 1452 17688
rect 2792 17678 2820 17734
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2884 16794 2912 18702
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2976 16522 3004 18702
rect 3988 18426 4016 18702
rect 4436 18624 4488 18630
rect 4436 18566 4488 18572
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 4448 18154 4476 18566
rect 4724 18222 4752 18906
rect 4816 18290 4844 19314
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4908 18698 4936 19110
rect 4896 18692 4948 18698
rect 4896 18634 4948 18640
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4436 18148 4488 18154
rect 4436 18090 4488 18096
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4620 16720 4672 16726
rect 4620 16662 4672 16668
rect 2964 16516 3016 16522
rect 2964 16458 3016 16464
rect 2136 15156 2188 15162
rect 2136 15098 2188 15104
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1688 14074 1716 14554
rect 2148 14414 2176 15098
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2700 14278 2728 14894
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1872 13938 1900 14214
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 2792 13870 2820 14350
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2792 13530 2820 13806
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1872 9042 1900 9318
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1596 8634 1624 8910
rect 2792 8838 2820 13262
rect 2884 13258 2912 14010
rect 2872 13252 2924 13258
rect 2872 13194 2924 13200
rect 2976 9586 3004 16458
rect 3240 16176 3292 16182
rect 3240 16118 3292 16124
rect 3148 14952 3200 14958
rect 3148 14894 3200 14900
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 3068 14482 3096 14554
rect 3160 14482 3188 14894
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 3068 13394 3096 14214
rect 3160 13954 3188 14418
rect 3252 14414 3280 16118
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3252 14278 3280 14350
rect 3804 14346 3832 14758
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 3792 14340 3844 14346
rect 3792 14282 3844 14288
rect 3240 14272 3292 14278
rect 3240 14214 3292 14220
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3160 13926 3280 13954
rect 3148 13864 3200 13870
rect 3148 13806 3200 13812
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 3160 13326 3188 13806
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3160 12850 3188 13262
rect 3252 13258 3280 13926
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 3252 12918 3280 13194
rect 3240 12912 3292 12918
rect 3240 12854 3292 12860
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3436 12646 3464 14010
rect 3804 13870 3832 14282
rect 3988 13938 4016 14554
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 3804 13734 3832 13806
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3988 13530 4016 13874
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 4632 13258 4660 16662
rect 4724 16522 4752 18158
rect 5092 17678 5120 19314
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 5092 16794 5120 17614
rect 5276 17134 5304 20742
rect 5368 17202 5396 23054
rect 5736 22642 5764 25842
rect 5724 22636 5776 22642
rect 5724 22578 5776 22584
rect 6932 21894 6960 26250
rect 7116 25906 7144 27406
rect 7104 25900 7156 25906
rect 7104 25842 7156 25848
rect 7564 25900 7616 25906
rect 7564 25842 7616 25848
rect 7576 22982 7604 25842
rect 7760 25158 7788 27814
rect 7840 25492 7892 25498
rect 7840 25434 7892 25440
rect 7852 25294 7880 25434
rect 7840 25288 7892 25294
rect 7840 25230 7892 25236
rect 7748 25152 7800 25158
rect 7748 25094 7800 25100
rect 7852 23322 7880 25230
rect 7944 24818 7972 28970
rect 8312 28626 8340 29158
rect 8300 28620 8352 28626
rect 8300 28562 8352 28568
rect 8404 28082 8432 29242
rect 8392 28076 8444 28082
rect 8392 28018 8444 28024
rect 8496 26586 8524 29582
rect 8484 26580 8536 26586
rect 8484 26522 8536 26528
rect 8576 25832 8628 25838
rect 8576 25774 8628 25780
rect 8300 25696 8352 25702
rect 8300 25638 8352 25644
rect 8312 25294 8340 25638
rect 8588 25362 8616 25774
rect 8576 25356 8628 25362
rect 8576 25298 8628 25304
rect 8300 25288 8352 25294
rect 8300 25230 8352 25236
rect 7932 24812 7984 24818
rect 7932 24754 7984 24760
rect 8864 24698 8892 30126
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 9324 29306 9352 29582
rect 9312 29300 9364 29306
rect 9312 29242 9364 29248
rect 9220 29096 9272 29102
rect 9220 29038 9272 29044
rect 9232 28762 9260 29038
rect 9220 28756 9272 28762
rect 9220 28698 9272 28704
rect 9416 28558 9444 30534
rect 9784 30326 9812 30602
rect 9772 30320 9824 30326
rect 9772 30262 9824 30268
rect 9680 29776 9732 29782
rect 9680 29718 9732 29724
rect 9692 28558 9720 29718
rect 9784 29714 9812 30262
rect 9772 29708 9824 29714
rect 9772 29650 9824 29656
rect 10336 29646 10364 30738
rect 12084 30734 12112 31078
rect 12072 30728 12124 30734
rect 12072 30670 12124 30676
rect 10968 30252 11020 30258
rect 10968 30194 11020 30200
rect 10784 30184 10836 30190
rect 10784 30126 10836 30132
rect 10796 29850 10824 30126
rect 10784 29844 10836 29850
rect 10784 29786 10836 29792
rect 10324 29640 10376 29646
rect 10324 29582 10376 29588
rect 10232 29572 10284 29578
rect 10232 29514 10284 29520
rect 10244 28762 10272 29514
rect 10336 29306 10364 29582
rect 10324 29300 10376 29306
rect 10324 29242 10376 29248
rect 10600 28960 10652 28966
rect 10600 28902 10652 28908
rect 10232 28756 10284 28762
rect 10232 28698 10284 28704
rect 10612 28558 10640 28902
rect 10796 28694 10824 29786
rect 10980 29782 11008 30194
rect 11152 30116 11204 30122
rect 11152 30058 11204 30064
rect 11060 30048 11112 30054
rect 11060 29990 11112 29996
rect 10968 29776 11020 29782
rect 10968 29718 11020 29724
rect 10980 29646 11008 29718
rect 10968 29640 11020 29646
rect 10968 29582 11020 29588
rect 11072 28762 11100 29990
rect 11164 29782 11192 30058
rect 11152 29776 11204 29782
rect 11152 29718 11204 29724
rect 11060 28756 11112 28762
rect 11060 28698 11112 28704
rect 10784 28688 10836 28694
rect 10784 28630 10836 28636
rect 9404 28552 9456 28558
rect 9404 28494 9456 28500
rect 9680 28552 9732 28558
rect 9680 28494 9732 28500
rect 9864 28552 9916 28558
rect 9864 28494 9916 28500
rect 10324 28552 10376 28558
rect 10324 28494 10376 28500
rect 10600 28552 10652 28558
rect 10600 28494 10652 28500
rect 9876 28218 9904 28494
rect 9864 28212 9916 28218
rect 9864 28154 9916 28160
rect 10336 28082 10364 28494
rect 10324 28076 10376 28082
rect 10324 28018 10376 28024
rect 8944 26376 8996 26382
rect 8944 26318 8996 26324
rect 9588 26376 9640 26382
rect 9588 26318 9640 26324
rect 10140 26376 10192 26382
rect 10140 26318 10192 26324
rect 8956 25974 8984 26318
rect 9496 26240 9548 26246
rect 9496 26182 9548 26188
rect 8944 25968 8996 25974
rect 8944 25910 8996 25916
rect 9508 25770 9536 26182
rect 9496 25764 9548 25770
rect 9496 25706 9548 25712
rect 9600 25498 9628 26318
rect 9864 26308 9916 26314
rect 9864 26250 9916 26256
rect 9876 25906 9904 26250
rect 10152 25922 10180 26318
rect 10232 26240 10284 26246
rect 10232 26182 10284 26188
rect 10060 25906 10180 25922
rect 9864 25900 9916 25906
rect 9864 25842 9916 25848
rect 10048 25900 10180 25906
rect 10100 25894 10180 25900
rect 10048 25842 10100 25848
rect 9680 25696 9732 25702
rect 9680 25638 9732 25644
rect 9588 25492 9640 25498
rect 9588 25434 9640 25440
rect 9692 25362 9720 25638
rect 9680 25356 9732 25362
rect 9680 25298 9732 25304
rect 9680 25220 9732 25226
rect 9680 25162 9732 25168
rect 9128 25152 9180 25158
rect 9128 25094 9180 25100
rect 9140 24818 9168 25094
rect 9128 24812 9180 24818
rect 9128 24754 9180 24760
rect 9588 24744 9640 24750
rect 8864 24682 9168 24698
rect 9588 24686 9640 24692
rect 8864 24676 9180 24682
rect 8864 24670 9128 24676
rect 9128 24618 9180 24624
rect 8208 24608 8260 24614
rect 8208 24550 8260 24556
rect 8024 23520 8076 23526
rect 8024 23462 8076 23468
rect 7840 23316 7892 23322
rect 7840 23258 7892 23264
rect 7656 23044 7708 23050
rect 7656 22986 7708 22992
rect 7932 23044 7984 23050
rect 7932 22986 7984 22992
rect 7564 22976 7616 22982
rect 7564 22918 7616 22924
rect 7668 22778 7696 22986
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 7656 22772 7708 22778
rect 7656 22714 7708 22720
rect 7012 22636 7064 22642
rect 7012 22578 7064 22584
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 6920 21888 6972 21894
rect 6920 21830 6972 21836
rect 5448 21480 5500 21486
rect 5448 21422 5500 21428
rect 5460 20874 5488 21422
rect 6932 21146 6960 21830
rect 7024 21690 7052 22578
rect 7104 22500 7156 22506
rect 7104 22442 7156 22448
rect 7012 21684 7064 21690
rect 7012 21626 7064 21632
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 7024 20992 7052 21626
rect 7116 21010 7144 22442
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7300 21486 7328 21966
rect 7392 21690 7420 22578
rect 7760 22438 7788 22918
rect 7748 22432 7800 22438
rect 7748 22374 7800 22380
rect 7564 22160 7616 22166
rect 7564 22102 7616 22108
rect 7472 21956 7524 21962
rect 7472 21898 7524 21904
rect 7380 21684 7432 21690
rect 7380 21626 7432 21632
rect 7288 21480 7340 21486
rect 7288 21422 7340 21428
rect 6932 20964 7052 20992
rect 7104 21004 7156 21010
rect 5448 20868 5500 20874
rect 5448 20810 5500 20816
rect 6932 20602 6960 20964
rect 7104 20946 7156 20952
rect 7012 20868 7064 20874
rect 7012 20810 7064 20816
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6932 19378 6960 20538
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6092 19168 6144 19174
rect 6092 19110 6144 19116
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5460 18086 5488 18226
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5368 16658 5396 17002
rect 5460 16674 5488 18022
rect 5736 17338 5764 18566
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5908 17264 5960 17270
rect 5908 17206 5960 17212
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 5356 16652 5408 16658
rect 5460 16646 5580 16674
rect 5356 16594 5408 16600
rect 4712 16516 4764 16522
rect 4712 16458 4764 16464
rect 4724 14958 4752 16458
rect 5092 16250 5120 16594
rect 5368 16538 5396 16594
rect 5184 16510 5396 16538
rect 5080 16244 5132 16250
rect 5080 16186 5132 16192
rect 4712 14952 4764 14958
rect 4712 14894 4764 14900
rect 4160 13252 4212 13258
rect 4160 13194 4212 13200
rect 4620 13252 4672 13258
rect 4672 13212 4752 13240
rect 4620 13194 4672 13200
rect 4172 12986 4200 13194
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4356 12918 4384 13126
rect 3976 12912 4028 12918
rect 3976 12854 4028 12860
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3988 10130 4016 12854
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4080 12238 4108 12786
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12306 4660 12582
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4724 12238 4752 13212
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2976 9178 3004 9522
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 2792 8498 2820 8774
rect 2976 8566 3004 8910
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 4080 7886 4108 9114
rect 4632 8498 4660 12038
rect 5184 10674 5212 16510
rect 5552 16114 5580 16646
rect 5920 16114 5948 17206
rect 6000 16516 6052 16522
rect 6000 16458 6052 16464
rect 6012 16182 6040 16458
rect 6000 16176 6052 16182
rect 6000 16118 6052 16124
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 5460 12850 5488 15982
rect 5552 15502 5580 16050
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 6012 12986 6040 13126
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5460 12374 5488 12786
rect 5448 12368 5500 12374
rect 5448 12310 5500 12316
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 5276 10674 5304 12174
rect 5460 11098 5488 12310
rect 5368 11070 5488 11098
rect 5724 11076 5776 11082
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 4724 9994 4752 10610
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5778 4660 7754
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4724 4146 4752 9930
rect 5368 8566 5396 11070
rect 5724 11018 5776 11024
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5460 10266 5488 10950
rect 5736 10810 5764 11018
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5368 7818 5396 8502
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5460 7274 5488 8434
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5552 5302 5580 8570
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5552 4622 5580 5238
rect 5644 5234 5672 8774
rect 6104 6866 6132 19110
rect 6748 18698 6776 19314
rect 7024 19310 7052 20810
rect 7116 19514 7144 20946
rect 7392 20466 7420 21626
rect 7484 21554 7512 21898
rect 7576 21554 7604 22102
rect 7760 21622 7788 22374
rect 7944 22234 7972 22986
rect 8036 22710 8064 23462
rect 8220 22930 8248 24550
rect 8220 22902 8432 22930
rect 8404 22778 8432 22902
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8392 22772 8444 22778
rect 8392 22714 8444 22720
rect 8024 22704 8076 22710
rect 8024 22646 8076 22652
rect 7932 22228 7984 22234
rect 7932 22170 7984 22176
rect 8036 21962 8064 22646
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 8220 22094 8248 22578
rect 8128 22066 8248 22094
rect 8024 21956 8076 21962
rect 8024 21898 8076 21904
rect 8128 21622 8156 22066
rect 8312 22030 8340 22714
rect 8392 22568 8444 22574
rect 8392 22510 8444 22516
rect 8404 22166 8432 22510
rect 8576 22432 8628 22438
rect 8576 22374 8628 22380
rect 8392 22160 8444 22166
rect 8392 22102 8444 22108
rect 8588 22098 8616 22374
rect 8576 22092 8628 22098
rect 8576 22034 8628 22040
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 8220 21894 8248 21925
rect 8208 21888 8260 21894
rect 8496 21842 8524 21966
rect 8260 21836 8524 21842
rect 8208 21830 8524 21836
rect 8220 21814 8524 21830
rect 7748 21616 7800 21622
rect 7748 21558 7800 21564
rect 8116 21616 8168 21622
rect 8116 21558 8168 21564
rect 7472 21548 7524 21554
rect 7472 21490 7524 21496
rect 7564 21548 7616 21554
rect 7564 21490 7616 21496
rect 7484 21010 7512 21490
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7380 20460 7432 20466
rect 7380 20402 7432 20408
rect 7484 20262 7512 20946
rect 7576 20942 7604 21490
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7576 20534 7604 20878
rect 7564 20528 7616 20534
rect 7564 20470 7616 20476
rect 8220 20330 8248 21814
rect 9140 21554 9168 24618
rect 9600 24614 9628 24686
rect 9220 24608 9272 24614
rect 9220 24550 9272 24556
rect 9588 24608 9640 24614
rect 9588 24550 9640 24556
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 8300 21344 8352 21350
rect 8300 21286 8352 21292
rect 8208 20324 8260 20330
rect 8208 20266 8260 20272
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7748 20256 7800 20262
rect 7748 20198 7800 20204
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 7024 18970 7052 19246
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 7116 18766 7144 19450
rect 7760 19174 7788 20198
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 6736 18692 6788 18698
rect 6736 18634 6788 18640
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6184 16448 6236 16454
rect 6184 16390 6236 16396
rect 6196 11150 6224 16390
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6564 11082 6592 16934
rect 6840 16182 6868 17478
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 6840 16046 6868 16118
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 7116 15162 7144 18702
rect 8312 17610 8340 21286
rect 9140 21162 9168 21490
rect 9232 21350 9260 24550
rect 9588 22568 9640 22574
rect 9692 22522 9720 25162
rect 9876 24954 9904 25842
rect 10060 25294 10088 25842
rect 10244 25838 10272 26182
rect 10232 25832 10284 25838
rect 10232 25774 10284 25780
rect 10048 25288 10100 25294
rect 10048 25230 10100 25236
rect 9864 24948 9916 24954
rect 9864 24890 9916 24896
rect 9640 22516 9720 22522
rect 9588 22510 9720 22516
rect 9600 22494 9720 22510
rect 9692 22030 9720 22494
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9784 22166 9812 22374
rect 9772 22160 9824 22166
rect 9772 22102 9824 22108
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 9680 22024 9732 22030
rect 9680 21966 9732 21972
rect 9324 21690 9352 21966
rect 9312 21684 9364 21690
rect 9312 21626 9364 21632
rect 9404 21480 9456 21486
rect 9404 21422 9456 21428
rect 9220 21344 9272 21350
rect 9220 21286 9272 21292
rect 9140 21134 9260 21162
rect 9036 20868 9088 20874
rect 9036 20810 9088 20816
rect 9048 20466 9076 20810
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8300 17604 8352 17610
rect 8300 17546 8352 17552
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7668 16522 7696 17138
rect 7656 16516 7708 16522
rect 7656 16458 7708 16464
rect 7288 16176 7340 16182
rect 7288 16118 7340 16124
rect 7300 15570 7328 16118
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7668 15502 7696 16458
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8220 15638 8248 15846
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6656 11218 6684 13262
rect 8220 13258 8248 15574
rect 8312 13258 8340 17546
rect 8496 17338 8524 17614
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 7564 13252 7616 13258
rect 7564 13194 7616 13200
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 8300 13252 8352 13258
rect 8300 13194 8352 13200
rect 7484 12442 7512 13194
rect 7576 12850 7604 13194
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 7576 11150 7604 12786
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 5724 5636 5776 5642
rect 5724 5578 5776 5584
rect 5736 5302 5764 5578
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5644 4690 5672 5170
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 5920 3602 5948 4082
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 6380 3058 6408 4558
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 848 2984 900 2990
rect 848 2926 900 2932
rect 860 800 888 2926
rect 6472 2774 6500 10950
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6748 8498 6776 8774
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6564 7886 6592 8230
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6748 7750 6776 8434
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6932 7478 6960 8026
rect 7024 7546 7052 8298
rect 8312 8090 8340 8366
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6564 6798 6592 7142
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6564 2990 6592 4558
rect 6656 3738 6684 6598
rect 7024 5914 7052 6802
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8220 4622 8248 5102
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6932 3466 6960 4490
rect 7944 4282 7972 4490
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 8220 3738 8248 4558
rect 8312 3942 8340 7210
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8312 3534 8340 3878
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 8496 3126 8524 13126
rect 8772 12918 8800 13806
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8772 11218 8800 12854
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8956 7954 8984 19314
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9140 17678 9168 18566
rect 9232 18290 9260 21134
rect 9416 20806 9444 21422
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 9692 20466 9720 21966
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9784 20942 9812 21830
rect 9876 21622 9904 21830
rect 9864 21616 9916 21622
rect 9864 21558 9916 21564
rect 9876 21010 9904 21558
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 9864 21004 9916 21010
rect 9864 20946 9916 20952
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9140 16250 9168 17614
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9140 16114 9168 16186
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9140 10674 9168 12174
rect 9232 10742 9260 18226
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9416 17610 9444 18158
rect 9404 17604 9456 17610
rect 9404 17546 9456 17552
rect 9416 11150 9444 17546
rect 10152 17542 10180 18566
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10244 17066 10272 21490
rect 10336 17338 10364 28018
rect 10612 26874 10640 28494
rect 10612 26846 10732 26874
rect 10600 26784 10652 26790
rect 10600 26726 10652 26732
rect 10508 25492 10560 25498
rect 10508 25434 10560 25440
rect 10520 24954 10548 25434
rect 10612 25294 10640 26726
rect 10704 25294 10732 26846
rect 10796 26042 10824 28630
rect 12084 26382 12112 30670
rect 12728 30190 12756 31300
rect 12716 30184 12768 30190
rect 12716 30126 12768 30132
rect 12532 26920 12584 26926
rect 12532 26862 12584 26868
rect 12544 26586 12572 26862
rect 12532 26580 12584 26586
rect 12532 26522 12584 26528
rect 12072 26376 12124 26382
rect 12072 26318 12124 26324
rect 12440 26376 12492 26382
rect 12440 26318 12492 26324
rect 12452 26042 12480 26318
rect 10784 26036 10836 26042
rect 10784 25978 10836 25984
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 10600 25288 10652 25294
rect 10600 25230 10652 25236
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 10508 24948 10560 24954
rect 10508 24890 10560 24896
rect 10416 20800 10468 20806
rect 10416 20742 10468 20748
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9508 16046 9536 16934
rect 9956 16176 10008 16182
rect 9956 16118 10008 16124
rect 9496 16040 9548 16046
rect 9496 15982 9548 15988
rect 9508 13938 9536 15982
rect 9968 15570 9996 16118
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9772 15496 9824 15502
rect 9692 15444 9772 15450
rect 9692 15438 9824 15444
rect 9692 15422 9812 15438
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9508 12170 9536 13874
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9220 10736 9272 10742
rect 9220 10678 9272 10684
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9140 10130 9168 10610
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9416 9994 9444 11086
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9404 9988 9456 9994
rect 9404 9930 9456 9936
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8956 4146 8984 7890
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8956 3398 8984 4082
rect 9140 3602 9168 4422
rect 9232 4078 9260 9930
rect 9508 7954 9536 12106
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9508 7392 9536 7890
rect 9588 7404 9640 7410
rect 9508 7364 9588 7392
rect 9588 7346 9640 7352
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9232 3466 9260 4014
rect 9220 3460 9272 3466
rect 9220 3402 9272 3408
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8484 3120 8536 3126
rect 8484 3062 8536 3068
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 9692 2922 9720 15422
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9784 12322 9812 13330
rect 10152 12986 10180 13670
rect 10244 12986 10272 17002
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 10428 12850 10456 20742
rect 10612 18766 10640 25230
rect 10704 21554 10732 25230
rect 10796 25226 10824 25978
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 10784 25220 10836 25226
rect 10784 25162 10836 25168
rect 12636 24818 12664 25230
rect 12624 24812 12676 24818
rect 12624 24754 12676 24760
rect 12728 23730 12756 30126
rect 13832 29714 13860 31418
rect 14108 30190 14136 35430
rect 14096 30184 14148 30190
rect 14096 30126 14148 30132
rect 13820 29708 13872 29714
rect 13820 29650 13872 29656
rect 13360 29504 13412 29510
rect 13360 29446 13412 29452
rect 13372 26926 13400 29446
rect 13820 29028 13872 29034
rect 13820 28970 13872 28976
rect 13832 26994 13860 28970
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 13360 26920 13412 26926
rect 13360 26862 13412 26868
rect 12900 25220 12952 25226
rect 12900 25162 12952 25168
rect 12912 24818 12940 25162
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 12716 23724 12768 23730
rect 12716 23666 12768 23672
rect 11888 23248 11940 23254
rect 11888 23190 11940 23196
rect 10968 23180 11020 23186
rect 10968 23122 11020 23128
rect 10980 22098 11008 23122
rect 11900 22778 11928 23190
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 11900 22642 11928 22714
rect 11888 22636 11940 22642
rect 11888 22578 11940 22584
rect 12072 22568 12124 22574
rect 12072 22510 12124 22516
rect 10968 22092 11020 22098
rect 10968 22034 11020 22040
rect 12084 22030 12112 22510
rect 12728 22234 12756 23666
rect 12992 23112 13044 23118
rect 12992 23054 13044 23060
rect 13176 23112 13228 23118
rect 13176 23054 13228 23060
rect 12808 23044 12860 23050
rect 12808 22986 12860 22992
rect 12716 22228 12768 22234
rect 12716 22170 12768 22176
rect 12820 22094 12848 22986
rect 13004 22438 13032 23054
rect 12992 22432 13044 22438
rect 12992 22374 13044 22380
rect 12728 22066 12848 22094
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10876 21548 10928 21554
rect 10876 21490 10928 21496
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 10888 21146 10916 21490
rect 11980 21344 12032 21350
rect 11980 21286 12032 21292
rect 10876 21140 10928 21146
rect 10876 21082 10928 21088
rect 11992 20942 12020 21286
rect 12084 21146 12112 21490
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 12072 21140 12124 21146
rect 12072 21082 12124 21088
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 12084 20602 12112 21082
rect 12440 21004 12492 21010
rect 12440 20946 12492 20952
rect 12072 20596 12124 20602
rect 12072 20538 12124 20544
rect 12452 20466 12480 20946
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 12544 20398 12572 21422
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10692 18692 10744 18698
rect 10692 18634 10744 18640
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10612 17882 10640 18226
rect 10704 18086 10732 18634
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10612 17134 10640 17818
rect 10704 17202 10732 18022
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 10784 17604 10836 17610
rect 10784 17546 10836 17552
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10520 15434 10548 15846
rect 10508 15428 10560 15434
rect 10508 15370 10560 15376
rect 10520 12918 10548 15370
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10060 12442 10088 12786
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10244 12322 10272 12718
rect 9784 12294 10272 12322
rect 9784 10606 9812 12294
rect 10428 10674 10456 12786
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10520 10810 10548 10950
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9784 5574 9812 10542
rect 10060 10266 10088 10610
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9784 4758 9812 5510
rect 10152 5370 10180 8298
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9968 4282 9996 5170
rect 10244 4554 10272 8366
rect 10428 7546 10456 10610
rect 10612 8430 10640 17070
rect 10796 17066 10824 17546
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10980 17270 11008 17478
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10980 10674 11008 17206
rect 12176 17134 12204 17614
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 12176 15570 12204 17070
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10888 8090 10916 8434
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10428 6934 10456 7482
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10416 6928 10468 6934
rect 10416 6870 10468 6876
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10336 4622 10364 5646
rect 10428 4826 10456 6870
rect 10704 6866 10732 7142
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10888 6798 10916 8026
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10520 6390 10548 6598
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10232 4548 10284 4554
rect 10232 4490 10284 4496
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10152 3074 10180 3130
rect 9968 3058 10180 3074
rect 9956 3052 10180 3058
rect 10008 3046 10180 3052
rect 9956 2994 10008 3000
rect 10244 2990 10272 4150
rect 10520 3738 10548 4558
rect 10704 4282 10732 4558
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 11072 3466 11100 12582
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11164 9722 11192 10406
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 6380 2746 6500 2774
rect 6380 2650 6408 2746
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6380 2446 6408 2586
rect 11072 2582 11100 3402
rect 11164 2582 11192 9658
rect 12636 8294 12664 12582
rect 12728 8566 12756 22066
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 12912 18290 12940 19790
rect 13004 18970 13032 22374
rect 13188 21486 13216 23054
rect 13176 21480 13228 21486
rect 13176 21422 13228 21428
rect 13176 21344 13228 21350
rect 13176 21286 13228 21292
rect 13188 19854 13216 21286
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 13372 18426 13400 26862
rect 13832 26382 13860 26930
rect 14200 26926 14228 36246
rect 14292 35834 14320 37334
rect 14464 36712 14516 36718
rect 14464 36654 14516 36660
rect 14476 36106 14504 36654
rect 14936 36242 14964 37334
rect 15028 37244 15056 39200
rect 17224 37460 17276 37466
rect 17224 37402 17276 37408
rect 15200 37256 15252 37262
rect 15028 37216 15200 37244
rect 15200 37198 15252 37204
rect 15292 37120 15344 37126
rect 15292 37062 15344 37068
rect 14924 36236 14976 36242
rect 14924 36178 14976 36184
rect 14464 36100 14516 36106
rect 14464 36042 14516 36048
rect 14280 35828 14332 35834
rect 14280 35770 14332 35776
rect 14476 35630 14504 36042
rect 15304 36038 15332 37062
rect 15752 36304 15804 36310
rect 15752 36246 15804 36252
rect 15292 36032 15344 36038
rect 15292 35974 15344 35980
rect 14464 35624 14516 35630
rect 14464 35566 14516 35572
rect 15108 31748 15160 31754
rect 15108 31690 15160 31696
rect 15120 31346 15148 31690
rect 15108 31340 15160 31346
rect 15108 31282 15160 31288
rect 14372 30864 14424 30870
rect 14372 30806 14424 30812
rect 14384 30326 14412 30806
rect 15120 30734 15148 31282
rect 14556 30728 14608 30734
rect 14556 30670 14608 30676
rect 15108 30728 15160 30734
rect 15108 30670 15160 30676
rect 14372 30320 14424 30326
rect 14372 30262 14424 30268
rect 14464 29640 14516 29646
rect 14464 29582 14516 29588
rect 14476 29510 14504 29582
rect 14280 29504 14332 29510
rect 14280 29446 14332 29452
rect 14464 29504 14516 29510
rect 14464 29446 14516 29452
rect 14292 29170 14320 29446
rect 14476 29238 14504 29446
rect 14464 29232 14516 29238
rect 14464 29174 14516 29180
rect 14280 29164 14332 29170
rect 14280 29106 14332 29112
rect 14372 27532 14424 27538
rect 14372 27474 14424 27480
rect 14280 27464 14332 27470
rect 14280 27406 14332 27412
rect 14292 26994 14320 27406
rect 14280 26988 14332 26994
rect 14280 26930 14332 26936
rect 14004 26920 14056 26926
rect 14004 26862 14056 26868
rect 14188 26920 14240 26926
rect 14188 26862 14240 26868
rect 14016 26790 14044 26862
rect 14004 26784 14056 26790
rect 14004 26726 14056 26732
rect 13820 26376 13872 26382
rect 13820 26318 13872 26324
rect 13832 25906 13860 26318
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 13452 25288 13504 25294
rect 13452 25230 13504 25236
rect 13464 24818 13492 25230
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13464 21010 13492 24754
rect 14016 22438 14044 26726
rect 14200 23662 14228 26862
rect 14188 23656 14240 23662
rect 14188 23598 14240 23604
rect 14292 23202 14320 26930
rect 14384 26382 14412 27474
rect 14476 27470 14504 29174
rect 14464 27464 14516 27470
rect 14464 27406 14516 27412
rect 14372 26376 14424 26382
rect 14372 26318 14424 26324
rect 14464 25424 14516 25430
rect 14464 25366 14516 25372
rect 14372 23792 14424 23798
rect 14372 23734 14424 23740
rect 14384 23322 14412 23734
rect 14372 23316 14424 23322
rect 14372 23258 14424 23264
rect 14200 23174 14320 23202
rect 14200 23050 14228 23174
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14188 23044 14240 23050
rect 14188 22986 14240 22992
rect 14292 22710 14320 23054
rect 14384 22778 14412 23054
rect 14372 22772 14424 22778
rect 14372 22714 14424 22720
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 14004 22432 14056 22438
rect 14004 22374 14056 22380
rect 14372 22024 14424 22030
rect 14372 21966 14424 21972
rect 14384 21690 14412 21966
rect 14372 21684 14424 21690
rect 14372 21626 14424 21632
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13452 21004 13504 21010
rect 13452 20946 13504 20952
rect 13912 20936 13964 20942
rect 13912 20878 13964 20884
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 13648 19718 13676 20334
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13464 18970 13492 19314
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 13360 17604 13412 17610
rect 13360 17546 13412 17552
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13280 16794 13308 17138
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13372 16250 13400 17546
rect 13648 16590 13676 19654
rect 13832 18358 13860 20198
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13360 16244 13412 16250
rect 13360 16186 13412 16192
rect 13464 15366 13492 16526
rect 13648 16182 13676 16526
rect 13636 16176 13688 16182
rect 13636 16118 13688 16124
rect 13740 16114 13768 17478
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13464 14414 13492 15302
rect 13740 15094 13768 16050
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 13924 15026 13952 20878
rect 14016 19514 14044 21490
rect 14476 20942 14504 25366
rect 14568 23118 14596 30670
rect 15200 30252 15252 30258
rect 15120 30212 15200 30240
rect 14832 30048 14884 30054
rect 14832 29990 14884 29996
rect 14844 29646 14872 29990
rect 14832 29640 14884 29646
rect 14832 29582 14884 29588
rect 14924 29572 14976 29578
rect 14924 29514 14976 29520
rect 14936 29034 14964 29514
rect 15120 29510 15148 30212
rect 15200 30194 15252 30200
rect 15764 29646 15792 36246
rect 17236 36242 17264 37402
rect 18340 37262 18368 39200
rect 21652 39114 21680 39200
rect 21744 39114 21772 39222
rect 21652 39086 21772 39114
rect 18328 37256 18380 37262
rect 18328 37198 18380 37204
rect 22020 37210 22048 39222
rect 24950 39200 25006 40000
rect 28262 39200 28318 40000
rect 31574 39200 31630 40000
rect 34886 39200 34942 40000
rect 38198 39200 38254 40000
rect 24964 37262 24992 39200
rect 28276 37262 28304 39200
rect 24952 37256 25004 37262
rect 22020 37194 22140 37210
rect 24952 37198 25004 37204
rect 28264 37256 28316 37262
rect 28264 37198 28316 37204
rect 31588 37210 31616 39200
rect 34900 37754 34928 39200
rect 34808 37726 34928 37754
rect 34808 37262 34836 37726
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 37188 37324 37240 37330
rect 37188 37266 37240 37272
rect 31760 37256 31812 37262
rect 31588 37204 31760 37210
rect 31588 37198 31812 37204
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 22020 37188 22152 37194
rect 22020 37182 22100 37188
rect 31588 37182 31800 37198
rect 22100 37130 22152 37136
rect 18604 37120 18656 37126
rect 18604 37062 18656 37068
rect 22192 37120 22244 37126
rect 22192 37062 22244 37068
rect 25228 37120 25280 37126
rect 25228 37062 25280 37068
rect 34520 37120 34572 37126
rect 34520 37062 34572 37068
rect 18616 36242 18644 37062
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 22204 36922 22232 37062
rect 22192 36916 22244 36922
rect 22192 36858 22244 36864
rect 19432 36848 19484 36854
rect 19432 36790 19484 36796
rect 18696 36780 18748 36786
rect 18696 36722 18748 36728
rect 17224 36236 17276 36242
rect 17224 36178 17276 36184
rect 18604 36236 18656 36242
rect 18604 36178 18656 36184
rect 17408 36168 17460 36174
rect 17328 36116 17408 36122
rect 17328 36110 17460 36116
rect 17328 36094 17448 36110
rect 17776 36100 17828 36106
rect 17224 34536 17276 34542
rect 17224 34478 17276 34484
rect 17236 33998 17264 34478
rect 17224 33992 17276 33998
rect 17224 33934 17276 33940
rect 17236 33522 17264 33934
rect 17224 33516 17276 33522
rect 17224 33458 17276 33464
rect 17236 33114 17264 33458
rect 17224 33108 17276 33114
rect 17224 33050 17276 33056
rect 17328 32450 17356 36094
rect 17776 36042 17828 36048
rect 17408 34604 17460 34610
rect 17408 34546 17460 34552
rect 17420 33998 17448 34546
rect 17408 33992 17460 33998
rect 17408 33934 17460 33940
rect 17420 33590 17448 33934
rect 17408 33584 17460 33590
rect 17408 33526 17460 33532
rect 17500 33516 17552 33522
rect 17500 33458 17552 33464
rect 17592 33516 17644 33522
rect 17592 33458 17644 33464
rect 17512 33386 17540 33458
rect 17500 33380 17552 33386
rect 17500 33322 17552 33328
rect 17512 32570 17540 33322
rect 17604 32570 17632 33458
rect 17684 32836 17736 32842
rect 17684 32778 17736 32784
rect 17500 32564 17552 32570
rect 17500 32506 17552 32512
rect 17592 32564 17644 32570
rect 17592 32506 17644 32512
rect 17328 32422 17540 32450
rect 17224 31884 17276 31890
rect 17224 31826 17276 31832
rect 17132 31340 17184 31346
rect 17132 31282 17184 31288
rect 15844 31272 15896 31278
rect 15844 31214 15896 31220
rect 15856 30666 15884 31214
rect 15844 30660 15896 30666
rect 15844 30602 15896 30608
rect 15752 29640 15804 29646
rect 15752 29582 15804 29588
rect 15108 29504 15160 29510
rect 15108 29446 15160 29452
rect 14924 29028 14976 29034
rect 14924 28970 14976 28976
rect 14936 28762 14964 28970
rect 14924 28756 14976 28762
rect 14924 28698 14976 28704
rect 14740 28552 14792 28558
rect 14740 28494 14792 28500
rect 14752 27470 14780 28494
rect 15752 27872 15804 27878
rect 15752 27814 15804 27820
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 15476 27464 15528 27470
rect 15476 27406 15528 27412
rect 14648 25356 14700 25362
rect 14648 25298 14700 25304
rect 14660 25158 14688 25298
rect 14648 25152 14700 25158
rect 14648 25094 14700 25100
rect 14556 23112 14608 23118
rect 14556 23054 14608 23060
rect 14556 21004 14608 21010
rect 14556 20946 14608 20952
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14568 19854 14596 20946
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 14016 15502 14044 19450
rect 14568 19378 14596 19790
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14660 17202 14688 25094
rect 14752 18902 14780 27406
rect 14924 26784 14976 26790
rect 14924 26726 14976 26732
rect 14936 26450 14964 26726
rect 14924 26444 14976 26450
rect 14924 26386 14976 26392
rect 15488 24206 15516 27406
rect 15660 25900 15712 25906
rect 15660 25842 15712 25848
rect 15672 24886 15700 25842
rect 15660 24880 15712 24886
rect 15660 24822 15712 24828
rect 15476 24200 15528 24206
rect 15476 24142 15528 24148
rect 15488 22710 15516 24142
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 15672 22094 15700 24822
rect 15764 24206 15792 27814
rect 15856 27062 15884 30602
rect 17144 30258 17172 31282
rect 16672 30252 16724 30258
rect 16672 30194 16724 30200
rect 17132 30252 17184 30258
rect 17132 30194 17184 30200
rect 16684 28150 16712 30194
rect 16672 28144 16724 28150
rect 16672 28086 16724 28092
rect 16488 28076 16540 28082
rect 16488 28018 16540 28024
rect 16028 28008 16080 28014
rect 16028 27950 16080 27956
rect 15844 27056 15896 27062
rect 15844 26998 15896 27004
rect 15936 27056 15988 27062
rect 15936 26998 15988 27004
rect 15752 24200 15804 24206
rect 15752 24142 15804 24148
rect 15856 23050 15884 26998
rect 15844 23044 15896 23050
rect 15844 22986 15896 22992
rect 15672 22066 15792 22094
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 14832 21956 14884 21962
rect 14832 21898 14884 21904
rect 14844 21554 14872 21898
rect 14832 21548 14884 21554
rect 14832 21490 14884 21496
rect 14844 20466 14872 21490
rect 14924 21412 14976 21418
rect 14924 21354 14976 21360
rect 14936 21010 14964 21354
rect 14924 21004 14976 21010
rect 14924 20946 14976 20952
rect 15580 20466 15608 21966
rect 15660 21616 15712 21622
rect 15660 21558 15712 21564
rect 15672 20466 15700 21558
rect 14832 20460 14884 20466
rect 14832 20402 14884 20408
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 14740 18896 14792 18902
rect 14740 18838 14792 18844
rect 14844 18748 14872 20402
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 14752 18720 14872 18748
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14108 16454 14136 16934
rect 14096 16448 14148 16454
rect 14096 16390 14148 16396
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14660 16114 14688 16390
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14752 15994 14780 18720
rect 14832 18624 14884 18630
rect 14832 18566 14884 18572
rect 14844 16182 14872 18566
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 15028 16250 15056 17070
rect 15212 16250 15240 19246
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 15200 16244 15252 16250
rect 15200 16186 15252 16192
rect 14832 16176 14884 16182
rect 14832 16118 14884 16124
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 14752 15966 14872 15994
rect 14004 15496 14056 15502
rect 14004 15438 14056 15444
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14200 14414 14228 14894
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13280 14006 13308 14214
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12912 13326 12940 13806
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 12820 12646 12848 13194
rect 12912 12850 12940 13262
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 13004 10742 13032 13126
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13280 11218 13308 12038
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 12992 10736 13044 10742
rect 12992 10678 13044 10684
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 13004 8362 13032 9522
rect 13464 8498 13492 14350
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14292 14074 14320 14214
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14188 12912 14240 12918
rect 14188 12854 14240 12860
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13648 11354 13676 12038
rect 14200 11694 14228 12854
rect 14752 12850 14780 13670
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14844 12238 14872 15966
rect 14936 14074 14964 16050
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 15028 13870 15056 16186
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15120 12986 15148 13874
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15396 12850 15424 19314
rect 15580 18426 15608 20402
rect 15672 19854 15700 20402
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15488 13938 15516 14350
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15488 12918 15516 13874
rect 15764 13530 15792 22066
rect 15948 18426 15976 26998
rect 16040 25974 16068 27950
rect 16120 27124 16172 27130
rect 16120 27066 16172 27072
rect 16132 26790 16160 27066
rect 16120 26784 16172 26790
rect 16120 26726 16172 26732
rect 16304 26784 16356 26790
rect 16304 26726 16356 26732
rect 16316 26382 16344 26726
rect 16304 26376 16356 26382
rect 16304 26318 16356 26324
rect 16028 25968 16080 25974
rect 16028 25910 16080 25916
rect 16500 25498 16528 28018
rect 16488 25492 16540 25498
rect 16488 25434 16540 25440
rect 16500 24886 16528 25434
rect 16580 25220 16632 25226
rect 16580 25162 16632 25168
rect 16488 24880 16540 24886
rect 16488 24822 16540 24828
rect 16212 22228 16264 22234
rect 16212 22170 16264 22176
rect 16224 22030 16252 22170
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 16304 22024 16356 22030
rect 16304 21966 16356 21972
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 16040 21434 16068 21490
rect 16040 21406 16252 21434
rect 16224 21350 16252 21406
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 16212 21344 16264 21350
rect 16212 21286 16264 21292
rect 16132 19854 16160 21286
rect 16316 20398 16344 21966
rect 16500 21554 16528 24822
rect 16592 22642 16620 25162
rect 16684 24410 16712 28086
rect 16764 28076 16816 28082
rect 16764 28018 16816 28024
rect 16776 25362 16804 28018
rect 17040 27872 17092 27878
rect 17040 27814 17092 27820
rect 16856 27464 16908 27470
rect 16856 27406 16908 27412
rect 16764 25356 16816 25362
rect 16764 25298 16816 25304
rect 16868 24818 16896 27406
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 16960 25838 16988 26930
rect 16948 25832 17000 25838
rect 16948 25774 17000 25780
rect 16960 25498 16988 25774
rect 16948 25492 17000 25498
rect 16948 25434 17000 25440
rect 17052 24818 17080 27814
rect 17236 27334 17264 31826
rect 17408 31816 17460 31822
rect 17408 31758 17460 31764
rect 17420 30258 17448 31758
rect 17408 30252 17460 30258
rect 17408 30194 17460 30200
rect 17420 29034 17448 30194
rect 17408 29028 17460 29034
rect 17408 28970 17460 28976
rect 17224 27328 17276 27334
rect 17224 27270 17276 27276
rect 17132 25968 17184 25974
rect 17132 25910 17184 25916
rect 17144 24954 17172 25910
rect 17132 24948 17184 24954
rect 17132 24890 17184 24896
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 16672 24404 16724 24410
rect 16672 24346 16724 24352
rect 17052 23594 17080 24754
rect 17040 23588 17092 23594
rect 17040 23530 17092 23536
rect 16856 22772 16908 22778
rect 16856 22714 16908 22720
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16868 22166 16896 22714
rect 16856 22160 16908 22166
rect 16856 22102 16908 22108
rect 16672 22092 16724 22098
rect 16672 22034 16724 22040
rect 16580 21956 16632 21962
rect 16580 21898 16632 21904
rect 16592 21622 16620 21898
rect 16580 21616 16632 21622
rect 16580 21558 16632 21564
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 16488 20868 16540 20874
rect 16488 20810 16540 20816
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 16316 19718 16344 20334
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 16500 18154 16528 20810
rect 16488 18148 16540 18154
rect 16488 18090 16540 18096
rect 16500 17542 16528 18090
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 16040 14278 16068 16050
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 16408 14618 16436 15982
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 14292 11150 14320 12174
rect 15212 12170 15240 12582
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14292 10810 14320 11086
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14292 9042 14320 9318
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 12992 8356 13044 8362
rect 12992 8298 13044 8304
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12636 7410 12664 8230
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12176 6458 12204 7142
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11716 5914 11744 6054
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 12268 5710 12296 6190
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12728 4826 12756 8026
rect 13004 5302 13032 8298
rect 14292 7954 14320 8978
rect 15120 8566 15148 11630
rect 15304 9586 15332 12174
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15108 8560 15160 8566
rect 14752 8498 14964 8514
rect 15108 8502 15160 8508
rect 14740 8492 14976 8498
rect 14792 8486 14924 8492
rect 14740 8434 14792 8440
rect 14924 8434 14976 8440
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14280 7948 14332 7954
rect 14280 7890 14332 7896
rect 14660 7478 14688 8366
rect 15120 8090 15148 8502
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15212 7886 15240 9318
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15304 7546 15332 8366
rect 15396 7970 15424 12786
rect 15488 12442 15516 12854
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15580 12442 15608 12786
rect 16040 12646 16068 14214
rect 16224 14074 16252 14350
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15488 9586 15516 12378
rect 15568 12164 15620 12170
rect 15568 12106 15620 12112
rect 15580 9654 15608 12106
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15580 8090 15608 9590
rect 16316 8974 16344 13806
rect 16500 11762 16528 17478
rect 16684 16182 16712 22034
rect 16868 20330 16896 22102
rect 17144 22094 17172 24890
rect 17236 24818 17264 27270
rect 17224 24812 17276 24818
rect 17224 24754 17276 24760
rect 17052 22066 17172 22094
rect 16948 21956 17000 21962
rect 16948 21898 17000 21904
rect 16960 20602 16988 21898
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 17052 20466 17080 22066
rect 17224 21616 17276 21622
rect 17224 21558 17276 21564
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 16856 20324 16908 20330
rect 16856 20266 16908 20272
rect 16868 18630 16896 20266
rect 17052 19786 17080 20402
rect 17236 20058 17264 21558
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 16856 18624 16908 18630
rect 16856 18566 16908 18572
rect 16856 17060 16908 17066
rect 16856 17002 16908 17008
rect 16868 16522 16896 17002
rect 16856 16516 16908 16522
rect 16856 16458 16908 16464
rect 16672 16176 16724 16182
rect 16672 16118 16724 16124
rect 16868 16130 16896 16458
rect 16868 16114 16988 16130
rect 16856 16108 16988 16114
rect 16908 16102 16988 16108
rect 16856 16050 16908 16056
rect 16856 15972 16908 15978
rect 16856 15914 16908 15920
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16684 14482 16712 15506
rect 16868 15502 16896 15914
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 16764 15428 16816 15434
rect 16764 15370 16816 15376
rect 16776 14958 16804 15370
rect 16868 15026 16896 15438
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16776 14414 16804 14894
rect 16868 14414 16896 14962
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16960 14006 16988 16102
rect 17052 15366 17080 19722
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 17236 18290 17264 18634
rect 17316 18624 17368 18630
rect 17316 18566 17368 18572
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17236 16114 17264 18226
rect 17328 17542 17356 18566
rect 17408 17672 17460 17678
rect 17408 17614 17460 17620
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 17328 16114 17356 17138
rect 17420 16998 17448 17614
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17420 16590 17448 16934
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 16960 13326 16988 13942
rect 17328 13938 17356 16050
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17328 13326 17356 13874
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 16960 12850 16988 12922
rect 17144 12850 17172 12922
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17144 12646 17172 12786
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16500 11626 16528 11698
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 17236 11286 17264 12786
rect 16396 11280 16448 11286
rect 16396 11222 16448 11228
rect 17224 11280 17276 11286
rect 17224 11222 17276 11228
rect 16408 9178 16436 11222
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16408 8974 16436 9114
rect 16500 9110 16528 9522
rect 16488 9104 16540 9110
rect 16488 9046 16540 9052
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15396 7942 15516 7970
rect 15488 7886 15516 7942
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15764 7546 15792 8570
rect 16316 8362 16344 8910
rect 16500 8430 16528 9046
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16304 8356 16356 8362
rect 16304 8298 16356 8304
rect 16500 8022 16528 8366
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 16684 7886 16712 8774
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14476 6798 14504 7346
rect 16316 6798 16344 7686
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 14476 5370 14504 6734
rect 16684 6662 16712 7822
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12728 4622 12756 4762
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12636 4146 12664 4422
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12728 3194 12756 4558
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14568 4146 14596 4422
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14108 3194 14136 4082
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14476 3194 14504 3878
rect 14752 3738 14780 4082
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 15120 3602 15148 4558
rect 17132 4004 17184 4010
rect 17132 3946 17184 3952
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16592 3602 16620 3878
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 15120 2990 15148 3538
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16868 3194 16896 3402
rect 17144 3398 17172 3946
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 15108 2984 15160 2990
rect 15108 2926 15160 2932
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 15672 2446 15700 3130
rect 17144 2446 17172 3334
rect 17236 3194 17264 9658
rect 17512 4826 17540 32422
rect 17592 32020 17644 32026
rect 17592 31962 17644 31968
rect 17604 31822 17632 31962
rect 17696 31958 17724 32778
rect 17684 31952 17736 31958
rect 17684 31894 17736 31900
rect 17592 31816 17644 31822
rect 17592 31758 17644 31764
rect 17592 26240 17644 26246
rect 17592 26182 17644 26188
rect 17604 25226 17632 26182
rect 17592 25220 17644 25226
rect 17592 25162 17644 25168
rect 17788 23254 17816 36042
rect 18708 35086 18736 36722
rect 19444 35698 19472 36790
rect 20076 36780 20128 36786
rect 20076 36722 20128 36728
rect 25136 36780 25188 36786
rect 25136 36722 25188 36728
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 18788 35692 18840 35698
rect 18788 35634 18840 35640
rect 19432 35692 19484 35698
rect 19432 35634 19484 35640
rect 18696 35080 18748 35086
rect 18696 35022 18748 35028
rect 18144 34604 18196 34610
rect 18144 34546 18196 34552
rect 18052 33992 18104 33998
rect 18052 33934 18104 33940
rect 18064 33522 18092 33934
rect 18156 33930 18184 34546
rect 18328 33992 18380 33998
rect 18328 33934 18380 33940
rect 18144 33924 18196 33930
rect 18144 33866 18196 33872
rect 18052 33516 18104 33522
rect 18052 33458 18104 33464
rect 18156 33454 18184 33866
rect 18144 33448 18196 33454
rect 18144 33390 18196 33396
rect 18156 32978 18184 33390
rect 18144 32972 18196 32978
rect 18144 32914 18196 32920
rect 18340 32502 18368 33934
rect 18708 33590 18736 35022
rect 18800 34066 18828 35634
rect 20088 35290 20116 36722
rect 25044 36712 25096 36718
rect 25044 36654 25096 36660
rect 24768 36168 24820 36174
rect 24768 36110 24820 36116
rect 22836 35760 22888 35766
rect 23112 35760 23164 35766
rect 22888 35708 23112 35714
rect 22836 35702 23164 35708
rect 21180 35692 21232 35698
rect 21180 35634 21232 35640
rect 22008 35692 22060 35698
rect 22848 35686 23152 35702
rect 23204 35692 23256 35698
rect 22008 35634 22060 35640
rect 23204 35634 23256 35640
rect 23388 35692 23440 35698
rect 23388 35634 23440 35640
rect 20536 35624 20588 35630
rect 20536 35566 20588 35572
rect 20076 35284 20128 35290
rect 20076 35226 20128 35232
rect 20352 35216 20404 35222
rect 20352 35158 20404 35164
rect 20260 35080 20312 35086
rect 20166 35048 20222 35057
rect 19064 35012 19116 35018
rect 20260 35022 20312 35028
rect 20166 34983 20168 34992
rect 19064 34954 19116 34960
rect 20220 34983 20222 34992
rect 20168 34954 20220 34960
rect 18880 34604 18932 34610
rect 18880 34546 18932 34552
rect 18892 34134 18920 34546
rect 18880 34128 18932 34134
rect 18880 34070 18932 34076
rect 18788 34060 18840 34066
rect 18788 34002 18840 34008
rect 18696 33584 18748 33590
rect 18696 33526 18748 33532
rect 18328 32496 18380 32502
rect 18328 32438 18380 32444
rect 18340 32366 18368 32438
rect 17868 32360 17920 32366
rect 17868 32302 17920 32308
rect 18328 32360 18380 32366
rect 18328 32302 18380 32308
rect 17880 32230 17908 32302
rect 17868 32224 17920 32230
rect 17868 32166 17920 32172
rect 17880 31482 17908 32166
rect 17868 31476 17920 31482
rect 17868 31418 17920 31424
rect 18236 30864 18288 30870
rect 18236 30806 18288 30812
rect 18144 30728 18196 30734
rect 18144 30670 18196 30676
rect 17960 30592 18012 30598
rect 17960 30534 18012 30540
rect 17972 30258 18000 30534
rect 18156 30326 18184 30670
rect 18144 30320 18196 30326
rect 18144 30262 18196 30268
rect 17960 30252 18012 30258
rect 17960 30194 18012 30200
rect 18156 29714 18184 30262
rect 18144 29708 18196 29714
rect 18144 29650 18196 29656
rect 18248 29646 18276 30806
rect 18420 30728 18472 30734
rect 18420 30670 18472 30676
rect 18328 30592 18380 30598
rect 18328 30534 18380 30540
rect 18236 29640 18288 29646
rect 18236 29582 18288 29588
rect 18340 29510 18368 30534
rect 18432 29850 18460 30670
rect 18708 30190 18736 33526
rect 19076 33522 19104 34954
rect 20076 34944 20128 34950
rect 20076 34886 20128 34892
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 20088 34678 20116 34886
rect 20076 34672 20128 34678
rect 20076 34614 20128 34620
rect 20272 34610 20300 35022
rect 20364 34950 20392 35158
rect 20352 34944 20404 34950
rect 20352 34886 20404 34892
rect 20364 34610 20392 34886
rect 20260 34604 20312 34610
rect 20260 34546 20312 34552
rect 20352 34604 20404 34610
rect 20352 34546 20404 34552
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19064 33516 19116 33522
rect 19064 33458 19116 33464
rect 18880 32496 18932 32502
rect 18880 32438 18932 32444
rect 18892 31278 18920 32438
rect 18880 31272 18932 31278
rect 18880 31214 18932 31220
rect 18788 30388 18840 30394
rect 18788 30330 18840 30336
rect 18696 30184 18748 30190
rect 18696 30126 18748 30132
rect 18604 30116 18656 30122
rect 18604 30058 18656 30064
rect 18420 29844 18472 29850
rect 18420 29786 18472 29792
rect 18328 29504 18380 29510
rect 18328 29446 18380 29452
rect 18616 29102 18644 30058
rect 18800 29714 18828 30330
rect 18892 30190 18920 31214
rect 19076 30394 19104 33458
rect 19340 33040 19392 33046
rect 19340 32982 19392 32988
rect 19156 32360 19208 32366
rect 19156 32302 19208 32308
rect 19064 30388 19116 30394
rect 19064 30330 19116 30336
rect 18880 30184 18932 30190
rect 18880 30126 18932 30132
rect 18788 29708 18840 29714
rect 18788 29650 18840 29656
rect 18800 29306 18828 29650
rect 18788 29300 18840 29306
rect 18788 29242 18840 29248
rect 18604 29096 18656 29102
rect 18604 29038 18656 29044
rect 18420 28552 18472 28558
rect 18420 28494 18472 28500
rect 18144 27600 18196 27606
rect 18144 27542 18196 27548
rect 18052 27328 18104 27334
rect 18052 27270 18104 27276
rect 18064 27062 18092 27270
rect 18156 27130 18184 27542
rect 18432 27334 18460 28494
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18420 27328 18472 27334
rect 18420 27270 18472 27276
rect 18432 27130 18460 27270
rect 18144 27124 18196 27130
rect 18144 27066 18196 27072
rect 18420 27124 18472 27130
rect 18420 27066 18472 27072
rect 18052 27056 18104 27062
rect 18052 26998 18104 27004
rect 18432 26790 18460 27066
rect 18420 26784 18472 26790
rect 18420 26726 18472 26732
rect 17868 25900 17920 25906
rect 17868 25842 17920 25848
rect 17880 25498 17908 25842
rect 17868 25492 17920 25498
rect 17868 25434 17920 25440
rect 18524 25294 18552 27406
rect 18696 27396 18748 27402
rect 18696 27338 18748 27344
rect 18052 25288 18104 25294
rect 18052 25230 18104 25236
rect 18512 25288 18564 25294
rect 18512 25230 18564 25236
rect 17776 23248 17828 23254
rect 17776 23190 17828 23196
rect 17592 23044 17644 23050
rect 17592 22986 17644 22992
rect 17604 22710 17632 22986
rect 17592 22704 17644 22710
rect 17592 22646 17644 22652
rect 17604 21962 17632 22646
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 17592 21956 17644 21962
rect 17592 21898 17644 21904
rect 17604 21010 17632 21898
rect 17972 21622 18000 22374
rect 17960 21616 18012 21622
rect 17960 21558 18012 21564
rect 18064 21350 18092 25230
rect 18708 24818 18736 27338
rect 18696 24812 18748 24818
rect 18696 24754 18748 24760
rect 18892 22710 18920 30126
rect 19168 29170 19196 32302
rect 19248 31272 19300 31278
rect 19248 31214 19300 31220
rect 19260 30802 19288 31214
rect 19248 30796 19300 30802
rect 19248 30738 19300 30744
rect 19352 29646 19380 32982
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 20548 31346 20576 35566
rect 20628 35284 20680 35290
rect 20628 35226 20680 35232
rect 20640 34610 20668 35226
rect 20720 35216 20772 35222
rect 20720 35158 20772 35164
rect 20628 34604 20680 34610
rect 20628 34546 20680 34552
rect 20640 34066 20668 34546
rect 20732 34202 20760 35158
rect 21192 35086 21220 35634
rect 20812 35080 20864 35086
rect 20810 35048 20812 35057
rect 21180 35080 21232 35086
rect 20864 35048 20866 35057
rect 21180 35022 21232 35028
rect 21916 35080 21968 35086
rect 21916 35022 21968 35028
rect 20810 34983 20866 34992
rect 21192 34678 21220 35022
rect 21180 34672 21232 34678
rect 21180 34614 21232 34620
rect 20720 34196 20772 34202
rect 20720 34138 20772 34144
rect 20628 34060 20680 34066
rect 20628 34002 20680 34008
rect 20640 33590 20668 34002
rect 20628 33584 20680 33590
rect 20628 33526 20680 33532
rect 20812 32428 20864 32434
rect 20812 32370 20864 32376
rect 20720 31408 20772 31414
rect 20720 31350 20772 31356
rect 19984 31340 20036 31346
rect 19984 31282 20036 31288
rect 20536 31340 20588 31346
rect 20536 31282 20588 31288
rect 19996 30870 20024 31282
rect 20260 31272 20312 31278
rect 20260 31214 20312 31220
rect 19984 30864 20036 30870
rect 19984 30806 20036 30812
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 20272 30190 20300 31214
rect 20732 30666 20760 31350
rect 20824 30802 20852 32370
rect 21192 30870 21220 34614
rect 21364 34604 21416 34610
rect 21364 34546 21416 34552
rect 21376 33998 21404 34546
rect 21548 34400 21600 34406
rect 21548 34342 21600 34348
rect 21560 34134 21588 34342
rect 21548 34128 21600 34134
rect 21548 34070 21600 34076
rect 21364 33992 21416 33998
rect 21364 33934 21416 33940
rect 21272 32768 21324 32774
rect 21272 32710 21324 32716
rect 21284 32434 21312 32710
rect 21376 32502 21404 33934
rect 21364 32496 21416 32502
rect 21364 32438 21416 32444
rect 21272 32428 21324 32434
rect 21272 32370 21324 32376
rect 21180 30864 21232 30870
rect 21180 30806 21232 30812
rect 20812 30796 20864 30802
rect 20812 30738 20864 30744
rect 20720 30660 20772 30666
rect 20720 30602 20772 30608
rect 20732 30394 20760 30602
rect 20720 30388 20772 30394
rect 20720 30330 20772 30336
rect 20824 30274 20852 30738
rect 20904 30728 20956 30734
rect 20904 30670 20956 30676
rect 20732 30258 20852 30274
rect 20720 30252 20852 30258
rect 20772 30246 20852 30252
rect 20720 30194 20772 30200
rect 20260 30184 20312 30190
rect 20260 30126 20312 30132
rect 19984 29776 20036 29782
rect 19984 29718 20036 29724
rect 20168 29776 20220 29782
rect 20168 29718 20220 29724
rect 19996 29646 20024 29718
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19432 29300 19484 29306
rect 19432 29242 19484 29248
rect 19156 29164 19208 29170
rect 19156 29106 19208 29112
rect 19168 28490 19196 29106
rect 19248 29096 19300 29102
rect 19248 29038 19300 29044
rect 19260 28762 19288 29038
rect 19340 28960 19392 28966
rect 19340 28902 19392 28908
rect 19248 28756 19300 28762
rect 19248 28698 19300 28704
rect 19156 28484 19208 28490
rect 19156 28426 19208 28432
rect 19352 27334 19380 28902
rect 19444 27606 19472 29242
rect 19996 28762 20024 29582
rect 20076 29572 20128 29578
rect 20076 29514 20128 29520
rect 20088 29102 20116 29514
rect 20076 29096 20128 29102
rect 20076 29038 20128 29044
rect 20180 29034 20208 29718
rect 20272 29306 20300 30126
rect 20352 29572 20404 29578
rect 20352 29514 20404 29520
rect 20260 29300 20312 29306
rect 20260 29242 20312 29248
rect 20364 29170 20392 29514
rect 20732 29322 20760 30194
rect 20916 29714 20944 30670
rect 21284 30258 21312 32370
rect 21272 30252 21324 30258
rect 21272 30194 21324 30200
rect 20904 29708 20956 29714
rect 20904 29650 20956 29656
rect 20548 29294 20760 29322
rect 20352 29164 20404 29170
rect 20352 29106 20404 29112
rect 20168 29028 20220 29034
rect 20168 28970 20220 28976
rect 20444 29028 20496 29034
rect 20444 28970 20496 28976
rect 19984 28756 20036 28762
rect 19984 28698 20036 28704
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19996 28218 20024 28698
rect 20180 28642 20208 28970
rect 20456 28762 20484 28970
rect 20444 28756 20496 28762
rect 20444 28698 20496 28704
rect 20180 28614 20484 28642
rect 19984 28212 20036 28218
rect 19984 28154 20036 28160
rect 19432 27600 19484 27606
rect 19432 27542 19484 27548
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19352 26874 19380 27270
rect 19444 26994 19472 27542
rect 19996 27470 20024 28154
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19432 26988 19484 26994
rect 19432 26930 19484 26936
rect 19616 26920 19668 26926
rect 19352 26868 19616 26874
rect 19352 26862 19668 26868
rect 19352 26846 19656 26862
rect 19996 26314 20024 27406
rect 20076 26852 20128 26858
rect 20076 26794 20128 26800
rect 19984 26308 20036 26314
rect 19984 26250 20036 26256
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19340 26036 19392 26042
rect 19340 25978 19392 25984
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 19260 25106 19288 25230
rect 19352 25226 19380 25978
rect 20088 25242 20116 26794
rect 20260 26512 20312 26518
rect 20260 26454 20312 26460
rect 20272 25786 20300 26454
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 20456 26330 20484 28614
rect 20548 26518 20576 29294
rect 20628 29164 20680 29170
rect 20628 29106 20680 29112
rect 20640 27402 20668 29106
rect 21284 29102 21312 30194
rect 21272 29096 21324 29102
rect 21272 29038 21324 29044
rect 20628 27396 20680 27402
rect 20628 27338 20680 27344
rect 20536 26512 20588 26518
rect 20536 26454 20588 26460
rect 20640 26450 20668 27338
rect 20628 26444 20680 26450
rect 20628 26386 20680 26392
rect 20364 26042 20392 26318
rect 20456 26302 20668 26330
rect 20536 26246 20588 26252
rect 20536 26188 20588 26194
rect 20352 26036 20404 26042
rect 20352 25978 20404 25984
rect 20180 25758 20300 25786
rect 20180 25362 20208 25758
rect 20260 25696 20312 25702
rect 20260 25638 20312 25644
rect 20168 25356 20220 25362
rect 20168 25298 20220 25304
rect 20272 25294 20300 25638
rect 20260 25288 20312 25294
rect 19340 25220 19392 25226
rect 20088 25214 20208 25242
rect 20260 25230 20312 25236
rect 19340 25162 19392 25168
rect 20076 25152 20128 25158
rect 19260 25078 19380 25106
rect 20076 25094 20128 25100
rect 19352 24886 19380 25078
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19340 24880 19392 24886
rect 19340 24822 19392 24828
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19800 23656 19852 23662
rect 19800 23598 19852 23604
rect 19812 23186 19840 23598
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 19800 23180 19852 23186
rect 19800 23122 19852 23128
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 18880 22704 18932 22710
rect 18880 22646 18932 22652
rect 19064 22636 19116 22642
rect 19064 22578 19116 22584
rect 18880 22500 18932 22506
rect 18880 22442 18932 22448
rect 18788 22432 18840 22438
rect 18788 22374 18840 22380
rect 18328 21888 18380 21894
rect 18328 21830 18380 21836
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 18064 20262 18092 21286
rect 18340 20602 18368 21830
rect 18328 20596 18380 20602
rect 18328 20538 18380 20544
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17604 18290 17632 18566
rect 17880 18358 17908 18702
rect 17868 18352 17920 18358
rect 17868 18294 17920 18300
rect 17592 18284 17644 18290
rect 17592 18226 17644 18232
rect 17604 15570 17632 18226
rect 17880 17678 17908 18294
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 18156 17338 18184 19110
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17696 16182 17724 16526
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 17684 16176 17736 16182
rect 17684 16118 17736 16124
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17592 15564 17644 15570
rect 17592 15506 17644 15512
rect 17880 15026 17908 16050
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17972 14482 18000 16458
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17972 13938 18000 14418
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 17868 8560 17920 8566
rect 17868 8502 17920 8508
rect 17880 5234 17908 8502
rect 18064 7546 18092 17206
rect 18340 17202 18368 20538
rect 18800 19378 18828 22374
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18512 18896 18564 18902
rect 18512 18838 18564 18844
rect 18524 18290 18552 18838
rect 18696 18692 18748 18698
rect 18696 18634 18748 18640
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18432 17134 18460 17478
rect 18420 17128 18472 17134
rect 18420 17070 18472 17076
rect 18524 16114 18552 18226
rect 18616 16522 18644 18226
rect 18708 17678 18736 18634
rect 18892 18358 18920 22442
rect 19076 22234 19104 22578
rect 19064 22228 19116 22234
rect 19064 22170 19116 22176
rect 19352 22098 19380 23054
rect 19996 22982 20024 23462
rect 20088 23186 20116 25094
rect 20180 23254 20208 25214
rect 20444 24880 20496 24886
rect 20444 24822 20496 24828
rect 20260 23724 20312 23730
rect 20260 23666 20312 23672
rect 20168 23248 20220 23254
rect 20168 23190 20220 23196
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 19984 22976 20036 22982
rect 19984 22918 20036 22924
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19996 22710 20024 22918
rect 19984 22704 20036 22710
rect 19984 22646 20036 22652
rect 19984 22432 20036 22438
rect 19984 22374 20036 22380
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19996 22030 20024 22374
rect 20272 22030 20300 23666
rect 20352 23316 20404 23322
rect 20352 23258 20404 23264
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19984 22024 20036 22030
rect 19984 21966 20036 21972
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19352 20534 19380 21286
rect 19444 20602 19472 21966
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19444 19922 19472 20538
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 18880 18352 18932 18358
rect 18880 18294 18932 18300
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18604 16516 18656 16522
rect 18604 16458 18656 16464
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 18524 15026 18552 16050
rect 18708 15570 18736 17138
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18524 14482 18552 14962
rect 18512 14476 18564 14482
rect 18512 14418 18564 14424
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18616 14074 18644 14350
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 18524 13326 18552 13874
rect 18616 13326 18644 14010
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18708 12850 18736 15506
rect 19260 15502 19288 17614
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19156 15496 19208 15502
rect 19156 15438 19208 15444
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19168 15026 19196 15438
rect 19156 15020 19208 15026
rect 19156 14962 19208 14968
rect 19064 14544 19116 14550
rect 19064 14486 19116 14492
rect 19076 13190 19104 14486
rect 19168 13938 19196 14962
rect 19260 14890 19288 15438
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19168 13394 19196 13874
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19260 13326 19288 14826
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 18708 12434 18736 12786
rect 18892 12646 18920 12854
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18524 12406 18736 12434
rect 18524 12238 18552 12406
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18236 11620 18288 11626
rect 18236 11562 18288 11568
rect 18248 10742 18276 11562
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 18524 8974 18552 12174
rect 18984 9178 19012 12786
rect 19076 12306 19104 13126
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19168 12442 19196 12786
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 19260 12170 19288 12582
rect 19248 12164 19300 12170
rect 19248 12106 19300 12112
rect 19352 10130 19380 14758
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19984 13456 20036 13462
rect 19984 13398 20036 13404
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19444 12850 19472 13126
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19996 12238 20024 13398
rect 20180 12434 20208 20402
rect 20272 18834 20300 21966
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 20364 17218 20392 23258
rect 20456 22642 20484 24822
rect 20548 23730 20576 26188
rect 20640 25362 20668 26302
rect 21284 25838 21312 29038
rect 21560 26382 21588 34070
rect 21928 33998 21956 35022
rect 22020 34610 22048 35634
rect 22652 35624 22704 35630
rect 22652 35566 22704 35572
rect 22664 35290 22692 35566
rect 23216 35290 23244 35634
rect 22652 35284 22704 35290
rect 22652 35226 22704 35232
rect 23204 35284 23256 35290
rect 23204 35226 23256 35232
rect 23400 35154 23428 35634
rect 24780 35630 24808 36110
rect 23756 35624 23808 35630
rect 23756 35566 23808 35572
rect 24768 35624 24820 35630
rect 24768 35566 24820 35572
rect 24952 35624 25004 35630
rect 24952 35566 25004 35572
rect 23480 35556 23532 35562
rect 23480 35498 23532 35504
rect 23388 35148 23440 35154
rect 23388 35090 23440 35096
rect 23492 35086 23520 35498
rect 22468 35080 22520 35086
rect 22468 35022 22520 35028
rect 22652 35080 22704 35086
rect 22652 35022 22704 35028
rect 23296 35080 23348 35086
rect 23296 35022 23348 35028
rect 23480 35080 23532 35086
rect 23480 35022 23532 35028
rect 22480 34950 22508 35022
rect 22468 34944 22520 34950
rect 22468 34886 22520 34892
rect 22664 34746 22692 35022
rect 23308 34950 23336 35022
rect 23296 34944 23348 34950
rect 23296 34886 23348 34892
rect 22652 34740 22704 34746
rect 22652 34682 22704 34688
rect 22008 34604 22060 34610
rect 22008 34546 22060 34552
rect 23308 34542 23336 34886
rect 23768 34678 23796 35566
rect 24216 35556 24268 35562
rect 24216 35498 24268 35504
rect 23756 34672 23808 34678
rect 23756 34614 23808 34620
rect 24228 34610 24256 35498
rect 24492 35012 24544 35018
rect 24492 34954 24544 34960
rect 24768 35012 24820 35018
rect 24768 34954 24820 34960
rect 24504 34610 24532 34954
rect 24676 34944 24728 34950
rect 24676 34886 24728 34892
rect 24688 34610 24716 34886
rect 24216 34604 24268 34610
rect 24216 34546 24268 34552
rect 24492 34604 24544 34610
rect 24492 34546 24544 34552
rect 24676 34604 24728 34610
rect 24676 34546 24728 34552
rect 22100 34536 22152 34542
rect 22100 34478 22152 34484
rect 23296 34536 23348 34542
rect 23296 34478 23348 34484
rect 22112 34082 22140 34478
rect 24228 34474 24256 34546
rect 22192 34468 22244 34474
rect 22192 34410 22244 34416
rect 24216 34468 24268 34474
rect 24216 34410 24268 34416
rect 22020 34054 22140 34082
rect 21916 33992 21968 33998
rect 21916 33934 21968 33940
rect 22020 32774 22048 34054
rect 22204 33998 22232 34410
rect 24780 34066 24808 34954
rect 24768 34060 24820 34066
rect 24768 34002 24820 34008
rect 22192 33992 22244 33998
rect 22192 33934 22244 33940
rect 23020 33924 23072 33930
rect 23020 33866 23072 33872
rect 23032 32910 23060 33866
rect 24780 33114 24808 34002
rect 24964 33998 24992 35566
rect 25056 35290 25084 36654
rect 25148 35834 25176 36722
rect 25136 35828 25188 35834
rect 25136 35770 25188 35776
rect 25240 35766 25268 37062
rect 25504 36780 25556 36786
rect 25504 36722 25556 36728
rect 26148 36780 26200 36786
rect 26148 36722 26200 36728
rect 31024 36780 31076 36786
rect 31024 36722 31076 36728
rect 25228 35760 25280 35766
rect 25228 35702 25280 35708
rect 25516 35630 25544 36722
rect 26056 36644 26108 36650
rect 26056 36586 26108 36592
rect 25872 36576 25924 36582
rect 25872 36518 25924 36524
rect 25884 36242 25912 36518
rect 26068 36242 26096 36586
rect 26160 36378 26188 36722
rect 30104 36576 30156 36582
rect 30104 36518 30156 36524
rect 26148 36372 26200 36378
rect 26148 36314 26200 36320
rect 25872 36236 25924 36242
rect 25872 36178 25924 36184
rect 26056 36236 26108 36242
rect 26056 36178 26108 36184
rect 26160 36106 26188 36314
rect 29092 36168 29144 36174
rect 29092 36110 29144 36116
rect 26148 36100 26200 36106
rect 26148 36042 26200 36048
rect 25504 35624 25556 35630
rect 25504 35566 25556 35572
rect 29000 35624 29052 35630
rect 29104 35612 29132 36110
rect 29460 36100 29512 36106
rect 29460 36042 29512 36048
rect 29184 36032 29236 36038
rect 29184 35974 29236 35980
rect 29052 35584 29132 35612
rect 29000 35566 29052 35572
rect 25516 35494 25544 35566
rect 25504 35488 25556 35494
rect 25504 35430 25556 35436
rect 25044 35284 25096 35290
rect 25044 35226 25096 35232
rect 29012 35154 29040 35566
rect 29000 35148 29052 35154
rect 29000 35090 29052 35096
rect 29196 35086 29224 35974
rect 29472 35698 29500 36042
rect 29460 35692 29512 35698
rect 29460 35634 29512 35640
rect 25780 35080 25832 35086
rect 25780 35022 25832 35028
rect 26792 35080 26844 35086
rect 26792 35022 26844 35028
rect 29184 35080 29236 35086
rect 29184 35022 29236 35028
rect 25044 34672 25096 34678
rect 25044 34614 25096 34620
rect 24952 33992 25004 33998
rect 24952 33934 25004 33940
rect 25056 33658 25084 34614
rect 25688 34400 25740 34406
rect 25688 34342 25740 34348
rect 25700 33998 25728 34342
rect 25688 33992 25740 33998
rect 25688 33934 25740 33940
rect 25044 33652 25096 33658
rect 25044 33594 25096 33600
rect 25412 33448 25464 33454
rect 25412 33390 25464 33396
rect 24952 33380 25004 33386
rect 24952 33322 25004 33328
rect 24768 33108 24820 33114
rect 24768 33050 24820 33056
rect 23112 33040 23164 33046
rect 23112 32982 23164 32988
rect 23020 32904 23072 32910
rect 23020 32846 23072 32852
rect 22008 32768 22060 32774
rect 22008 32710 22060 32716
rect 23032 32502 23060 32846
rect 23020 32496 23072 32502
rect 23020 32438 23072 32444
rect 23124 32434 23152 32982
rect 24860 32904 24912 32910
rect 24860 32846 24912 32852
rect 23388 32496 23440 32502
rect 23388 32438 23440 32444
rect 23112 32428 23164 32434
rect 23112 32370 23164 32376
rect 23124 31890 23152 32370
rect 23204 32020 23256 32026
rect 23204 31962 23256 31968
rect 23112 31884 23164 31890
rect 23112 31826 23164 31832
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22296 30326 22324 31282
rect 23216 31210 23244 31962
rect 23400 31958 23428 32438
rect 24872 32026 24900 32846
rect 24964 32502 24992 33322
rect 25424 33046 25452 33390
rect 25792 33114 25820 35022
rect 26424 34536 26476 34542
rect 26424 34478 26476 34484
rect 26436 33998 26464 34478
rect 26804 34134 26832 35022
rect 26792 34128 26844 34134
rect 26792 34070 26844 34076
rect 26424 33992 26476 33998
rect 26424 33934 26476 33940
rect 26148 33924 26200 33930
rect 26148 33866 26200 33872
rect 27252 33924 27304 33930
rect 27252 33866 27304 33872
rect 25964 33448 26016 33454
rect 25964 33390 26016 33396
rect 25780 33108 25832 33114
rect 25780 33050 25832 33056
rect 25412 33040 25464 33046
rect 25412 32982 25464 32988
rect 25976 32910 26004 33390
rect 26160 33130 26188 33866
rect 26424 33516 26476 33522
rect 26424 33458 26476 33464
rect 26160 33102 26280 33130
rect 26252 33046 26280 33102
rect 26148 33040 26200 33046
rect 26148 32982 26200 32988
rect 26240 33040 26292 33046
rect 26240 32982 26292 32988
rect 26160 32910 26188 32982
rect 25320 32904 25372 32910
rect 25320 32846 25372 32852
rect 25964 32904 26016 32910
rect 25964 32846 26016 32852
rect 26148 32904 26200 32910
rect 26148 32846 26200 32852
rect 24952 32496 25004 32502
rect 24952 32438 25004 32444
rect 24860 32020 24912 32026
rect 24860 31962 24912 31968
rect 23388 31952 23440 31958
rect 23388 31894 23440 31900
rect 23572 31340 23624 31346
rect 23572 31282 23624 31288
rect 23204 31204 23256 31210
rect 23204 31146 23256 31152
rect 22376 31136 22428 31142
rect 22376 31078 22428 31084
rect 22284 30320 22336 30326
rect 22284 30262 22336 30268
rect 22100 29776 22152 29782
rect 22100 29718 22152 29724
rect 22112 27946 22140 29718
rect 22192 28076 22244 28082
rect 22192 28018 22244 28024
rect 22100 27940 22152 27946
rect 22100 27882 22152 27888
rect 22204 27130 22232 28018
rect 22192 27124 22244 27130
rect 22192 27066 22244 27072
rect 22100 26988 22152 26994
rect 22100 26930 22152 26936
rect 21364 26376 21416 26382
rect 21364 26318 21416 26324
rect 21548 26376 21600 26382
rect 21548 26318 21600 26324
rect 21272 25832 21324 25838
rect 21272 25774 21324 25780
rect 20628 25356 20680 25362
rect 20628 25298 20680 25304
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 20536 23588 20588 23594
rect 20536 23530 20588 23536
rect 20548 22930 20576 23530
rect 20640 23322 20668 25298
rect 20720 24132 20772 24138
rect 20720 24074 20772 24080
rect 20628 23316 20680 23322
rect 20628 23258 20680 23264
rect 20640 23118 20668 23258
rect 20628 23112 20680 23118
rect 20628 23054 20680 23060
rect 20548 22902 20668 22930
rect 20640 22778 20668 22902
rect 20628 22772 20680 22778
rect 20628 22714 20680 22720
rect 20444 22636 20496 22642
rect 20444 22578 20496 22584
rect 20456 21622 20484 22578
rect 20444 21616 20496 21622
rect 20444 21558 20496 21564
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20548 20058 20576 20402
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20640 17678 20668 22714
rect 20732 21690 20760 24074
rect 21376 23798 21404 26318
rect 22008 26240 22060 26246
rect 22008 26182 22060 26188
rect 21364 23792 21416 23798
rect 21364 23734 21416 23740
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 20720 21684 20772 21690
rect 20720 21626 20772 21632
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 20824 21486 20852 21626
rect 20812 21480 20864 21486
rect 20812 21422 20864 21428
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20812 20528 20864 20534
rect 20812 20470 20864 20476
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 20364 17190 20576 17218
rect 20260 15428 20312 15434
rect 20260 15370 20312 15376
rect 20272 14414 20300 15370
rect 20260 14408 20312 14414
rect 20260 14350 20312 14356
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20352 14340 20404 14346
rect 20352 14282 20404 14288
rect 20180 12406 20300 12434
rect 19524 12232 19576 12238
rect 19444 12180 19524 12186
rect 19444 12174 19576 12180
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19444 12158 19564 12174
rect 20168 12164 20220 12170
rect 19444 11354 19472 12158
rect 20168 12106 20220 12112
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19260 9586 19288 9998
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19352 9466 19380 10066
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 19444 9654 19472 9862
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19260 9438 19380 9466
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 18616 8974 18644 9114
rect 18880 9036 18932 9042
rect 18880 8978 18932 8984
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18248 8634 18276 8910
rect 18328 8900 18380 8906
rect 18380 8860 18460 8888
rect 18328 8842 18380 8848
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18432 8566 18460 8860
rect 18420 8560 18472 8566
rect 18420 8502 18472 8508
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 18524 8090 18552 8230
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18892 7750 18920 8978
rect 19260 7886 19288 9438
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19352 8498 19380 9318
rect 19996 8906 20024 10542
rect 20180 9994 20208 12106
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 20180 9722 20208 9930
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20272 9382 20300 12406
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 19432 8900 19484 8906
rect 19432 8842 19484 8848
rect 19984 8900 20036 8906
rect 19984 8842 20036 8848
rect 19444 8634 19472 8842
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 18432 6390 18460 7686
rect 18892 6458 18920 7686
rect 19352 7546 19380 8434
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 18420 6384 18472 6390
rect 18420 6326 18472 6332
rect 19352 5302 19380 7346
rect 19444 6118 19472 7822
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 20088 7478 20116 8774
rect 20364 8634 20392 14282
rect 20456 13462 20484 14350
rect 20444 13456 20496 13462
rect 20444 13398 20496 13404
rect 20444 13252 20496 13258
rect 20444 13194 20496 13200
rect 20456 9738 20484 13194
rect 20548 12306 20576 17190
rect 20732 16590 20760 20402
rect 20824 20058 20852 20470
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20916 19854 20944 21286
rect 21008 20602 21036 23054
rect 21088 22704 21140 22710
rect 21088 22646 21140 22652
rect 21100 21894 21128 22646
rect 21916 21956 21968 21962
rect 21916 21898 21968 21904
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 21364 21888 21416 21894
rect 21364 21830 21416 21836
rect 21456 21888 21508 21894
rect 21456 21830 21508 21836
rect 21272 21548 21324 21554
rect 21272 21490 21324 21496
rect 20996 20596 21048 20602
rect 20996 20538 21048 20544
rect 21284 20534 21312 21490
rect 21272 20528 21324 20534
rect 21272 20470 21324 20476
rect 21376 19854 21404 21830
rect 21468 21690 21496 21830
rect 21456 21684 21508 21690
rect 21456 21626 21508 21632
rect 21548 21548 21600 21554
rect 21548 21490 21600 21496
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 21272 19848 21324 19854
rect 21272 19790 21324 19796
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21180 19780 21232 19786
rect 21180 19722 21232 19728
rect 20812 18080 20864 18086
rect 20812 18022 20864 18028
rect 20824 17610 20852 18022
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20824 13326 20852 17546
rect 21192 17202 21220 19722
rect 21180 17196 21232 17202
rect 21180 17138 21232 17144
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 21100 16590 21128 16934
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 20916 15094 20944 16526
rect 21284 16250 21312 19790
rect 21468 19786 21496 20402
rect 21456 19780 21508 19786
rect 21456 19722 21508 19728
rect 21560 17814 21588 21490
rect 21640 20528 21692 20534
rect 21640 20470 21692 20476
rect 21652 19854 21680 20470
rect 21640 19848 21692 19854
rect 21640 19790 21692 19796
rect 21928 18698 21956 21898
rect 22020 20058 22048 26182
rect 22008 20052 22060 20058
rect 22008 19994 22060 20000
rect 22112 19514 22140 26930
rect 22296 25294 22324 30262
rect 22388 30190 22416 31078
rect 22376 30184 22428 30190
rect 22376 30126 22428 30132
rect 22388 29238 22416 30126
rect 23584 29782 23612 31282
rect 24308 30252 24360 30258
rect 24308 30194 24360 30200
rect 24952 30252 25004 30258
rect 24952 30194 25004 30200
rect 23940 30048 23992 30054
rect 23940 29990 23992 29996
rect 23572 29776 23624 29782
rect 23572 29718 23624 29724
rect 23480 29640 23532 29646
rect 23480 29582 23532 29588
rect 23388 29572 23440 29578
rect 23388 29514 23440 29520
rect 22836 29504 22888 29510
rect 22836 29446 22888 29452
rect 22376 29232 22428 29238
rect 22376 29174 22428 29180
rect 22848 29034 22876 29446
rect 22836 29028 22888 29034
rect 22836 28970 22888 28976
rect 22376 28960 22428 28966
rect 22376 28902 22428 28908
rect 22388 28082 22416 28902
rect 22744 28552 22796 28558
rect 22744 28494 22796 28500
rect 22560 28416 22612 28422
rect 22560 28358 22612 28364
rect 22572 28150 22600 28358
rect 22560 28144 22612 28150
rect 22560 28086 22612 28092
rect 22376 28076 22428 28082
rect 22376 28018 22428 28024
rect 22756 27538 22784 28494
rect 22744 27532 22796 27538
rect 22744 27474 22796 27480
rect 22468 27464 22520 27470
rect 22468 27406 22520 27412
rect 22376 26988 22428 26994
rect 22376 26930 22428 26936
rect 22388 26382 22416 26930
rect 22480 26382 22508 27406
rect 23400 27130 23428 29514
rect 23388 27124 23440 27130
rect 23388 27066 23440 27072
rect 23492 26926 23520 29582
rect 23584 28558 23612 29718
rect 23952 29714 23980 29990
rect 23756 29708 23808 29714
rect 23756 29650 23808 29656
rect 23940 29708 23992 29714
rect 23940 29650 23992 29656
rect 23664 29640 23716 29646
rect 23664 29582 23716 29588
rect 23676 29238 23704 29582
rect 23768 29306 23796 29650
rect 23848 29640 23900 29646
rect 23848 29582 23900 29588
rect 23756 29300 23808 29306
rect 23756 29242 23808 29248
rect 23664 29232 23716 29238
rect 23664 29174 23716 29180
rect 23860 29186 23888 29582
rect 23952 29306 23980 29650
rect 23940 29300 23992 29306
rect 23940 29242 23992 29248
rect 23860 29158 23980 29186
rect 23952 29102 23980 29158
rect 23940 29096 23992 29102
rect 23940 29038 23992 29044
rect 24032 29096 24084 29102
rect 24032 29038 24084 29044
rect 23952 28762 23980 29038
rect 23940 28756 23992 28762
rect 23940 28698 23992 28704
rect 23572 28552 23624 28558
rect 23572 28494 23624 28500
rect 23480 26920 23532 26926
rect 23480 26862 23532 26868
rect 23492 26450 23520 26862
rect 23480 26444 23532 26450
rect 23480 26386 23532 26392
rect 22376 26376 22428 26382
rect 22376 26318 22428 26324
rect 22468 26376 22520 26382
rect 22468 26318 22520 26324
rect 23584 26234 23612 28494
rect 24044 27470 24072 29038
rect 24320 29034 24348 30194
rect 24964 29850 24992 30194
rect 25332 30190 25360 32846
rect 26160 32570 26188 32846
rect 26436 32842 26464 33458
rect 27264 32910 27292 33866
rect 28908 33584 28960 33590
rect 28908 33526 28960 33532
rect 27896 33516 27948 33522
rect 27896 33458 27948 33464
rect 27436 33312 27488 33318
rect 27436 33254 27488 33260
rect 27448 32910 27476 33254
rect 27908 33114 27936 33458
rect 27896 33108 27948 33114
rect 27896 33050 27948 33056
rect 27160 32904 27212 32910
rect 27160 32846 27212 32852
rect 27252 32904 27304 32910
rect 27252 32846 27304 32852
rect 27436 32904 27488 32910
rect 27436 32846 27488 32852
rect 27528 32904 27580 32910
rect 27528 32846 27580 32852
rect 28080 32904 28132 32910
rect 28080 32846 28132 32852
rect 28632 32904 28684 32910
rect 28632 32846 28684 32852
rect 26424 32836 26476 32842
rect 26424 32778 26476 32784
rect 26148 32564 26200 32570
rect 26148 32506 26200 32512
rect 26436 32298 26464 32778
rect 26424 32292 26476 32298
rect 26424 32234 26476 32240
rect 27172 31822 27200 32846
rect 27264 32774 27292 32846
rect 27252 32768 27304 32774
rect 27252 32710 27304 32716
rect 27540 32570 27568 32846
rect 27804 32768 27856 32774
rect 27804 32710 27856 32716
rect 27528 32564 27580 32570
rect 27528 32506 27580 32512
rect 27344 32428 27396 32434
rect 27344 32370 27396 32376
rect 27160 31816 27212 31822
rect 27160 31758 27212 31764
rect 25320 30184 25372 30190
rect 25320 30126 25372 30132
rect 25964 30184 26016 30190
rect 25964 30126 26016 30132
rect 24952 29844 25004 29850
rect 24952 29786 25004 29792
rect 24584 29708 24636 29714
rect 24584 29650 24636 29656
rect 24492 29096 24544 29102
rect 24490 29064 24492 29073
rect 24544 29064 24546 29073
rect 24308 29028 24360 29034
rect 24490 28999 24546 29008
rect 24308 28970 24360 28976
rect 24400 28552 24452 28558
rect 24400 28494 24452 28500
rect 24412 28082 24440 28494
rect 24400 28076 24452 28082
rect 24400 28018 24452 28024
rect 24412 27538 24440 28018
rect 24400 27532 24452 27538
rect 24400 27474 24452 27480
rect 24032 27464 24084 27470
rect 24032 27406 24084 27412
rect 24216 26988 24268 26994
rect 24216 26930 24268 26936
rect 24228 26518 24256 26930
rect 24216 26512 24268 26518
rect 24216 26454 24268 26460
rect 23756 26444 23808 26450
rect 23756 26386 23808 26392
rect 23584 26206 23704 26234
rect 23572 25832 23624 25838
rect 23572 25774 23624 25780
rect 22284 25288 22336 25294
rect 22284 25230 22336 25236
rect 22296 24886 22324 25230
rect 23480 25220 23532 25226
rect 23480 25162 23532 25168
rect 22284 24880 22336 24886
rect 22284 24822 22336 24828
rect 22376 24812 22428 24818
rect 22376 24754 22428 24760
rect 22836 24812 22888 24818
rect 22836 24754 22888 24760
rect 22928 24812 22980 24818
rect 22928 24754 22980 24760
rect 22192 24132 22244 24138
rect 22192 24074 22244 24080
rect 22204 23118 22232 24074
rect 22192 23112 22244 23118
rect 22192 23054 22244 23060
rect 22388 21486 22416 24754
rect 22848 24410 22876 24754
rect 22836 24404 22888 24410
rect 22836 24346 22888 24352
rect 22652 24200 22704 24206
rect 22652 24142 22704 24148
rect 22468 24132 22520 24138
rect 22468 24074 22520 24080
rect 22480 23866 22508 24074
rect 22468 23860 22520 23866
rect 22468 23802 22520 23808
rect 22560 22976 22612 22982
rect 22560 22918 22612 22924
rect 22572 22094 22600 22918
rect 22480 22066 22600 22094
rect 22376 21480 22428 21486
rect 22376 21422 22428 21428
rect 22192 19984 22244 19990
rect 22192 19926 22244 19932
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 21916 18692 21968 18698
rect 21916 18634 21968 18640
rect 21548 17808 21600 17814
rect 21548 17750 21600 17756
rect 21560 17202 21588 17750
rect 21928 17610 21956 18634
rect 22020 17882 22048 19314
rect 22204 18698 22232 19926
rect 22388 18766 22416 21422
rect 22480 19922 22508 22066
rect 22664 21570 22692 24142
rect 22744 24064 22796 24070
rect 22744 24006 22796 24012
rect 22756 23662 22784 24006
rect 22940 23730 22968 24754
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 22928 23724 22980 23730
rect 22928 23666 22980 23672
rect 22744 23656 22796 23662
rect 22744 23598 22796 23604
rect 22940 23186 22968 23666
rect 22928 23180 22980 23186
rect 22928 23122 22980 23128
rect 23400 21622 23428 24550
rect 23492 23866 23520 25162
rect 23480 23860 23532 23866
rect 23480 23802 23532 23808
rect 23584 23118 23612 25774
rect 23676 25226 23704 26206
rect 23768 25362 23796 26386
rect 24032 26376 24084 26382
rect 24032 26318 24084 26324
rect 23756 25356 23808 25362
rect 23756 25298 23808 25304
rect 23664 25220 23716 25226
rect 23664 25162 23716 25168
rect 23664 24744 23716 24750
rect 23664 24686 23716 24692
rect 23676 23322 23704 24686
rect 24044 24410 24072 26318
rect 24596 26234 24624 29650
rect 24676 29572 24728 29578
rect 24676 29514 24728 29520
rect 24688 29458 24716 29514
rect 24688 29430 24900 29458
rect 24872 29306 24900 29430
rect 24768 29300 24820 29306
rect 24768 29242 24820 29248
rect 24860 29300 24912 29306
rect 24860 29242 24912 29248
rect 24676 29164 24728 29170
rect 24676 29106 24728 29112
rect 24688 28490 24716 29106
rect 24676 28484 24728 28490
rect 24676 28426 24728 28432
rect 24780 28218 24808 29242
rect 24964 29170 24992 29786
rect 25596 29776 25648 29782
rect 25596 29718 25648 29724
rect 25608 29238 25636 29718
rect 25976 29646 26004 30126
rect 26056 29708 26108 29714
rect 26056 29650 26108 29656
rect 25964 29640 26016 29646
rect 25964 29582 26016 29588
rect 25872 29504 25924 29510
rect 25872 29446 25924 29452
rect 25884 29306 25912 29446
rect 25872 29300 25924 29306
rect 25872 29242 25924 29248
rect 25596 29232 25648 29238
rect 25596 29174 25648 29180
rect 25884 29170 25912 29242
rect 24952 29164 25004 29170
rect 24952 29106 25004 29112
rect 25872 29164 25924 29170
rect 25872 29106 25924 29112
rect 26068 29102 26096 29650
rect 26056 29096 26108 29102
rect 26056 29038 26108 29044
rect 24860 28960 24912 28966
rect 24860 28902 24912 28908
rect 24768 28212 24820 28218
rect 24768 28154 24820 28160
rect 24768 27328 24820 27334
rect 24768 27270 24820 27276
rect 24780 26994 24808 27270
rect 24872 26994 24900 28902
rect 27356 28694 27384 32370
rect 27712 31884 27764 31890
rect 27712 31826 27764 31832
rect 27724 31793 27752 31826
rect 27816 31822 27844 32710
rect 28092 32348 28120 32846
rect 28644 32774 28672 32846
rect 28632 32768 28684 32774
rect 28632 32710 28684 32716
rect 28920 32586 28948 33526
rect 28828 32558 28948 32586
rect 28828 32434 28856 32558
rect 28816 32428 28868 32434
rect 28816 32370 28868 32376
rect 28356 32360 28408 32366
rect 28092 32320 28356 32348
rect 28092 31958 28120 32320
rect 28356 32302 28408 32308
rect 28080 31952 28132 31958
rect 28080 31894 28132 31900
rect 27804 31816 27856 31822
rect 27710 31784 27766 31793
rect 27804 31758 27856 31764
rect 27710 31719 27766 31728
rect 28080 30660 28132 30666
rect 28080 30602 28132 30608
rect 28092 30190 28120 30602
rect 28172 30252 28224 30258
rect 28172 30194 28224 30200
rect 28080 30184 28132 30190
rect 28080 30126 28132 30132
rect 27988 30048 28040 30054
rect 27988 29990 28040 29996
rect 28000 29646 28028 29990
rect 27988 29640 28040 29646
rect 27988 29582 28040 29588
rect 27712 29504 27764 29510
rect 27712 29446 27764 29452
rect 27804 29504 27856 29510
rect 27804 29446 27856 29452
rect 27618 29064 27674 29073
rect 27618 28999 27674 29008
rect 27344 28688 27396 28694
rect 27344 28630 27396 28636
rect 25044 28416 25096 28422
rect 25044 28358 25096 28364
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24860 26988 24912 26994
rect 24860 26930 24912 26936
rect 24860 26852 24912 26858
rect 24860 26794 24912 26800
rect 24872 26382 24900 26794
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 24596 26206 24716 26234
rect 24584 24812 24636 24818
rect 24584 24754 24636 24760
rect 24032 24404 24084 24410
rect 24032 24346 24084 24352
rect 24492 24200 24544 24206
rect 24492 24142 24544 24148
rect 23664 23316 23716 23322
rect 23664 23258 23716 23264
rect 23572 23112 23624 23118
rect 23572 23054 23624 23060
rect 24032 23112 24084 23118
rect 24032 23054 24084 23060
rect 22572 21542 22692 21570
rect 23388 21616 23440 21622
rect 23388 21558 23440 21564
rect 22572 21486 22600 21542
rect 22560 21480 22612 21486
rect 22560 21422 22612 21428
rect 22572 21010 22600 21422
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 22560 21004 22612 21010
rect 22560 20946 22612 20952
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 23400 19718 23428 20402
rect 23572 20256 23624 20262
rect 23572 20198 23624 20204
rect 22928 19712 22980 19718
rect 22928 19654 22980 19660
rect 23388 19712 23440 19718
rect 23388 19654 23440 19660
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22192 18692 22244 18698
rect 22192 18634 22244 18640
rect 22008 17876 22060 17882
rect 22008 17818 22060 17824
rect 21916 17604 21968 17610
rect 21916 17546 21968 17552
rect 21916 17264 21968 17270
rect 21916 17206 21968 17212
rect 21548 17196 21600 17202
rect 21548 17138 21600 17144
rect 21824 17128 21876 17134
rect 21824 17070 21876 17076
rect 21836 16590 21864 17070
rect 21928 16794 21956 17206
rect 22020 17202 22048 17818
rect 22008 17196 22060 17202
rect 22008 17138 22060 17144
rect 22008 17060 22060 17066
rect 22008 17002 22060 17008
rect 22020 16794 22048 17002
rect 21916 16788 21968 16794
rect 21916 16730 21968 16736
rect 22008 16788 22060 16794
rect 22008 16730 22060 16736
rect 21824 16584 21876 16590
rect 21824 16526 21876 16532
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21272 16108 21324 16114
rect 21272 16050 21324 16056
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 20904 15088 20956 15094
rect 20904 15030 20956 15036
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 21088 14884 21140 14890
rect 21088 14826 21140 14832
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 20536 12300 20588 12306
rect 20536 12242 20588 12248
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20456 9722 20576 9738
rect 20456 9716 20588 9722
rect 20456 9710 20536 9716
rect 20536 9658 20588 9664
rect 20444 9648 20496 9654
rect 20444 9590 20496 9596
rect 20456 9178 20484 9590
rect 20916 9586 20944 12174
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 21008 11218 21036 12038
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20548 7818 20576 9522
rect 20812 9444 20864 9450
rect 20812 9386 20864 9392
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 20640 7886 20668 8230
rect 20732 8022 20760 8230
rect 20824 8090 20852 9386
rect 20916 8498 20944 9522
rect 21100 9450 21128 14826
rect 21192 14550 21220 14962
rect 21180 14544 21232 14550
rect 21180 14486 21232 14492
rect 21284 12986 21312 16050
rect 21376 15162 21404 16050
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21928 13530 21956 16730
rect 22008 16652 22060 16658
rect 22008 16594 22060 16600
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 22020 12434 22048 16594
rect 22204 16046 22232 18634
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 22572 18358 22600 18566
rect 22560 18352 22612 18358
rect 22560 18294 22612 18300
rect 22376 17332 22428 17338
rect 22376 17274 22428 17280
rect 22388 16454 22416 17274
rect 22376 16448 22428 16454
rect 22376 16390 22428 16396
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 22204 15434 22232 15982
rect 22192 15428 22244 15434
rect 22192 15370 22244 15376
rect 22284 15088 22336 15094
rect 22284 15030 22336 15036
rect 22296 14006 22324 15030
rect 22388 14482 22416 16390
rect 22376 14476 22428 14482
rect 22376 14418 22428 14424
rect 22940 14414 22968 19654
rect 23204 19372 23256 19378
rect 23204 19314 23256 19320
rect 23216 18970 23244 19314
rect 23204 18964 23256 18970
rect 23204 18906 23256 18912
rect 23480 17808 23532 17814
rect 23480 17750 23532 17756
rect 23492 17678 23520 17750
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23020 17536 23072 17542
rect 23020 17478 23072 17484
rect 23388 17536 23440 17542
rect 23388 17478 23440 17484
rect 23032 17202 23060 17478
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 23400 16998 23428 17478
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 23400 16182 23428 16934
rect 23584 16590 23612 20198
rect 23676 19854 23704 21082
rect 24044 20398 24072 23054
rect 24504 21690 24532 24142
rect 24596 23118 24624 24754
rect 24688 24206 24716 26206
rect 24860 25900 24912 25906
rect 24860 25842 24912 25848
rect 24872 24954 24900 25842
rect 24860 24948 24912 24954
rect 24860 24890 24912 24896
rect 24872 24342 24900 24890
rect 24860 24336 24912 24342
rect 24860 24278 24912 24284
rect 24676 24200 24728 24206
rect 24676 24142 24728 24148
rect 24676 23792 24728 23798
rect 24676 23734 24728 23740
rect 24584 23112 24636 23118
rect 24584 23054 24636 23060
rect 24492 21684 24544 21690
rect 24492 21626 24544 21632
rect 24596 21146 24624 23054
rect 24688 22030 24716 23734
rect 24860 22636 24912 22642
rect 24860 22578 24912 22584
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24676 22024 24728 22030
rect 24676 21966 24728 21972
rect 24584 21140 24636 21146
rect 24584 21082 24636 21088
rect 24780 20942 24808 22374
rect 24872 22166 24900 22578
rect 24860 22160 24912 22166
rect 24860 22102 24912 22108
rect 24768 20936 24820 20942
rect 24768 20878 24820 20884
rect 24032 20392 24084 20398
rect 24032 20334 24084 20340
rect 23756 20324 23808 20330
rect 23756 20266 23808 20272
rect 23664 19848 23716 19854
rect 23664 19790 23716 19796
rect 23768 19334 23796 20266
rect 24860 20052 24912 20058
rect 24860 19994 24912 20000
rect 23848 19780 23900 19786
rect 23848 19722 23900 19728
rect 23860 19514 23888 19722
rect 23848 19508 23900 19514
rect 23848 19450 23900 19456
rect 23676 19306 23796 19334
rect 23676 18766 23704 19306
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 23676 16590 23704 18702
rect 23860 18698 23888 19450
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 24872 17610 24900 19994
rect 25056 17882 25084 28358
rect 27356 27606 27384 28630
rect 27632 28422 27660 28999
rect 27724 28558 27752 29446
rect 27712 28552 27764 28558
rect 27712 28494 27764 28500
rect 27620 28416 27672 28422
rect 27620 28358 27672 28364
rect 27620 28076 27672 28082
rect 27620 28018 27672 28024
rect 26240 27600 26292 27606
rect 26240 27542 26292 27548
rect 27344 27600 27396 27606
rect 27632 27554 27660 28018
rect 27344 27542 27396 27548
rect 25320 27464 25372 27470
rect 25320 27406 25372 27412
rect 25332 27130 25360 27406
rect 25320 27124 25372 27130
rect 25320 27066 25372 27072
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 25148 26858 25176 26930
rect 25136 26852 25188 26858
rect 25136 26794 25188 26800
rect 26252 26382 26280 27542
rect 26240 26376 26292 26382
rect 26240 26318 26292 26324
rect 26608 26376 26660 26382
rect 26608 26318 26660 26324
rect 25780 24880 25832 24886
rect 25780 24822 25832 24828
rect 25228 23724 25280 23730
rect 25228 23666 25280 23672
rect 25240 23322 25268 23666
rect 25228 23316 25280 23322
rect 25228 23258 25280 23264
rect 25792 22642 25820 24822
rect 26424 24268 26476 24274
rect 26424 24210 26476 24216
rect 25964 24200 26016 24206
rect 25964 24142 26016 24148
rect 25976 23254 26004 24142
rect 26148 24132 26200 24138
rect 26148 24074 26200 24080
rect 26056 23316 26108 23322
rect 26056 23258 26108 23264
rect 25964 23248 26016 23254
rect 25964 23190 26016 23196
rect 25872 23044 25924 23050
rect 25872 22986 25924 22992
rect 25884 22778 25912 22986
rect 25872 22772 25924 22778
rect 25872 22714 25924 22720
rect 25780 22636 25832 22642
rect 25780 22578 25832 22584
rect 25964 20460 26016 20466
rect 25964 20402 26016 20408
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 25884 19446 25912 20198
rect 25872 19440 25924 19446
rect 25872 19382 25924 19388
rect 25228 19304 25280 19310
rect 25228 19246 25280 19252
rect 25240 18766 25268 19246
rect 25872 19168 25924 19174
rect 25872 19110 25924 19116
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 25884 18630 25912 19110
rect 25872 18624 25924 18630
rect 25872 18566 25924 18572
rect 25044 17876 25096 17882
rect 25044 17818 25096 17824
rect 25412 17876 25464 17882
rect 25412 17818 25464 17824
rect 24860 17604 24912 17610
rect 24860 17546 24912 17552
rect 25136 17536 25188 17542
rect 25136 17478 25188 17484
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 23952 16794 23980 17138
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 24860 16516 24912 16522
rect 24860 16458 24912 16464
rect 23388 16176 23440 16182
rect 23388 16118 23440 16124
rect 24676 16040 24728 16046
rect 24676 15982 24728 15988
rect 24688 15570 24716 15982
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24136 14550 24164 14962
rect 24124 14544 24176 14550
rect 24124 14486 24176 14492
rect 23204 14476 23256 14482
rect 23204 14418 23256 14424
rect 22928 14408 22980 14414
rect 22928 14350 22980 14356
rect 22284 14000 22336 14006
rect 22284 13942 22336 13948
rect 23216 13938 23244 14418
rect 23296 14000 23348 14006
rect 23296 13942 23348 13948
rect 23204 13932 23256 13938
rect 23204 13874 23256 13880
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 21928 12406 22048 12434
rect 21364 12368 21416 12374
rect 21364 12310 21416 12316
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 21192 10130 21220 12174
rect 21376 12102 21404 12310
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21376 11354 21404 12038
rect 21468 11762 21496 12174
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21180 10124 21232 10130
rect 21180 10066 21232 10072
rect 21192 9926 21220 10066
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 21088 9444 21140 9450
rect 21088 9386 21140 9392
rect 21928 8974 21956 12406
rect 22296 12170 22324 13806
rect 23308 12442 23336 13942
rect 23388 13524 23440 13530
rect 23388 13466 23440 13472
rect 23400 12714 23428 13466
rect 23572 12776 23624 12782
rect 23572 12718 23624 12724
rect 23388 12708 23440 12714
rect 23388 12650 23440 12656
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23296 12436 23348 12442
rect 23296 12378 23348 12384
rect 22284 12164 22336 12170
rect 22284 12106 22336 12112
rect 23492 11694 23520 12582
rect 23584 11898 23612 12718
rect 23848 12436 23900 12442
rect 23848 12378 23900 12384
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 23860 11830 23888 12378
rect 24136 11898 24164 14486
rect 24584 13728 24636 13734
rect 24584 13670 24636 13676
rect 24596 13394 24624 13670
rect 24584 13388 24636 13394
rect 24584 13330 24636 13336
rect 24596 12306 24624 13330
rect 24688 12986 24716 15506
rect 24872 15502 24900 16458
rect 25044 15904 25096 15910
rect 25044 15846 25096 15852
rect 25056 15502 25084 15846
rect 25148 15502 25176 17478
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 25240 16522 25268 16934
rect 25228 16516 25280 16522
rect 25228 16458 25280 16464
rect 24860 15496 24912 15502
rect 24860 15438 24912 15444
rect 25044 15496 25096 15502
rect 25044 15438 25096 15444
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 25148 14822 25176 15438
rect 25320 15088 25372 15094
rect 25320 15030 25372 15036
rect 25136 14816 25188 14822
rect 25136 14758 25188 14764
rect 25332 14482 25360 15030
rect 25320 14476 25372 14482
rect 25320 14418 25372 14424
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24308 12164 24360 12170
rect 24308 12106 24360 12112
rect 24320 11898 24348 12106
rect 24872 12102 24900 13874
rect 25332 12442 25360 14418
rect 25320 12436 25372 12442
rect 25320 12378 25372 12384
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24124 11892 24176 11898
rect 24124 11834 24176 11840
rect 24308 11892 24360 11898
rect 24308 11834 24360 11840
rect 23848 11824 23900 11830
rect 23848 11766 23900 11772
rect 22008 11688 22060 11694
rect 22008 11630 22060 11636
rect 23480 11688 23532 11694
rect 23480 11630 23532 11636
rect 22020 11150 22048 11630
rect 23388 11620 23440 11626
rect 23388 11562 23440 11568
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22020 10266 22048 11086
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 23400 8906 23428 11562
rect 23572 11552 23624 11558
rect 23572 11494 23624 11500
rect 23584 9178 23612 11494
rect 24872 10062 24900 12038
rect 25228 11688 25280 11694
rect 25228 11630 25280 11636
rect 25240 10062 25268 11630
rect 25332 10062 25360 12378
rect 25424 11558 25452 17818
rect 25780 16448 25832 16454
rect 25780 16390 25832 16396
rect 25792 16182 25820 16390
rect 25780 16176 25832 16182
rect 25780 16118 25832 16124
rect 25884 15994 25912 18566
rect 25792 15966 25912 15994
rect 25792 12850 25820 15966
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 25780 12844 25832 12850
rect 25780 12786 25832 12792
rect 25884 11762 25912 15302
rect 25976 13870 26004 20402
rect 26068 19854 26096 23258
rect 26160 22982 26188 24074
rect 26436 23730 26464 24210
rect 26424 23724 26476 23730
rect 26424 23666 26476 23672
rect 26240 23656 26292 23662
rect 26240 23598 26292 23604
rect 26148 22976 26200 22982
rect 26148 22918 26200 22924
rect 26056 19848 26108 19854
rect 26056 19790 26108 19796
rect 26056 18760 26108 18766
rect 26056 18702 26108 18708
rect 26068 18426 26096 18702
rect 26056 18420 26108 18426
rect 26056 18362 26108 18368
rect 26160 16590 26188 22918
rect 26252 22778 26280 23598
rect 26516 23044 26568 23050
rect 26516 22986 26568 22992
rect 26240 22772 26292 22778
rect 26240 22714 26292 22720
rect 26332 22636 26384 22642
rect 26332 22578 26384 22584
rect 26240 22024 26292 22030
rect 26240 21966 26292 21972
rect 26252 18970 26280 21966
rect 26344 20466 26372 22578
rect 26528 22234 26556 22986
rect 26516 22228 26568 22234
rect 26516 22170 26568 22176
rect 26620 22098 26648 26318
rect 27356 24274 27384 27542
rect 27448 27526 27660 27554
rect 27448 26858 27476 27526
rect 27724 27470 27752 28494
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 27620 27396 27672 27402
rect 27620 27338 27672 27344
rect 27632 26994 27660 27338
rect 27620 26988 27672 26994
rect 27620 26930 27672 26936
rect 27436 26852 27488 26858
rect 27436 26794 27488 26800
rect 27344 24268 27396 24274
rect 27344 24210 27396 24216
rect 27448 23730 27476 26794
rect 27528 26308 27580 26314
rect 27528 26250 27580 26256
rect 27436 23724 27488 23730
rect 27436 23666 27488 23672
rect 26608 22092 26660 22098
rect 26608 22034 26660 22040
rect 26608 20528 26660 20534
rect 26608 20470 26660 20476
rect 26332 20460 26384 20466
rect 26332 20402 26384 20408
rect 26620 19514 26648 20470
rect 26884 19780 26936 19786
rect 26884 19722 26936 19728
rect 26608 19508 26660 19514
rect 26608 19450 26660 19456
rect 26896 19446 26924 19722
rect 26884 19440 26936 19446
rect 26884 19382 26936 19388
rect 26896 18970 26924 19382
rect 27160 19168 27212 19174
rect 27160 19110 27212 19116
rect 26240 18964 26292 18970
rect 26240 18906 26292 18912
rect 26884 18964 26936 18970
rect 26884 18906 26936 18912
rect 27172 18698 27200 19110
rect 27160 18692 27212 18698
rect 27160 18634 27212 18640
rect 26240 18284 26292 18290
rect 26240 18226 26292 18232
rect 26252 17542 26280 18226
rect 27448 18222 27476 23666
rect 27540 22778 27568 26250
rect 27620 25220 27672 25226
rect 27620 25162 27672 25168
rect 27632 24410 27660 25162
rect 27816 24834 27844 29446
rect 28092 29306 28120 30126
rect 28080 29300 28132 29306
rect 28080 29242 28132 29248
rect 28184 28082 28212 30194
rect 28356 30116 28408 30122
rect 28356 30058 28408 30064
rect 28368 29782 28396 30058
rect 28356 29776 28408 29782
rect 28356 29718 28408 29724
rect 28264 28688 28316 28694
rect 28264 28630 28316 28636
rect 28172 28076 28224 28082
rect 28172 28018 28224 28024
rect 28172 27872 28224 27878
rect 28172 27814 28224 27820
rect 28184 26994 28212 27814
rect 28276 27470 28304 28630
rect 28368 28422 28396 29718
rect 28724 29572 28776 29578
rect 28724 29514 28776 29520
rect 28736 29170 28764 29514
rect 28724 29164 28776 29170
rect 28724 29106 28776 29112
rect 28724 28484 28776 28490
rect 28724 28426 28776 28432
rect 28356 28416 28408 28422
rect 28356 28358 28408 28364
rect 28264 27464 28316 27470
rect 28264 27406 28316 27412
rect 28368 27402 28396 28358
rect 28448 28076 28500 28082
rect 28448 28018 28500 28024
rect 28460 27538 28488 28018
rect 28448 27532 28500 27538
rect 28448 27474 28500 27480
rect 28736 27470 28764 28426
rect 28816 28416 28868 28422
rect 28816 28358 28868 28364
rect 28828 28082 28856 28358
rect 28816 28076 28868 28082
rect 28816 28018 28868 28024
rect 28724 27464 28776 27470
rect 28724 27406 28776 27412
rect 28356 27396 28408 27402
rect 28356 27338 28408 27344
rect 28724 27124 28776 27130
rect 28724 27066 28776 27072
rect 27896 26988 27948 26994
rect 27896 26930 27948 26936
rect 27988 26988 28040 26994
rect 27988 26930 28040 26936
rect 28172 26988 28224 26994
rect 28172 26930 28224 26936
rect 28632 26988 28684 26994
rect 28632 26930 28684 26936
rect 27908 26518 27936 26930
rect 28000 26518 28028 26930
rect 27896 26512 27948 26518
rect 27896 26454 27948 26460
rect 27988 26512 28040 26518
rect 27988 26454 28040 26460
rect 27724 24806 27844 24834
rect 27620 24404 27672 24410
rect 27620 24346 27672 24352
rect 27620 24268 27672 24274
rect 27620 24210 27672 24216
rect 27528 22772 27580 22778
rect 27528 22714 27580 22720
rect 27632 22642 27660 24210
rect 27620 22636 27672 22642
rect 27620 22578 27672 22584
rect 27620 22432 27672 22438
rect 27620 22374 27672 22380
rect 27632 22030 27660 22374
rect 27724 22098 27752 24806
rect 27804 24744 27856 24750
rect 27804 24686 27856 24692
rect 27816 24206 27844 24686
rect 27804 24200 27856 24206
rect 27804 24142 27856 24148
rect 27908 22642 27936 26454
rect 28080 26444 28132 26450
rect 28080 26386 28132 26392
rect 28092 24274 28120 26386
rect 28080 24268 28132 24274
rect 28080 24210 28132 24216
rect 28170 22672 28226 22681
rect 27896 22636 27948 22642
rect 28170 22607 28172 22616
rect 27896 22578 27948 22584
rect 28224 22607 28226 22616
rect 28172 22578 28224 22584
rect 27988 22500 28040 22506
rect 27988 22442 28040 22448
rect 27804 22228 27856 22234
rect 27804 22170 27856 22176
rect 27712 22092 27764 22098
rect 27712 22034 27764 22040
rect 27620 22024 27672 22030
rect 27620 21966 27672 21972
rect 27620 20460 27672 20466
rect 27620 20402 27672 20408
rect 27528 19712 27580 19718
rect 27528 19654 27580 19660
rect 27540 18902 27568 19654
rect 27632 19378 27660 20402
rect 27620 19372 27672 19378
rect 27620 19314 27672 19320
rect 27528 18896 27580 18902
rect 27528 18838 27580 18844
rect 27436 18216 27488 18222
rect 27436 18158 27488 18164
rect 27816 17882 27844 22170
rect 28000 21944 28028 22442
rect 28080 21956 28132 21962
rect 28000 21916 28080 21944
rect 28000 21554 28028 21916
rect 28080 21898 28132 21904
rect 27988 21548 28040 21554
rect 27988 21490 28040 21496
rect 28172 21548 28224 21554
rect 28172 21490 28224 21496
rect 28184 20058 28212 21490
rect 28644 20058 28672 26930
rect 28736 25158 28764 27066
rect 28724 25152 28776 25158
rect 28724 25094 28776 25100
rect 28736 24138 28764 25094
rect 28920 24614 28948 32558
rect 29472 31754 29500 35634
rect 29644 35556 29696 35562
rect 29644 35498 29696 35504
rect 29552 35216 29604 35222
rect 29552 35158 29604 35164
rect 29564 34610 29592 35158
rect 29552 34604 29604 34610
rect 29552 34546 29604 34552
rect 29564 33522 29592 34546
rect 29552 33516 29604 33522
rect 29552 33458 29604 33464
rect 29656 32434 29684 35498
rect 30116 35154 30144 36518
rect 31036 36378 31064 36722
rect 31208 36712 31260 36718
rect 31208 36654 31260 36660
rect 30380 36372 30432 36378
rect 30380 36314 30432 36320
rect 31024 36372 31076 36378
rect 31024 36314 31076 36320
rect 30392 36174 30420 36314
rect 30380 36168 30432 36174
rect 30380 36110 30432 36116
rect 30288 36032 30340 36038
rect 30288 35974 30340 35980
rect 30300 35766 30328 35974
rect 30288 35760 30340 35766
rect 30288 35702 30340 35708
rect 30392 35698 30420 36110
rect 30472 36100 30524 36106
rect 30472 36042 30524 36048
rect 30484 35834 30512 36042
rect 30840 36032 30892 36038
rect 30840 35974 30892 35980
rect 30472 35828 30524 35834
rect 30472 35770 30524 35776
rect 30484 35698 30512 35770
rect 30380 35692 30432 35698
rect 30380 35634 30432 35640
rect 30472 35692 30524 35698
rect 30472 35634 30524 35640
rect 30012 35148 30064 35154
rect 30012 35090 30064 35096
rect 30104 35148 30156 35154
rect 30104 35090 30156 35096
rect 30024 34950 30052 35090
rect 30012 34944 30064 34950
rect 30012 34886 30064 34892
rect 30392 34746 30420 35634
rect 30380 34740 30432 34746
rect 30380 34682 30432 34688
rect 29736 33516 29788 33522
rect 29736 33458 29788 33464
rect 29748 33046 29776 33458
rect 29736 33040 29788 33046
rect 29736 32982 29788 32988
rect 29644 32428 29696 32434
rect 29644 32370 29696 32376
rect 29472 31726 29592 31754
rect 29184 30592 29236 30598
rect 29184 30534 29236 30540
rect 29276 30592 29328 30598
rect 29276 30534 29328 30540
rect 29196 30326 29224 30534
rect 29184 30320 29236 30326
rect 29184 30262 29236 30268
rect 29196 29714 29224 30262
rect 29288 30258 29316 30534
rect 29276 30252 29328 30258
rect 29276 30194 29328 30200
rect 29288 29850 29316 30194
rect 29276 29844 29328 29850
rect 29276 29786 29328 29792
rect 29184 29708 29236 29714
rect 29184 29650 29236 29656
rect 29564 29510 29592 31726
rect 29656 30938 29684 32370
rect 30484 31346 30512 35634
rect 30852 35630 30880 35974
rect 30840 35624 30892 35630
rect 30840 35566 30892 35572
rect 30852 35290 30880 35566
rect 31220 35494 31248 36654
rect 33232 36236 33284 36242
rect 33232 36178 33284 36184
rect 31392 36168 31444 36174
rect 31392 36110 31444 36116
rect 31404 35766 31432 36110
rect 31392 35760 31444 35766
rect 31392 35702 31444 35708
rect 32956 35692 33008 35698
rect 32956 35634 33008 35640
rect 32128 35624 32180 35630
rect 32128 35566 32180 35572
rect 31208 35488 31260 35494
rect 31208 35430 31260 35436
rect 30840 35284 30892 35290
rect 30840 35226 30892 35232
rect 32140 35086 32168 35566
rect 32968 35154 32996 35634
rect 33140 35488 33192 35494
rect 33140 35430 33192 35436
rect 32312 35148 32364 35154
rect 32312 35090 32364 35096
rect 32956 35148 33008 35154
rect 32956 35090 33008 35096
rect 32128 35080 32180 35086
rect 32128 35022 32180 35028
rect 30840 35012 30892 35018
rect 30840 34954 30892 34960
rect 30852 34610 30880 34954
rect 30840 34604 30892 34610
rect 30840 34546 30892 34552
rect 32140 34542 32168 35022
rect 32324 34610 32352 35090
rect 33048 35012 33100 35018
rect 33048 34954 33100 34960
rect 32956 34944 33008 34950
rect 32956 34886 33008 34892
rect 32404 34672 32456 34678
rect 32404 34614 32456 34620
rect 32312 34604 32364 34610
rect 32312 34546 32364 34552
rect 32128 34536 32180 34542
rect 32128 34478 32180 34484
rect 31668 33992 31720 33998
rect 31668 33934 31720 33940
rect 31680 33454 31708 33934
rect 32324 33658 32352 34546
rect 32416 34406 32444 34614
rect 32772 34536 32824 34542
rect 32772 34478 32824 34484
rect 32404 34400 32456 34406
rect 32404 34342 32456 34348
rect 32312 33652 32364 33658
rect 32312 33594 32364 33600
rect 32416 33590 32444 34342
rect 32784 34202 32812 34478
rect 32772 34196 32824 34202
rect 32772 34138 32824 34144
rect 32496 33924 32548 33930
rect 32496 33866 32548 33872
rect 32404 33584 32456 33590
rect 32404 33526 32456 33532
rect 32508 33522 32536 33866
rect 32496 33516 32548 33522
rect 32496 33458 32548 33464
rect 31668 33448 31720 33454
rect 31668 33390 31720 33396
rect 31680 32298 31708 33390
rect 31668 32292 31720 32298
rect 31668 32234 31720 32240
rect 31024 31408 31076 31414
rect 31024 31350 31076 31356
rect 30472 31340 30524 31346
rect 30472 31282 30524 31288
rect 30656 31340 30708 31346
rect 30656 31282 30708 31288
rect 29828 31136 29880 31142
rect 29828 31078 29880 31084
rect 29644 30932 29696 30938
rect 29644 30874 29696 30880
rect 29736 30796 29788 30802
rect 29736 30738 29788 30744
rect 29748 30054 29776 30738
rect 29840 30258 29868 31078
rect 29920 30864 29972 30870
rect 29920 30806 29972 30812
rect 29932 30598 29960 30806
rect 30484 30802 30512 31282
rect 30668 30818 30696 31282
rect 30472 30796 30524 30802
rect 30472 30738 30524 30744
rect 30576 30790 30696 30818
rect 30576 30734 30604 30790
rect 31036 30734 31064 31350
rect 30196 30728 30248 30734
rect 30196 30670 30248 30676
rect 30564 30728 30616 30734
rect 30564 30670 30616 30676
rect 31024 30728 31076 30734
rect 31024 30670 31076 30676
rect 29920 30592 29972 30598
rect 29920 30534 29972 30540
rect 29932 30326 29960 30534
rect 29920 30320 29972 30326
rect 29920 30262 29972 30268
rect 29828 30252 29880 30258
rect 29828 30194 29880 30200
rect 29736 30048 29788 30054
rect 29736 29990 29788 29996
rect 29748 29646 29776 29990
rect 30208 29850 30236 30670
rect 30576 30258 30604 30670
rect 31036 30326 31064 30670
rect 31024 30320 31076 30326
rect 31024 30262 31076 30268
rect 30564 30252 30616 30258
rect 30564 30194 30616 30200
rect 32220 30252 32272 30258
rect 32220 30194 32272 30200
rect 30576 29850 30604 30194
rect 30196 29844 30248 29850
rect 30196 29786 30248 29792
rect 30564 29844 30616 29850
rect 30564 29786 30616 29792
rect 32232 29646 32260 30194
rect 32404 30184 32456 30190
rect 32404 30126 32456 30132
rect 32416 29646 32444 30126
rect 29736 29640 29788 29646
rect 29736 29582 29788 29588
rect 32220 29640 32272 29646
rect 32220 29582 32272 29588
rect 32404 29640 32456 29646
rect 32404 29582 32456 29588
rect 31668 29572 31720 29578
rect 31668 29514 31720 29520
rect 29552 29504 29604 29510
rect 29552 29446 29604 29452
rect 29828 29504 29880 29510
rect 29828 29446 29880 29452
rect 29184 29096 29236 29102
rect 29184 29038 29236 29044
rect 29276 29096 29328 29102
rect 29276 29038 29328 29044
rect 29092 28960 29144 28966
rect 29092 28902 29144 28908
rect 29104 28218 29132 28902
rect 29196 28694 29224 29038
rect 29288 28966 29316 29038
rect 29276 28960 29328 28966
rect 29276 28902 29328 28908
rect 29736 28960 29788 28966
rect 29736 28902 29788 28908
rect 29184 28688 29236 28694
rect 29184 28630 29236 28636
rect 29092 28212 29144 28218
rect 29092 28154 29144 28160
rect 29288 28082 29316 28902
rect 29748 28490 29776 28902
rect 29736 28484 29788 28490
rect 29736 28426 29788 28432
rect 29552 28416 29604 28422
rect 29552 28358 29604 28364
rect 29564 28082 29592 28358
rect 29276 28076 29328 28082
rect 29276 28018 29328 28024
rect 29552 28076 29604 28082
rect 29552 28018 29604 28024
rect 29564 27674 29592 28018
rect 29552 27668 29604 27674
rect 29552 27610 29604 27616
rect 29736 24812 29788 24818
rect 29736 24754 29788 24760
rect 28908 24608 28960 24614
rect 28908 24550 28960 24556
rect 28724 24132 28776 24138
rect 28724 24074 28776 24080
rect 29748 23866 29776 24754
rect 29840 24342 29868 29446
rect 31116 29028 31168 29034
rect 31116 28970 31168 28976
rect 29920 28756 29972 28762
rect 29920 28698 29972 28704
rect 29932 28218 29960 28698
rect 29920 28212 29972 28218
rect 29920 28154 29972 28160
rect 31128 28082 31156 28970
rect 31680 28098 31708 29514
rect 31220 28082 31892 28098
rect 31116 28076 31168 28082
rect 31116 28018 31168 28024
rect 31220 28076 31904 28082
rect 31220 28070 31852 28076
rect 31220 25906 31248 28070
rect 31852 28018 31904 28024
rect 31760 28008 31812 28014
rect 31680 27956 31760 27962
rect 31680 27950 31812 27956
rect 31484 27940 31536 27946
rect 31484 27882 31536 27888
rect 31680 27934 31800 27950
rect 31496 27538 31524 27882
rect 31484 27532 31536 27538
rect 31484 27474 31536 27480
rect 31680 27334 31708 27934
rect 32036 27872 32088 27878
rect 32036 27814 32088 27820
rect 32312 27872 32364 27878
rect 32312 27814 32364 27820
rect 32048 27470 32076 27814
rect 32036 27464 32088 27470
rect 32036 27406 32088 27412
rect 32324 27402 32352 27814
rect 32312 27396 32364 27402
rect 32312 27338 32364 27344
rect 31392 27328 31444 27334
rect 31392 27270 31444 27276
rect 31668 27328 31720 27334
rect 31668 27270 31720 27276
rect 31404 26994 31432 27270
rect 32508 27062 32536 33458
rect 32968 32366 32996 34886
rect 33060 34678 33088 34954
rect 33048 34672 33100 34678
rect 33048 34614 33100 34620
rect 33152 34610 33180 35430
rect 33244 34746 33272 36178
rect 34532 36174 34560 37062
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 37200 36174 37228 37266
rect 38212 37262 38240 39200
rect 38200 37256 38252 37262
rect 38200 37198 38252 37204
rect 33416 36168 33468 36174
rect 33416 36110 33468 36116
rect 34520 36168 34572 36174
rect 34520 36110 34572 36116
rect 37188 36168 37240 36174
rect 37188 36110 37240 36116
rect 33428 35154 33456 36110
rect 34060 36032 34112 36038
rect 34060 35974 34112 35980
rect 34244 36032 34296 36038
rect 34244 35974 34296 35980
rect 33600 35556 33652 35562
rect 33600 35498 33652 35504
rect 33416 35148 33468 35154
rect 33416 35090 33468 35096
rect 33232 34740 33284 34746
rect 33232 34682 33284 34688
rect 33140 34604 33192 34610
rect 33140 34546 33192 34552
rect 32956 32360 33008 32366
rect 32956 32302 33008 32308
rect 33232 31884 33284 31890
rect 33232 31826 33284 31832
rect 32956 30252 33008 30258
rect 32956 30194 33008 30200
rect 33140 30252 33192 30258
rect 33140 30194 33192 30200
rect 32968 29782 32996 30194
rect 32956 29776 33008 29782
rect 32956 29718 33008 29724
rect 33152 29646 33180 30194
rect 33244 29850 33272 31826
rect 33428 30666 33456 35090
rect 33612 35018 33640 35498
rect 34072 35086 34100 35974
rect 34060 35080 34112 35086
rect 34060 35022 34112 35028
rect 33600 35012 33652 35018
rect 33600 34954 33652 34960
rect 33508 32224 33560 32230
rect 33508 32166 33560 32172
rect 33520 31822 33548 32166
rect 33508 31816 33560 31822
rect 33508 31758 33560 31764
rect 33416 30660 33468 30666
rect 33416 30602 33468 30608
rect 33324 30116 33376 30122
rect 33324 30058 33376 30064
rect 33232 29844 33284 29850
rect 33232 29786 33284 29792
rect 33140 29640 33192 29646
rect 33140 29582 33192 29588
rect 33232 29640 33284 29646
rect 33232 29582 33284 29588
rect 33048 28552 33100 28558
rect 33048 28494 33100 28500
rect 33060 28150 33088 28494
rect 33048 28144 33100 28150
rect 32968 28092 33048 28098
rect 32968 28086 33100 28092
rect 32968 28070 33088 28086
rect 32680 27600 32732 27606
rect 32680 27542 32732 27548
rect 32692 27418 32720 27542
rect 32968 27470 32996 28070
rect 33152 28014 33180 29582
rect 33244 28966 33272 29582
rect 33336 29578 33364 30058
rect 33324 29572 33376 29578
rect 33324 29514 33376 29520
rect 33336 29034 33364 29514
rect 33508 29504 33560 29510
rect 33508 29446 33560 29452
rect 33324 29028 33376 29034
rect 33324 28970 33376 28976
rect 33232 28960 33284 28966
rect 33232 28902 33284 28908
rect 33336 28490 33364 28970
rect 33520 28694 33548 29446
rect 33508 28688 33560 28694
rect 33508 28630 33560 28636
rect 33416 28552 33468 28558
rect 33416 28494 33468 28500
rect 33324 28484 33376 28490
rect 33324 28426 33376 28432
rect 33428 28082 33456 28494
rect 33416 28076 33468 28082
rect 33416 28018 33468 28024
rect 33140 28008 33192 28014
rect 33140 27950 33192 27956
rect 33048 27940 33100 27946
rect 33048 27882 33100 27888
rect 33060 27470 33088 27882
rect 33428 27674 33456 28018
rect 33416 27668 33468 27674
rect 33416 27610 33468 27616
rect 33612 27554 33640 34954
rect 33876 34468 33928 34474
rect 33876 34410 33928 34416
rect 33784 31816 33836 31822
rect 33784 31758 33836 31764
rect 33796 31278 33824 31758
rect 33784 31272 33836 31278
rect 33784 31214 33836 31220
rect 33692 30660 33744 30666
rect 33692 30602 33744 30608
rect 33704 30326 33732 30602
rect 33692 30320 33744 30326
rect 33692 30262 33744 30268
rect 33704 29646 33732 30262
rect 33692 29640 33744 29646
rect 33692 29582 33744 29588
rect 33704 28082 33732 29582
rect 33692 28076 33744 28082
rect 33692 28018 33744 28024
rect 33796 28014 33824 31214
rect 33888 30734 33916 34410
rect 34060 31680 34112 31686
rect 34060 31622 34112 31628
rect 34152 31680 34204 31686
rect 34152 31622 34204 31628
rect 34072 31346 34100 31622
rect 34164 31346 34192 31622
rect 34060 31340 34112 31346
rect 34060 31282 34112 31288
rect 34152 31340 34204 31346
rect 34152 31282 34204 31288
rect 34164 30938 34192 31282
rect 34152 30932 34204 30938
rect 34152 30874 34204 30880
rect 33876 30728 33928 30734
rect 33876 30670 33928 30676
rect 33888 30394 33916 30670
rect 33876 30388 33928 30394
rect 33876 30330 33928 30336
rect 34256 30054 34284 35974
rect 34428 35692 34480 35698
rect 34428 35634 34480 35640
rect 34440 32570 34468 35634
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35992 34944 36044 34950
rect 35992 34886 36044 34892
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34428 32564 34480 32570
rect 34428 32506 34480 32512
rect 34520 32496 34572 32502
rect 34520 32438 34572 32444
rect 34532 31414 34560 32438
rect 36004 32434 36032 34886
rect 35992 32428 36044 32434
rect 35992 32370 36044 32376
rect 35348 32360 35400 32366
rect 35348 32302 35400 32308
rect 34612 32224 34664 32230
rect 34612 32166 34664 32172
rect 34624 31822 34652 32166
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34796 31884 34848 31890
rect 34796 31826 34848 31832
rect 34612 31816 34664 31822
rect 34612 31758 34664 31764
rect 34612 31680 34664 31686
rect 34612 31622 34664 31628
rect 34520 31408 34572 31414
rect 34520 31350 34572 31356
rect 34428 31204 34480 31210
rect 34428 31146 34480 31152
rect 34440 30258 34468 31146
rect 34624 30802 34652 31622
rect 34808 30802 34836 31826
rect 35360 31686 35388 32302
rect 35440 31884 35492 31890
rect 35440 31826 35492 31832
rect 35348 31680 35400 31686
rect 35348 31622 35400 31628
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35452 30870 35480 31826
rect 35440 30864 35492 30870
rect 35440 30806 35492 30812
rect 34612 30796 34664 30802
rect 34612 30738 34664 30744
rect 34796 30796 34848 30802
rect 34796 30738 34848 30744
rect 34428 30252 34480 30258
rect 34428 30194 34480 30200
rect 34244 30048 34296 30054
rect 34244 29990 34296 29996
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34336 28620 34388 28626
rect 34336 28562 34388 28568
rect 34348 28082 34376 28562
rect 34336 28076 34388 28082
rect 34336 28018 34388 28024
rect 33784 28008 33836 28014
rect 33784 27950 33836 27956
rect 33428 27526 33640 27554
rect 32956 27464 33008 27470
rect 32692 27402 32812 27418
rect 32956 27406 33008 27412
rect 33048 27464 33100 27470
rect 33048 27406 33100 27412
rect 32692 27396 32824 27402
rect 32692 27390 32772 27396
rect 32496 27056 32548 27062
rect 32496 26998 32548 27004
rect 31392 26988 31444 26994
rect 31392 26930 31444 26936
rect 31852 26988 31904 26994
rect 31852 26930 31904 26936
rect 32588 26988 32640 26994
rect 32588 26930 32640 26936
rect 31864 26314 31892 26930
rect 32600 26518 32628 26930
rect 32588 26512 32640 26518
rect 32588 26454 32640 26460
rect 32692 26314 32720 27390
rect 32772 27338 32824 27344
rect 32968 27130 32996 27406
rect 33048 27328 33100 27334
rect 33048 27270 33100 27276
rect 32956 27124 33008 27130
rect 32956 27066 33008 27072
rect 32864 26920 32916 26926
rect 32864 26862 32916 26868
rect 32876 26382 32904 26862
rect 33060 26450 33088 27270
rect 33428 26926 33456 27526
rect 33416 26920 33468 26926
rect 33416 26862 33468 26868
rect 33428 26518 33456 26862
rect 34348 26586 34376 28018
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34336 26580 34388 26586
rect 34336 26522 34388 26528
rect 33416 26512 33468 26518
rect 33416 26454 33468 26460
rect 33048 26444 33100 26450
rect 33048 26386 33100 26392
rect 32864 26376 32916 26382
rect 32864 26318 32916 26324
rect 31852 26308 31904 26314
rect 31852 26250 31904 26256
rect 32680 26308 32732 26314
rect 32680 26250 32732 26256
rect 31300 26240 31352 26246
rect 31300 26182 31352 26188
rect 30932 25900 30984 25906
rect 30932 25842 30984 25848
rect 31024 25900 31076 25906
rect 31024 25842 31076 25848
rect 31208 25900 31260 25906
rect 31208 25842 31260 25848
rect 29920 25696 29972 25702
rect 29920 25638 29972 25644
rect 30840 25696 30892 25702
rect 30840 25638 30892 25644
rect 29932 25294 29960 25638
rect 29920 25288 29972 25294
rect 29920 25230 29972 25236
rect 29828 24336 29880 24342
rect 29828 24278 29880 24284
rect 30852 24138 30880 25638
rect 30944 24682 30972 25842
rect 30932 24676 30984 24682
rect 30932 24618 30984 24624
rect 30840 24132 30892 24138
rect 30840 24074 30892 24080
rect 29736 23860 29788 23866
rect 29736 23802 29788 23808
rect 30944 23118 30972 24618
rect 30932 23112 30984 23118
rect 30932 23054 30984 23060
rect 31036 22710 31064 25842
rect 31220 24410 31248 25842
rect 31312 25294 31340 26182
rect 31864 25498 31892 26250
rect 32588 26240 32640 26246
rect 32588 26182 32640 26188
rect 32312 25900 32364 25906
rect 32312 25842 32364 25848
rect 31852 25492 31904 25498
rect 31852 25434 31904 25440
rect 31300 25288 31352 25294
rect 31300 25230 31352 25236
rect 32324 24886 32352 25842
rect 32600 25158 32628 26182
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 32588 25152 32640 25158
rect 32588 25094 32640 25100
rect 32312 24880 32364 24886
rect 32312 24822 32364 24828
rect 31208 24404 31260 24410
rect 31208 24346 31260 24352
rect 31760 24064 31812 24070
rect 31760 24006 31812 24012
rect 31024 22704 31076 22710
rect 31024 22646 31076 22652
rect 29920 22636 29972 22642
rect 29920 22578 29972 22584
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 29552 22568 29604 22574
rect 29552 22510 29604 22516
rect 29564 22098 29592 22510
rect 29932 22234 29960 22578
rect 30748 22500 30800 22506
rect 30748 22442 30800 22448
rect 29920 22228 29972 22234
rect 29920 22170 29972 22176
rect 29552 22092 29604 22098
rect 29552 22034 29604 22040
rect 30760 22030 30788 22442
rect 30944 22030 30972 22578
rect 30748 22024 30800 22030
rect 30748 21966 30800 21972
rect 30932 22024 30984 22030
rect 30932 21966 30984 21972
rect 28908 21956 28960 21962
rect 28908 21898 28960 21904
rect 28920 21010 28948 21898
rect 29736 21480 29788 21486
rect 29736 21422 29788 21428
rect 28908 21004 28960 21010
rect 28908 20946 28960 20952
rect 29000 20800 29052 20806
rect 29000 20742 29052 20748
rect 28172 20052 28224 20058
rect 28172 19994 28224 20000
rect 28356 20052 28408 20058
rect 28356 19994 28408 20000
rect 28632 20052 28684 20058
rect 28632 19994 28684 20000
rect 28264 19848 28316 19854
rect 28264 19790 28316 19796
rect 28276 18970 28304 19790
rect 28264 18964 28316 18970
rect 28264 18906 28316 18912
rect 27804 17876 27856 17882
rect 27804 17818 27856 17824
rect 27252 17604 27304 17610
rect 27252 17546 27304 17552
rect 26240 17536 26292 17542
rect 26240 17478 26292 17484
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 26056 16516 26108 16522
rect 26056 16458 26108 16464
rect 26068 15094 26096 16458
rect 26148 16448 26200 16454
rect 26148 16390 26200 16396
rect 26160 15910 26188 16390
rect 26148 15904 26200 15910
rect 26148 15846 26200 15852
rect 26148 15428 26200 15434
rect 26148 15370 26200 15376
rect 26160 15162 26188 15370
rect 26148 15156 26200 15162
rect 26148 15098 26200 15104
rect 26056 15088 26108 15094
rect 26056 15030 26108 15036
rect 25964 13864 26016 13870
rect 25964 13806 26016 13812
rect 26252 12918 26280 17478
rect 26332 16652 26384 16658
rect 26332 16594 26384 16600
rect 26344 15026 26372 16594
rect 26516 15360 26568 15366
rect 26516 15302 26568 15308
rect 26528 15162 26556 15302
rect 26516 15156 26568 15162
rect 26516 15098 26568 15104
rect 26332 15020 26384 15026
rect 26332 14962 26384 14968
rect 26528 14906 26556 15098
rect 26344 14878 26556 14906
rect 26344 14414 26372 14878
rect 26424 14816 26476 14822
rect 26424 14758 26476 14764
rect 26332 14408 26384 14414
rect 26332 14350 26384 14356
rect 26436 14362 26464 14758
rect 26436 14346 26556 14362
rect 26436 14340 26568 14346
rect 26436 14334 26516 14340
rect 26516 14282 26568 14288
rect 26792 14340 26844 14346
rect 26792 14282 26844 14288
rect 26700 14272 26752 14278
rect 26700 14214 26752 14220
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 26332 13184 26384 13190
rect 26332 13126 26384 13132
rect 26344 12918 26372 13126
rect 26240 12912 26292 12918
rect 26240 12854 26292 12860
rect 26332 12912 26384 12918
rect 26332 12854 26384 12860
rect 26148 12776 26200 12782
rect 26148 12718 26200 12724
rect 26160 12458 26188 12718
rect 26068 12442 26188 12458
rect 26056 12436 26188 12442
rect 26108 12430 26188 12436
rect 26056 12378 26108 12384
rect 26068 12347 26096 12378
rect 26436 11762 26464 14010
rect 26608 13184 26660 13190
rect 26608 13126 26660 13132
rect 26620 12850 26648 13126
rect 26608 12844 26660 12850
rect 26608 12786 26660 12792
rect 25872 11756 25924 11762
rect 25872 11698 25924 11704
rect 26056 11756 26108 11762
rect 26056 11698 26108 11704
rect 26424 11756 26476 11762
rect 26424 11698 26476 11704
rect 25412 11552 25464 11558
rect 25412 11494 25464 11500
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 25228 10056 25280 10062
rect 25228 9998 25280 10004
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25964 10056 26016 10062
rect 25964 9998 26016 10004
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 23572 9172 23624 9178
rect 23572 9114 23624 9120
rect 22192 8900 22244 8906
rect 22192 8842 22244 8848
rect 23388 8900 23440 8906
rect 23388 8842 23440 8848
rect 21640 8832 21692 8838
rect 21640 8774 21692 8780
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 21652 8566 21680 8774
rect 22020 8634 22048 8774
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 21640 8560 21692 8566
rect 21640 8502 21692 8508
rect 20904 8492 20956 8498
rect 20904 8434 20956 8440
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 20720 8016 20772 8022
rect 20720 7958 20772 7964
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20536 7812 20588 7818
rect 20536 7754 20588 7760
rect 20456 7546 20484 7754
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20076 7472 20128 7478
rect 20076 7414 20128 7420
rect 20640 7410 20668 7822
rect 20824 7546 20852 8026
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20916 7410 20944 7686
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19444 5370 19472 6054
rect 21916 5908 21968 5914
rect 21916 5850 21968 5856
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17880 4622 17908 5170
rect 21928 4622 21956 5850
rect 22204 5234 22232 8842
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 22928 8492 22980 8498
rect 22928 8434 22980 8440
rect 22940 8090 22968 8434
rect 23112 8288 23164 8294
rect 23112 8230 23164 8236
rect 23204 8288 23256 8294
rect 23204 8230 23256 8236
rect 23124 8090 23152 8230
rect 22928 8084 22980 8090
rect 22928 8026 22980 8032
rect 23112 8084 23164 8090
rect 23112 8026 23164 8032
rect 23216 7818 23244 8230
rect 23204 7812 23256 7818
rect 23204 7754 23256 7760
rect 23400 7478 23428 8570
rect 23584 8090 23612 9114
rect 24872 8974 24900 9862
rect 25240 9178 25268 9998
rect 25228 9172 25280 9178
rect 25228 9114 25280 9120
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 24492 8560 24544 8566
rect 24596 8548 24624 8910
rect 24676 8832 24728 8838
rect 24676 8774 24728 8780
rect 24688 8566 24716 8774
rect 24544 8520 24624 8548
rect 24492 8502 24544 8508
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 24596 7546 24624 8520
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24584 7540 24636 7546
rect 24584 7482 24636 7488
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 23400 5302 23428 7414
rect 24688 6798 24716 7822
rect 25332 7750 25360 9998
rect 25412 9988 25464 9994
rect 25412 9930 25464 9936
rect 25424 9654 25452 9930
rect 25412 9648 25464 9654
rect 25412 9590 25464 9596
rect 25424 8906 25452 9590
rect 25412 8900 25464 8906
rect 25412 8842 25464 8848
rect 25596 7812 25648 7818
rect 25596 7754 25648 7760
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25332 7478 25360 7686
rect 25608 7546 25636 7754
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25320 7472 25372 7478
rect 25320 7414 25372 7420
rect 25688 7472 25740 7478
rect 25688 7414 25740 7420
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24688 5370 24716 6734
rect 25320 6724 25372 6730
rect 25320 6666 25372 6672
rect 25332 6458 25360 6666
rect 25320 6452 25372 6458
rect 25320 6394 25372 6400
rect 25700 6322 25728 7414
rect 25976 6662 26004 9998
rect 26068 9994 26096 11698
rect 26436 10962 26464 11698
rect 26436 10934 26556 10962
rect 26424 10464 26476 10470
rect 26424 10406 26476 10412
rect 26436 10062 26464 10406
rect 26528 10062 26556 10934
rect 26712 10266 26740 14214
rect 26804 12918 26832 14282
rect 27160 13252 27212 13258
rect 27160 13194 27212 13200
rect 27172 12986 27200 13194
rect 27160 12980 27212 12986
rect 27160 12922 27212 12928
rect 26792 12912 26844 12918
rect 26792 12854 26844 12860
rect 27264 12442 27292 17546
rect 28172 16720 28224 16726
rect 28172 16662 28224 16668
rect 28184 15162 28212 16662
rect 28172 15156 28224 15162
rect 28172 15098 28224 15104
rect 28368 13530 28396 19994
rect 29012 19854 29040 20742
rect 29552 20528 29604 20534
rect 29552 20470 29604 20476
rect 29564 20330 29592 20470
rect 29552 20324 29604 20330
rect 29552 20266 29604 20272
rect 29000 19848 29052 19854
rect 29000 19790 29052 19796
rect 28448 18760 28500 18766
rect 28448 18702 28500 18708
rect 28460 17746 28488 18702
rect 28632 18284 28684 18290
rect 28632 18226 28684 18232
rect 28448 17740 28500 17746
rect 28448 17682 28500 17688
rect 28460 15026 28488 17682
rect 28644 17542 28672 18226
rect 29000 18080 29052 18086
rect 29000 18022 29052 18028
rect 29012 17814 29040 18022
rect 29000 17808 29052 17814
rect 29000 17750 29052 17756
rect 28632 17536 28684 17542
rect 28632 17478 28684 17484
rect 28540 16516 28592 16522
rect 28540 16458 28592 16464
rect 28552 16250 28580 16458
rect 28540 16244 28592 16250
rect 28540 16186 28592 16192
rect 28448 15020 28500 15026
rect 28448 14962 28500 14968
rect 28356 13524 28408 13530
rect 28356 13466 28408 13472
rect 27344 12844 27396 12850
rect 27344 12786 27396 12792
rect 26792 12436 26844 12442
rect 26792 12378 26844 12384
rect 27252 12436 27304 12442
rect 27356 12434 27384 12786
rect 28080 12708 28132 12714
rect 28080 12650 28132 12656
rect 28092 12442 28120 12650
rect 28080 12436 28132 12442
rect 27356 12406 27476 12434
rect 27252 12378 27304 12384
rect 26804 11898 26832 12378
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 26700 10260 26752 10266
rect 26700 10202 26752 10208
rect 26424 10056 26476 10062
rect 26424 9998 26476 10004
rect 26516 10056 26568 10062
rect 26516 9998 26568 10004
rect 26056 9988 26108 9994
rect 26056 9930 26108 9936
rect 26528 9586 26556 9998
rect 26516 9580 26568 9586
rect 26516 9522 26568 9528
rect 26148 9512 26200 9518
rect 26148 9454 26200 9460
rect 26160 8090 26188 9454
rect 26148 8084 26200 8090
rect 26148 8026 26200 8032
rect 26160 7546 26188 8026
rect 27448 7886 27476 12406
rect 28080 12378 28132 12384
rect 28460 12306 28488 14962
rect 28644 12918 28672 17478
rect 29460 16584 29512 16590
rect 29460 16526 29512 16532
rect 29000 16108 29052 16114
rect 29000 16050 29052 16056
rect 29012 15570 29040 16050
rect 29472 16046 29500 16526
rect 29092 16040 29144 16046
rect 29092 15982 29144 15988
rect 29460 16040 29512 16046
rect 29460 15982 29512 15988
rect 29000 15564 29052 15570
rect 29000 15506 29052 15512
rect 28724 15020 28776 15026
rect 28724 14962 28776 14968
rect 28736 14618 28764 14962
rect 28724 14612 28776 14618
rect 28724 14554 28776 14560
rect 29104 13802 29132 15982
rect 29092 13796 29144 13802
rect 29092 13738 29144 13744
rect 29104 13326 29132 13738
rect 29092 13320 29144 13326
rect 29092 13262 29144 13268
rect 29472 12986 29500 15982
rect 29564 15502 29592 20266
rect 29644 19848 29696 19854
rect 29644 19790 29696 19796
rect 29656 19310 29684 19790
rect 29644 19304 29696 19310
rect 29644 19246 29696 19252
rect 29656 18426 29684 19246
rect 29644 18420 29696 18426
rect 29644 18362 29696 18368
rect 29748 17678 29776 21422
rect 29828 21344 29880 21350
rect 29828 21286 29880 21292
rect 29840 20942 29868 21286
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 30748 20460 30800 20466
rect 30748 20402 30800 20408
rect 30012 20256 30064 20262
rect 30012 20198 30064 20204
rect 30024 19922 30052 20198
rect 30760 20058 30788 20402
rect 30748 20052 30800 20058
rect 30748 19994 30800 20000
rect 30012 19916 30064 19922
rect 30012 19858 30064 19864
rect 30944 18834 30972 21966
rect 31772 20534 31800 24006
rect 31760 20528 31812 20534
rect 31760 20470 31812 20476
rect 32324 20398 32352 24822
rect 32404 24812 32456 24818
rect 32404 24754 32456 24760
rect 32416 24070 32444 24754
rect 32496 24200 32548 24206
rect 32496 24142 32548 24148
rect 32404 24064 32456 24070
rect 32404 24006 32456 24012
rect 32508 23322 32536 24142
rect 32496 23316 32548 23322
rect 32496 23258 32548 23264
rect 32600 22094 32628 25094
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35992 23724 36044 23730
rect 35992 23666 36044 23672
rect 32956 23656 33008 23662
rect 32956 23598 33008 23604
rect 34612 23656 34664 23662
rect 34612 23598 34664 23604
rect 32968 22098 32996 23598
rect 33324 22636 33376 22642
rect 33324 22578 33376 22584
rect 33416 22636 33468 22642
rect 33416 22578 33468 22584
rect 33336 22234 33364 22578
rect 33324 22228 33376 22234
rect 33324 22170 33376 22176
rect 32508 22066 32628 22094
rect 32956 22092 33008 22098
rect 31116 20392 31168 20398
rect 31116 20334 31168 20340
rect 32312 20392 32364 20398
rect 32312 20334 32364 20340
rect 30380 18828 30432 18834
rect 30380 18770 30432 18776
rect 30932 18828 30984 18834
rect 30932 18770 30984 18776
rect 30196 18624 30248 18630
rect 30196 18566 30248 18572
rect 29736 17672 29788 17678
rect 29736 17614 29788 17620
rect 30208 17338 30236 18566
rect 30392 17746 30420 18770
rect 31024 18760 31076 18766
rect 31024 18702 31076 18708
rect 30840 18692 30892 18698
rect 30840 18634 30892 18640
rect 30852 18290 30880 18634
rect 31036 18630 31064 18702
rect 31024 18624 31076 18630
rect 31024 18566 31076 18572
rect 31036 18290 31064 18566
rect 30840 18284 30892 18290
rect 30840 18226 30892 18232
rect 31024 18284 31076 18290
rect 31024 18226 31076 18232
rect 30380 17740 30432 17746
rect 30380 17682 30432 17688
rect 30196 17332 30248 17338
rect 30196 17274 30248 17280
rect 30932 16448 30984 16454
rect 30932 16390 30984 16396
rect 30944 16182 30972 16390
rect 30932 16176 30984 16182
rect 30932 16118 30984 16124
rect 30656 16108 30708 16114
rect 30656 16050 30708 16056
rect 30668 15706 30696 16050
rect 30656 15700 30708 15706
rect 30656 15642 30708 15648
rect 30196 15564 30248 15570
rect 30196 15506 30248 15512
rect 29552 15496 29604 15502
rect 29552 15438 29604 15444
rect 30208 13326 30236 15506
rect 30944 15026 30972 16118
rect 30564 15020 30616 15026
rect 30564 14962 30616 14968
rect 30932 15020 30984 15026
rect 30932 14962 30984 14968
rect 30576 14618 30604 14962
rect 30564 14612 30616 14618
rect 30564 14554 30616 14560
rect 30380 14544 30432 14550
rect 30380 14486 30432 14492
rect 30196 13320 30248 13326
rect 30196 13262 30248 13268
rect 29736 13184 29788 13190
rect 29736 13126 29788 13132
rect 29460 12980 29512 12986
rect 29460 12922 29512 12928
rect 28632 12912 28684 12918
rect 28632 12854 28684 12860
rect 28448 12300 28500 12306
rect 28448 12242 28500 12248
rect 28460 11898 28488 12242
rect 28540 12164 28592 12170
rect 28540 12106 28592 12112
rect 28448 11892 28500 11898
rect 28448 11834 28500 11840
rect 28264 11824 28316 11830
rect 28264 11766 28316 11772
rect 27988 11552 28040 11558
rect 27988 11494 28040 11500
rect 28000 10266 28028 11494
rect 27988 10260 28040 10266
rect 27988 10202 28040 10208
rect 28276 9994 28304 11766
rect 28552 11762 28580 12106
rect 29748 11762 29776 13126
rect 30208 12918 30236 13262
rect 30196 12912 30248 12918
rect 30196 12854 30248 12860
rect 30208 11830 30236 12854
rect 30392 12306 30420 14486
rect 30472 13252 30524 13258
rect 30472 13194 30524 13200
rect 30380 12300 30432 12306
rect 30380 12242 30432 12248
rect 30288 12232 30340 12238
rect 30288 12174 30340 12180
rect 30196 11824 30248 11830
rect 30196 11766 30248 11772
rect 28540 11756 28592 11762
rect 28540 11698 28592 11704
rect 29736 11756 29788 11762
rect 29736 11698 29788 11704
rect 29184 11688 29236 11694
rect 29184 11630 29236 11636
rect 29092 11620 29144 11626
rect 29092 11562 29144 11568
rect 29104 10062 29132 11562
rect 29196 10810 29224 11630
rect 29920 11144 29972 11150
rect 29920 11086 29972 11092
rect 29932 10810 29960 11086
rect 29184 10804 29236 10810
rect 29184 10746 29236 10752
rect 29920 10804 29972 10810
rect 29920 10746 29972 10752
rect 30208 10062 30236 11766
rect 29092 10056 29144 10062
rect 29092 9998 29144 10004
rect 30196 10056 30248 10062
rect 30196 9998 30248 10004
rect 27620 9988 27672 9994
rect 27620 9930 27672 9936
rect 28264 9988 28316 9994
rect 28264 9930 28316 9936
rect 29000 9988 29052 9994
rect 29000 9930 29052 9936
rect 27436 7880 27488 7886
rect 27436 7822 27488 7828
rect 26148 7540 26200 7546
rect 26148 7482 26200 7488
rect 25964 6656 26016 6662
rect 25964 6598 26016 6604
rect 25976 6458 26004 6598
rect 25964 6452 26016 6458
rect 25964 6394 26016 6400
rect 27448 6390 27476 7822
rect 27632 6882 27660 9930
rect 29012 9654 29040 9930
rect 29104 9722 29132 9998
rect 29644 9920 29696 9926
rect 29644 9862 29696 9868
rect 29092 9716 29144 9722
rect 29092 9658 29144 9664
rect 29656 9654 29684 9862
rect 27712 9648 27764 9654
rect 27712 9590 27764 9596
rect 29000 9648 29052 9654
rect 29000 9590 29052 9596
rect 29644 9648 29696 9654
rect 29644 9590 29696 9596
rect 27724 9178 27752 9590
rect 28816 9444 28868 9450
rect 28816 9386 28868 9392
rect 27712 9172 27764 9178
rect 27712 9114 27764 9120
rect 28828 7478 28856 9386
rect 29736 9376 29788 9382
rect 29736 9318 29788 9324
rect 29748 8974 29776 9318
rect 29092 8968 29144 8974
rect 29092 8910 29144 8916
rect 29736 8968 29788 8974
rect 29736 8910 29788 8916
rect 29104 8566 29132 8910
rect 29644 8900 29696 8906
rect 29644 8842 29696 8848
rect 29656 8634 29684 8842
rect 29644 8628 29696 8634
rect 29644 8570 29696 8576
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 29748 7546 29776 8910
rect 29828 8900 29880 8906
rect 29828 8842 29880 8848
rect 29840 8090 29868 8842
rect 30208 8566 30236 9998
rect 30300 9994 30328 12174
rect 30484 10062 30512 13194
rect 30576 13190 30604 14554
rect 30944 14550 30972 14962
rect 30932 14544 30984 14550
rect 30932 14486 30984 14492
rect 30564 13184 30616 13190
rect 30564 13126 30616 13132
rect 30576 12102 30604 13126
rect 31128 12850 31156 20334
rect 32324 19854 32352 20334
rect 32312 19848 32364 19854
rect 32312 19790 32364 19796
rect 32508 19786 32536 22066
rect 32956 22034 33008 22040
rect 33428 22030 33456 22578
rect 34520 22432 34572 22438
rect 34520 22374 34572 22380
rect 34532 22030 34560 22374
rect 34624 22166 34652 23598
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 36004 23186 36032 23666
rect 36084 23520 36136 23526
rect 36084 23462 36136 23468
rect 35992 23180 36044 23186
rect 35992 23122 36044 23128
rect 36096 22642 36124 23462
rect 36176 23248 36228 23254
rect 36176 23190 36228 23196
rect 36084 22636 36136 22642
rect 36084 22578 36136 22584
rect 35900 22568 35952 22574
rect 36188 22522 36216 23190
rect 36360 23112 36412 23118
rect 36360 23054 36412 23060
rect 36372 22778 36400 23054
rect 36360 22772 36412 22778
rect 36360 22714 36412 22720
rect 36268 22636 36320 22642
rect 36268 22578 36320 22584
rect 35900 22510 35952 22516
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34612 22160 34664 22166
rect 34612 22102 34664 22108
rect 33416 22024 33468 22030
rect 33416 21966 33468 21972
rect 34520 22024 34572 22030
rect 34520 21966 34572 21972
rect 33324 20052 33376 20058
rect 33324 19994 33376 20000
rect 33336 19922 33364 19994
rect 33324 19916 33376 19922
rect 33324 19858 33376 19864
rect 32496 19780 32548 19786
rect 32496 19722 32548 19728
rect 31208 19712 31260 19718
rect 31208 19654 31260 19660
rect 32220 19712 32272 19718
rect 32220 19654 32272 19660
rect 31220 19310 31248 19654
rect 32232 19446 32260 19654
rect 32220 19440 32272 19446
rect 32220 19382 32272 19388
rect 31208 19304 31260 19310
rect 31208 19246 31260 19252
rect 32232 18426 32260 19382
rect 32220 18420 32272 18426
rect 32220 18362 32272 18368
rect 32232 17678 32260 18362
rect 32220 17672 32272 17678
rect 32220 17614 32272 17620
rect 31208 15904 31260 15910
rect 31208 15846 31260 15852
rect 31220 15366 31248 15846
rect 31392 15428 31444 15434
rect 31392 15370 31444 15376
rect 31208 15360 31260 15366
rect 31208 15302 31260 15308
rect 31220 14958 31248 15302
rect 31208 14952 31260 14958
rect 31208 14894 31260 14900
rect 31220 14822 31248 14894
rect 31208 14816 31260 14822
rect 31208 14758 31260 14764
rect 31116 12844 31168 12850
rect 31116 12786 31168 12792
rect 30840 12164 30892 12170
rect 30840 12106 30892 12112
rect 30564 12096 30616 12102
rect 30564 12038 30616 12044
rect 30576 11694 30604 12038
rect 30852 11898 30880 12106
rect 30840 11892 30892 11898
rect 30840 11834 30892 11840
rect 31404 11762 31432 15370
rect 31852 15088 31904 15094
rect 31852 15030 31904 15036
rect 31864 14346 31892 15030
rect 31852 14340 31904 14346
rect 31852 14282 31904 14288
rect 31864 11830 31892 14282
rect 32404 13932 32456 13938
rect 32404 13874 32456 13880
rect 32312 13864 32364 13870
rect 32312 13806 32364 13812
rect 32324 13530 32352 13806
rect 32312 13524 32364 13530
rect 32312 13466 32364 13472
rect 32128 13252 32180 13258
rect 32128 13194 32180 13200
rect 32140 12102 32168 13194
rect 32324 12850 32352 13466
rect 32312 12844 32364 12850
rect 32312 12786 32364 12792
rect 32128 12096 32180 12102
rect 32128 12038 32180 12044
rect 31852 11824 31904 11830
rect 31852 11766 31904 11772
rect 31392 11756 31444 11762
rect 31392 11698 31444 11704
rect 30564 11688 30616 11694
rect 30564 11630 30616 11636
rect 31116 10464 31168 10470
rect 31116 10406 31168 10412
rect 30472 10056 30524 10062
rect 30472 9998 30524 10004
rect 30288 9988 30340 9994
rect 30288 9930 30340 9936
rect 29920 8560 29972 8566
rect 29920 8502 29972 8508
rect 30196 8560 30248 8566
rect 30196 8502 30248 8508
rect 29828 8084 29880 8090
rect 29828 8026 29880 8032
rect 29736 7540 29788 7546
rect 29736 7482 29788 7488
rect 28816 7472 28868 7478
rect 28816 7414 28868 7420
rect 27540 6854 27660 6882
rect 27436 6384 27488 6390
rect 27436 6326 27488 6332
rect 25688 6316 25740 6322
rect 25688 6258 25740 6264
rect 27540 5778 27568 6854
rect 27528 5772 27580 5778
rect 27528 5714 27580 5720
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 23388 5296 23440 5302
rect 23388 5238 23440 5244
rect 22192 5228 22244 5234
rect 22192 5170 22244 5176
rect 22100 5024 22152 5030
rect 22100 4966 22152 4972
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 21916 4616 21968 4622
rect 21916 4558 21968 4564
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17696 4146 17724 4422
rect 17880 4282 17908 4558
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 17868 4276 17920 4282
rect 17868 4218 17920 4224
rect 19444 4146 19472 4422
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 22112 4146 22140 4966
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19800 4140 19852 4146
rect 19800 4082 19852 4088
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17972 3194 18000 3334
rect 18432 3194 18460 4082
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 17972 2446 18000 3130
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 18800 2650 18828 2994
rect 19076 2990 19104 3538
rect 19352 3058 19380 3878
rect 19812 3738 19840 4082
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 20916 3534 20944 3878
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 18788 2644 18840 2650
rect 18788 2586 18840 2592
rect 20088 2446 20116 2994
rect 20916 2446 20944 3470
rect 22204 3058 22232 5170
rect 22284 4752 22336 4758
rect 22284 4694 22336 4700
rect 22296 4214 22324 4694
rect 27540 4622 27568 5714
rect 28080 5636 28132 5642
rect 28080 5578 28132 5584
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 27160 4616 27212 4622
rect 27160 4558 27212 4564
rect 27528 4616 27580 4622
rect 27528 4558 27580 4564
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 22836 4480 22888 4486
rect 22836 4422 22888 4428
rect 22664 4282 22692 4422
rect 22652 4276 22704 4282
rect 22652 4218 22704 4224
rect 22284 4208 22336 4214
rect 22284 4150 22336 4156
rect 22848 3534 22876 4422
rect 23020 4276 23072 4282
rect 23020 4218 23072 4224
rect 22560 3528 22612 3534
rect 22560 3470 22612 3476
rect 22836 3528 22888 3534
rect 22836 3470 22888 3476
rect 22572 3194 22600 3470
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 23032 2446 23060 4218
rect 23216 3738 23244 4558
rect 26792 4548 26844 4554
rect 26792 4490 26844 4496
rect 23572 4480 23624 4486
rect 23572 4422 23624 4428
rect 23848 4480 23900 4486
rect 23848 4422 23900 4428
rect 23584 3738 23612 4422
rect 23860 4146 23888 4422
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 24584 4140 24636 4146
rect 24584 4082 24636 4088
rect 24596 3738 24624 4082
rect 26424 4072 26476 4078
rect 26424 4014 26476 4020
rect 25044 3936 25096 3942
rect 25044 3878 25096 3884
rect 23204 3732 23256 3738
rect 23204 3674 23256 3680
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 23756 3732 23808 3738
rect 23756 3674 23808 3680
rect 24584 3732 24636 3738
rect 24584 3674 24636 3680
rect 23216 3534 23244 3674
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 23768 2446 23796 3674
rect 25056 3602 25084 3878
rect 25044 3596 25096 3602
rect 25044 3538 25096 3544
rect 25056 2446 25084 3538
rect 26436 3466 26464 4014
rect 26804 3738 26832 4490
rect 27172 4146 27200 4558
rect 27804 4480 27856 4486
rect 27804 4422 27856 4428
rect 27160 4140 27212 4146
rect 27160 4082 27212 4088
rect 27436 3936 27488 3942
rect 27436 3878 27488 3884
rect 27448 3738 27476 3878
rect 27816 3738 27844 4422
rect 26792 3732 26844 3738
rect 26792 3674 26844 3680
rect 27436 3732 27488 3738
rect 27436 3674 27488 3680
rect 27804 3732 27856 3738
rect 27804 3674 27856 3680
rect 26424 3460 26476 3466
rect 26424 3402 26476 3408
rect 26436 2922 26464 3402
rect 26424 2916 26476 2922
rect 26424 2858 26476 2864
rect 27448 2446 27476 3674
rect 27896 3596 27948 3602
rect 27896 3538 27948 3544
rect 27908 2922 27936 3538
rect 28092 3194 28120 5578
rect 28632 5568 28684 5574
rect 28632 5510 28684 5516
rect 28644 4758 28672 5510
rect 28828 5302 28856 7414
rect 29932 5370 29960 8502
rect 30208 7886 30236 8502
rect 30300 8362 30328 9930
rect 30656 9920 30708 9926
rect 30656 9862 30708 9868
rect 30668 8498 30696 9862
rect 31128 9178 31156 10406
rect 30932 9172 30984 9178
rect 30932 9114 30984 9120
rect 31116 9172 31168 9178
rect 31116 9114 31168 9120
rect 30944 8634 30972 9114
rect 30932 8628 30984 8634
rect 30932 8570 30984 8576
rect 30656 8492 30708 8498
rect 30656 8434 30708 8440
rect 30748 8492 30800 8498
rect 30748 8434 30800 8440
rect 30288 8356 30340 8362
rect 30288 8298 30340 8304
rect 30196 7880 30248 7886
rect 30196 7822 30248 7828
rect 30760 7342 30788 8434
rect 31128 7818 31156 9114
rect 31404 7954 31432 11698
rect 31484 11552 31536 11558
rect 31484 11494 31536 11500
rect 31496 11218 31524 11494
rect 31484 11212 31536 11218
rect 31484 11154 31536 11160
rect 32140 10742 32168 12038
rect 32416 11898 32444 13874
rect 32404 11892 32456 11898
rect 32404 11834 32456 11840
rect 32508 11762 32536 19722
rect 33140 18828 33192 18834
rect 33140 18770 33192 18776
rect 32772 18284 32824 18290
rect 32772 18226 32824 18232
rect 32588 18148 32640 18154
rect 32588 18090 32640 18096
rect 32600 17678 32628 18090
rect 32784 18086 32812 18226
rect 32864 18216 32916 18222
rect 32864 18158 32916 18164
rect 32772 18080 32824 18086
rect 32772 18022 32824 18028
rect 32588 17672 32640 17678
rect 32588 17614 32640 17620
rect 32680 17604 32732 17610
rect 32680 17546 32732 17552
rect 32692 17202 32720 17546
rect 32680 17196 32732 17202
rect 32680 17138 32732 17144
rect 32784 15162 32812 18022
rect 32876 16794 32904 18158
rect 33048 17672 33100 17678
rect 33048 17614 33100 17620
rect 32864 16788 32916 16794
rect 32864 16730 32916 16736
rect 32772 15156 32824 15162
rect 32772 15098 32824 15104
rect 33060 15026 33088 17614
rect 33152 17338 33180 18770
rect 33336 18290 33364 19858
rect 33324 18284 33376 18290
rect 33324 18226 33376 18232
rect 33428 17882 33456 21966
rect 34532 21486 34560 21966
rect 35348 21956 35400 21962
rect 35348 21898 35400 21904
rect 35072 21888 35124 21894
rect 35072 21830 35124 21836
rect 35084 21690 35112 21830
rect 35072 21684 35124 21690
rect 35072 21626 35124 21632
rect 35360 21486 35388 21898
rect 35912 21554 35940 22510
rect 36004 22506 36216 22522
rect 35992 22500 36216 22506
rect 36044 22494 36216 22500
rect 35992 22442 36044 22448
rect 36004 22094 36032 22442
rect 36004 22066 36124 22094
rect 35900 21548 35952 21554
rect 35900 21490 35952 21496
rect 34520 21480 34572 21486
rect 34520 21422 34572 21428
rect 34796 21480 34848 21486
rect 34796 21422 34848 21428
rect 35348 21480 35400 21486
rect 35348 21422 35400 21428
rect 35808 21480 35860 21486
rect 35808 21422 35860 21428
rect 34808 21010 34836 21422
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35360 21078 35388 21422
rect 35348 21072 35400 21078
rect 35348 21014 35400 21020
rect 35820 21010 35848 21422
rect 34796 21004 34848 21010
rect 34796 20946 34848 20952
rect 35808 21004 35860 21010
rect 35808 20946 35860 20952
rect 34808 20058 34836 20946
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34796 20052 34848 20058
rect 34796 19994 34848 20000
rect 35348 19848 35400 19854
rect 35348 19790 35400 19796
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 33784 18760 33836 18766
rect 33784 18702 33836 18708
rect 33600 18216 33652 18222
rect 33600 18158 33652 18164
rect 33416 17876 33468 17882
rect 33416 17818 33468 17824
rect 33612 17746 33640 18158
rect 33600 17740 33652 17746
rect 33600 17682 33652 17688
rect 33140 17332 33192 17338
rect 33140 17274 33192 17280
rect 33416 17264 33468 17270
rect 33612 17218 33640 17682
rect 33796 17678 33824 18702
rect 35360 18698 35388 19790
rect 35716 18760 35768 18766
rect 35716 18702 35768 18708
rect 35348 18692 35400 18698
rect 35348 18634 35400 18640
rect 34796 18216 34848 18222
rect 34796 18158 34848 18164
rect 34808 17678 34836 18158
rect 35360 18154 35388 18634
rect 35728 18358 35756 18702
rect 35716 18352 35768 18358
rect 35716 18294 35768 18300
rect 35716 18216 35768 18222
rect 35820 18170 35848 20946
rect 35912 20874 35940 21490
rect 36096 21146 36124 22066
rect 36176 21480 36228 21486
rect 36176 21422 36228 21428
rect 36084 21140 36136 21146
rect 36084 21082 36136 21088
rect 36188 20942 36216 21422
rect 36176 20936 36228 20942
rect 36176 20878 36228 20884
rect 35900 20868 35952 20874
rect 35900 20810 35952 20816
rect 35912 19514 35940 20810
rect 36188 19922 36216 20878
rect 36280 20058 36308 22578
rect 37188 22024 37240 22030
rect 37188 21966 37240 21972
rect 38016 22024 38068 22030
rect 38016 21966 38068 21972
rect 36728 21956 36780 21962
rect 36728 21898 36780 21904
rect 36636 21616 36688 21622
rect 36636 21558 36688 21564
rect 36648 21010 36676 21558
rect 36636 21004 36688 21010
rect 36636 20946 36688 20952
rect 36740 20874 36768 21898
rect 37200 21894 37228 21966
rect 37188 21888 37240 21894
rect 37188 21830 37240 21836
rect 38028 21622 38056 21966
rect 38016 21616 38068 21622
rect 38016 21558 38068 21564
rect 36728 20868 36780 20874
rect 36728 20810 36780 20816
rect 36268 20052 36320 20058
rect 36268 19994 36320 20000
rect 36176 19916 36228 19922
rect 36176 19858 36228 19864
rect 35992 19848 36044 19854
rect 35992 19790 36044 19796
rect 36544 19848 36596 19854
rect 36544 19790 36596 19796
rect 35900 19508 35952 19514
rect 35900 19450 35952 19456
rect 36004 18766 36032 19790
rect 36452 19780 36504 19786
rect 36452 19722 36504 19728
rect 36176 19372 36228 19378
rect 36176 19314 36228 19320
rect 36084 19304 36136 19310
rect 36084 19246 36136 19252
rect 36096 18902 36124 19246
rect 36084 18896 36136 18902
rect 36084 18838 36136 18844
rect 35992 18760 36044 18766
rect 35992 18702 36044 18708
rect 36004 18426 36032 18702
rect 36188 18426 36216 19314
rect 36464 18766 36492 19722
rect 36556 19242 36584 19790
rect 36544 19236 36596 19242
rect 36544 19178 36596 19184
rect 36452 18760 36504 18766
rect 36452 18702 36504 18708
rect 35992 18420 36044 18426
rect 35992 18362 36044 18368
rect 36176 18420 36228 18426
rect 36176 18362 36228 18368
rect 36464 18358 36492 18702
rect 36452 18352 36504 18358
rect 36452 18294 36504 18300
rect 35768 18164 35848 18170
rect 35716 18158 35848 18164
rect 35348 18148 35400 18154
rect 35728 18142 35848 18158
rect 35348 18090 35400 18096
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 33784 17672 33836 17678
rect 33784 17614 33836 17620
rect 34796 17672 34848 17678
rect 34796 17614 34848 17620
rect 33416 17206 33468 17212
rect 33232 17128 33284 17134
rect 33232 17070 33284 17076
rect 33244 16590 33272 17070
rect 33232 16584 33284 16590
rect 33232 16526 33284 16532
rect 33428 16454 33456 17206
rect 33520 17202 33640 17218
rect 33508 17196 33640 17202
rect 33560 17190 33640 17196
rect 33508 17138 33560 17144
rect 33508 17060 33560 17066
rect 33508 17002 33560 17008
rect 33520 16590 33548 17002
rect 33796 16794 33824 17614
rect 34808 17202 34836 17614
rect 34796 17196 34848 17202
rect 34796 17138 34848 17144
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 33784 16788 33836 16794
rect 33784 16730 33836 16736
rect 33508 16584 33560 16590
rect 33508 16526 33560 16532
rect 34336 16584 34388 16590
rect 34336 16526 34388 16532
rect 33416 16448 33468 16454
rect 33416 16390 33468 16396
rect 33428 15706 33456 16390
rect 34348 15706 34376 16526
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 33416 15700 33468 15706
rect 33416 15642 33468 15648
rect 34336 15700 34388 15706
rect 34336 15642 34388 15648
rect 34888 15564 34940 15570
rect 34888 15506 34940 15512
rect 33692 15496 33744 15502
rect 33692 15438 33744 15444
rect 34704 15496 34756 15502
rect 34704 15438 34756 15444
rect 33048 15020 33100 15026
rect 33048 14962 33100 14968
rect 33508 15020 33560 15026
rect 33508 14962 33560 14968
rect 33060 14618 33088 14962
rect 33520 14906 33548 14962
rect 33704 14906 33732 15438
rect 34520 15156 34572 15162
rect 34520 15098 34572 15104
rect 33520 14878 33732 14906
rect 34532 14890 34560 15098
rect 34612 15088 34664 15094
rect 34612 15030 34664 15036
rect 33704 14822 33732 14878
rect 34520 14884 34572 14890
rect 34520 14826 34572 14832
rect 33600 14816 33652 14822
rect 33600 14758 33652 14764
rect 33692 14816 33744 14822
rect 33692 14758 33744 14764
rect 33048 14612 33100 14618
rect 33048 14554 33100 14560
rect 33612 14278 33640 14758
rect 34532 14414 34560 14826
rect 34520 14408 34572 14414
rect 34520 14350 34572 14356
rect 34624 14346 34652 15030
rect 34716 14958 34744 15438
rect 34796 15428 34848 15434
rect 34796 15370 34848 15376
rect 34704 14952 34756 14958
rect 34704 14894 34756 14900
rect 34808 14618 34836 15370
rect 34900 15026 34928 15506
rect 35164 15360 35216 15366
rect 35164 15302 35216 15308
rect 35176 15094 35204 15302
rect 35164 15088 35216 15094
rect 35164 15030 35216 15036
rect 34888 15020 34940 15026
rect 34888 14962 34940 14968
rect 34900 14822 34928 14962
rect 35360 14958 35388 18090
rect 35900 16516 35952 16522
rect 35900 16458 35952 16464
rect 35912 16250 35940 16458
rect 35900 16244 35952 16250
rect 35900 16186 35952 16192
rect 36360 16108 36412 16114
rect 36360 16050 36412 16056
rect 35900 15972 35952 15978
rect 35900 15914 35952 15920
rect 35912 15026 35940 15914
rect 36372 15570 36400 16050
rect 36464 16046 36492 18294
rect 36740 16794 36768 20810
rect 38108 20392 38160 20398
rect 38108 20334 38160 20340
rect 38120 19961 38148 20334
rect 38106 19952 38162 19961
rect 38106 19887 38162 19896
rect 36912 19848 36964 19854
rect 36912 19790 36964 19796
rect 36924 19378 36952 19790
rect 36912 19372 36964 19378
rect 36912 19314 36964 19320
rect 36728 16788 36780 16794
rect 36728 16730 36780 16736
rect 36924 16590 36952 19314
rect 36912 16584 36964 16590
rect 36912 16526 36964 16532
rect 37188 16584 37240 16590
rect 37188 16526 37240 16532
rect 36636 16108 36688 16114
rect 36636 16050 36688 16056
rect 36452 16040 36504 16046
rect 36452 15982 36504 15988
rect 36464 15858 36492 15982
rect 36648 15978 36676 16050
rect 36636 15972 36688 15978
rect 36636 15914 36688 15920
rect 36464 15830 36584 15858
rect 36360 15564 36412 15570
rect 36360 15506 36412 15512
rect 36556 15502 36584 15830
rect 36924 15638 36952 16526
rect 37200 16250 37228 16526
rect 37832 16516 37884 16522
rect 37832 16458 37884 16464
rect 37844 16250 37872 16458
rect 37188 16244 37240 16250
rect 37188 16186 37240 16192
rect 37832 16244 37884 16250
rect 37832 16186 37884 16192
rect 37372 16176 37424 16182
rect 37372 16118 37424 16124
rect 37384 15706 37412 16118
rect 37372 15700 37424 15706
rect 37372 15642 37424 15648
rect 36912 15632 36964 15638
rect 36912 15574 36964 15580
rect 36544 15496 36596 15502
rect 36544 15438 36596 15444
rect 36912 15496 36964 15502
rect 36912 15438 36964 15444
rect 37188 15496 37240 15502
rect 37188 15438 37240 15444
rect 35900 15020 35952 15026
rect 35900 14962 35952 14968
rect 35348 14952 35400 14958
rect 35348 14894 35400 14900
rect 34888 14816 34940 14822
rect 34888 14758 34940 14764
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35360 14634 35388 14894
rect 35808 14816 35860 14822
rect 35808 14758 35860 14764
rect 34796 14612 34848 14618
rect 34796 14554 34848 14560
rect 35268 14606 35388 14634
rect 35268 14414 35296 14606
rect 35820 14414 35848 14758
rect 35256 14408 35308 14414
rect 35256 14350 35308 14356
rect 35808 14408 35860 14414
rect 35808 14350 35860 14356
rect 34612 14340 34664 14346
rect 34612 14282 34664 14288
rect 33600 14272 33652 14278
rect 33600 14214 33652 14220
rect 35268 14074 35296 14350
rect 35912 14278 35940 14962
rect 36556 14822 36584 15438
rect 36924 15162 36952 15438
rect 36912 15156 36964 15162
rect 36912 15098 36964 15104
rect 36176 14816 36228 14822
rect 36176 14758 36228 14764
rect 36544 14816 36596 14822
rect 36544 14758 36596 14764
rect 36188 14414 36216 14758
rect 37200 14618 37228 15438
rect 37188 14612 37240 14618
rect 37188 14554 37240 14560
rect 36176 14408 36228 14414
rect 36176 14350 36228 14356
rect 35900 14272 35952 14278
rect 35900 14214 35952 14220
rect 32680 14068 32732 14074
rect 32680 14010 32732 14016
rect 35256 14068 35308 14074
rect 35256 14010 35308 14016
rect 32692 11898 32720 14010
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 36188 12986 36216 14350
rect 36176 12980 36228 12986
rect 36176 12922 36228 12928
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 32680 11892 32732 11898
rect 32680 11834 32732 11840
rect 32588 11824 32640 11830
rect 32588 11766 32640 11772
rect 32496 11756 32548 11762
rect 32496 11698 32548 11704
rect 32128 10736 32180 10742
rect 32128 10678 32180 10684
rect 32508 8430 32536 11698
rect 32600 11354 32628 11766
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 32588 11348 32640 11354
rect 32588 11290 32640 11296
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 32496 8424 32548 8430
rect 32496 8366 32548 8372
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 31392 7948 31444 7954
rect 31392 7890 31444 7896
rect 31116 7812 31168 7818
rect 31116 7754 31168 7760
rect 30748 7336 30800 7342
rect 30748 7278 30800 7284
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 29920 5364 29972 5370
rect 29920 5306 29972 5312
rect 28816 5296 28868 5302
rect 28816 5238 28868 5244
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 28632 4752 28684 4758
rect 28632 4694 28684 4700
rect 28724 4752 28776 4758
rect 28724 4694 28776 4700
rect 28644 3738 28672 4694
rect 28736 3942 28764 4694
rect 28816 4684 28868 4690
rect 28816 4626 28868 4632
rect 28828 4282 28856 4626
rect 28816 4276 28868 4282
rect 28816 4218 28868 4224
rect 28724 3936 28776 3942
rect 28724 3878 28776 3884
rect 28632 3732 28684 3738
rect 28632 3674 28684 3680
rect 28736 3670 28764 3878
rect 28724 3664 28776 3670
rect 28724 3606 28776 3612
rect 28828 3602 28856 4218
rect 29092 4140 29144 4146
rect 29092 4082 29144 4088
rect 29104 3738 29132 4082
rect 32312 3936 32364 3942
rect 32312 3878 32364 3884
rect 29092 3732 29144 3738
rect 29092 3674 29144 3680
rect 28908 3664 28960 3670
rect 28908 3606 28960 3612
rect 28816 3596 28868 3602
rect 28816 3538 28868 3544
rect 28920 3534 28948 3606
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 28080 3188 28132 3194
rect 28080 3130 28132 3136
rect 27896 2916 27948 2922
rect 27896 2858 27948 2864
rect 27908 2446 27936 2858
rect 28920 2514 28948 3470
rect 28908 2508 28960 2514
rect 28908 2450 28960 2456
rect 32324 2446 32352 3878
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 39120 2984 39172 2990
rect 39120 2926 39172 2932
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 20904 2440 20956 2446
rect 20904 2382 20956 2388
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 25044 2440 25096 2446
rect 25044 2382 25096 2388
rect 27436 2440 27488 2446
rect 27436 2382 27488 2388
rect 27896 2440 27948 2446
rect 27896 2382 27948 2388
rect 32312 2440 32364 2446
rect 32312 2382 32364 2388
rect 33232 2440 33284 2446
rect 33232 2382 33284 2388
rect 34704 2440 34756 2446
rect 34704 2382 34756 2388
rect 36176 2440 36228 2446
rect 36176 2382 36228 2388
rect 37648 2440 37700 2446
rect 37648 2382 37700 2388
rect 2320 2372 2372 2378
rect 2320 2314 2372 2320
rect 3792 2372 3844 2378
rect 3792 2314 3844 2320
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 2332 800 2360 2314
rect 3804 800 3832 2314
rect 5276 800 5304 2314
rect 6748 800 6776 2382
rect 8220 800 8248 2382
rect 9692 800 9720 2382
rect 11164 800 11192 2382
rect 12636 800 12664 2382
rect 14108 800 14136 2382
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 17040 2372 17092 2378
rect 17040 2314 17092 2320
rect 18512 2372 18564 2378
rect 18512 2314 18564 2320
rect 19984 2372 20036 2378
rect 19984 2314 20036 2320
rect 21456 2372 21508 2378
rect 21456 2314 21508 2320
rect 22928 2372 22980 2378
rect 22928 2314 22980 2320
rect 24400 2372 24452 2378
rect 24400 2314 24452 2320
rect 25872 2372 25924 2378
rect 25872 2314 25924 2320
rect 27344 2372 27396 2378
rect 27344 2314 27396 2320
rect 28816 2372 28868 2378
rect 28816 2314 28868 2320
rect 30288 2372 30340 2378
rect 30288 2314 30340 2320
rect 31760 2372 31812 2378
rect 31760 2314 31812 2320
rect 15580 800 15608 2314
rect 17052 800 17080 2314
rect 18524 800 18552 2314
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2314
rect 21468 800 21496 2314
rect 22940 800 22968 2314
rect 24412 800 24440 2314
rect 25884 800 25912 2314
rect 27356 800 27384 2314
rect 28828 800 28856 2314
rect 30300 800 30328 2314
rect 31772 800 31800 2314
rect 33244 800 33272 2382
rect 34716 800 34744 2382
rect 36188 800 36216 2382
rect 37660 800 37688 2382
rect 39132 800 39160 2926
rect 846 0 902 800
rect 2318 0 2374 800
rect 3790 0 3846 800
rect 5262 0 5318 800
rect 6734 0 6790 800
rect 8206 0 8262 800
rect 9678 0 9734 800
rect 11150 0 11206 800
rect 12622 0 12678 800
rect 14094 0 14150 800
rect 15566 0 15622 800
rect 17038 0 17094 800
rect 18510 0 18566 800
rect 19982 0 20038 800
rect 21454 0 21510 800
rect 22926 0 22982 800
rect 24398 0 24454 800
rect 25870 0 25926 800
rect 27342 0 27398 800
rect 28814 0 28870 800
rect 30286 0 30342 800
rect 31758 0 31814 800
rect 33230 0 33286 800
rect 34702 0 34758 800
rect 36174 0 36230 800
rect 37646 0 37702 800
rect 39118 0 39174 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 20166 35012 20222 35048
rect 20166 34992 20168 35012
rect 20168 34992 20220 35012
rect 20220 34992 20222 35012
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 20810 35028 20812 35048
rect 20812 35028 20864 35048
rect 20864 35028 20866 35048
rect 20810 34992 20866 35028
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 24490 29044 24492 29064
rect 24492 29044 24544 29064
rect 24544 29044 24546 29064
rect 24490 29008 24546 29044
rect 27710 31728 27766 31784
rect 27618 29008 27674 29064
rect 28170 22636 28226 22672
rect 28170 22616 28172 22636
rect 28172 22616 28224 22636
rect 28224 22616 28226 22636
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 38106 19896 38162 19952
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 20161 35050 20227 35053
rect 20805 35050 20871 35053
rect 20161 35048 20871 35050
rect 20161 34992 20166 35048
rect 20222 34992 20810 35048
rect 20866 34992 20871 35048
rect 20161 34990 20871 34992
rect 20161 34987 20227 34990
rect 20805 34987 20871 34990
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 27705 31786 27771 31789
rect 28206 31786 28212 31788
rect 27705 31784 28212 31786
rect 27705 31728 27710 31784
rect 27766 31728 28212 31784
rect 27705 31726 28212 31728
rect 27705 31723 27771 31726
rect 28206 31724 28212 31726
rect 28276 31724 28282 31788
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 24485 29066 24551 29069
rect 27613 29066 27679 29069
rect 24485 29064 27679 29066
rect 24485 29008 24490 29064
rect 24546 29008 27618 29064
rect 27674 29008 27679 29064
rect 24485 29006 27679 29008
rect 24485 29003 24551 29006
rect 27613 29003 27679 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 28165 22676 28231 22677
rect 28165 22674 28212 22676
rect 28120 22672 28212 22674
rect 28120 22616 28170 22672
rect 28120 22614 28212 22616
rect 28165 22612 28212 22614
rect 28276 22612 28282 22676
rect 28165 22611 28231 22612
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 38101 19954 38167 19957
rect 39200 19954 40000 19984
rect 38101 19952 40000 19954
rect 38101 19896 38106 19952
rect 38162 19896 40000 19952
rect 38101 19894 40000 19896
rect 38101 19891 38167 19894
rect 39200 19864 40000 19894
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 28212 31724 28276 31788
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 28212 22672 28276 22676
rect 28212 22616 28226 22672
rect 28226 22616 28276 22672
rect 28212 22612 28276 22616
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 28211 31788 28277 31789
rect 28211 31724 28212 31788
rect 28276 31724 28277 31788
rect 28211 31723 28277 31724
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 28214 22677 28274 31723
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 28211 22676 28277 22677
rect 28211 22612 28212 22676
rect 28276 22612 28277 22676
rect 28211 22611 28277 22612
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25576 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1666464484
transform 1 0 18400 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20
timestamp 1666464484
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37
timestamp 1666464484
transform 1 0 4508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1666464484
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77
timestamp 1666464484
transform 1 0 8188 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93
timestamp 1666464484
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118
timestamp 1666464484
transform 1 0 11960 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129
timestamp 1666464484
transform 1 0 12972 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146
timestamp 1666464484
transform 1 0 14536 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1666464484
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1666464484
transform 1 0 17020 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_180
timestamp 1666464484
transform 1 0 17664 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1666464484
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1666464484
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_212
timestamp 1666464484
transform 1 0 20608 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1666464484
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_237
timestamp 1666464484
transform 1 0 22908 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_244
timestamp 1666464484
transform 1 0 23552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_261
timestamp 1666464484
transform 1 0 25116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_269
timestamp 1666464484
transform 1 0 25852 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1666464484
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_285
timestamp 1666464484
transform 1 0 27324 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_292
timestamp 1666464484
transform 1 0 27968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1666464484
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1666464484
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_317
timestamp 1666464484
transform 1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_327
timestamp 1666464484
transform 1 0 31188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1666464484
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1666464484
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_345
timestamp 1666464484
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_349
timestamp 1666464484
transform 1 0 33212 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_353
timestamp 1666464484
transform 1 0 33580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1666464484
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1666464484
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_370
timestamp 1666464484
transform 1 0 35144 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1666464484
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_393
timestamp 1666464484
transform 1 0 37260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_397
timestamp 1666464484
transform 1 0 37628 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_401
timestamp 1666464484
transform 1 0 37996 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_11
timestamp 1666464484
transform 1 0 2116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_23
timestamp 1666464484
transform 1 0 3220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_35
timestamp 1666464484
transform 1 0 4324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 1666464484
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_100
timestamp 1666464484
transform 1 0 10304 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_150
timestamp 1666464484
transform 1 0 14904 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1666464484
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_180
timestamp 1666464484
transform 1 0 17664 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_197
timestamp 1666464484
transform 1 0 19228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_209
timestamp 1666464484
transform 1 0 20332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp 1666464484
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_233
timestamp 1666464484
transform 1 0 22540 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1666464484
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1666464484
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1666464484
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1666464484
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1666464484
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1666464484
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1666464484
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1666464484
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1666464484
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1666464484
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1666464484
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1666464484
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1666464484
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1666464484
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1666464484
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1666464484
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 1666464484
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_401
timestamp 1666464484
transform 1 0 37996 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1666464484
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_69
timestamp 1666464484
transform 1 0 7452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1666464484
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_107
timestamp 1666464484
transform 1 0 10948 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_119
timestamp 1666464484
transform 1 0 12052 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_131
timestamp 1666464484
transform 1 0 13156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_158
timestamp 1666464484
transform 1 0 15640 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_166
timestamp 1666464484
transform 1 0 16376 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_184
timestamp 1666464484
transform 1 0 18032 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_212
timestamp 1666464484
transform 1 0 20608 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_224
timestamp 1666464484
transform 1 0 21712 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_232
timestamp 1666464484
transform 1 0 22448 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp 1666464484
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_264
timestamp 1666464484
transform 1 0 25392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_268
timestamp 1666464484
transform 1 0 25760 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_274
timestamp 1666464484
transform 1 0 26312 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_280
timestamp 1666464484
transform 1 0 26864 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_295
timestamp 1666464484
transform 1 0 28244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp 1666464484
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1666464484
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1666464484
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1666464484
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1666464484
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1666464484
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1666464484
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1666464484
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1666464484
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1666464484
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_401
timestamp 1666464484
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1666464484
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1666464484
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666464484
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_75
timestamp 1666464484
transform 1 0 8004 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_83
timestamp 1666464484
transform 1 0 8740 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_141
timestamp 1666464484
transform 1 0 14076 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_174
timestamp 1666464484
transform 1 0 17112 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_196
timestamp 1666464484
transform 1 0 19136 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1666464484
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1666464484
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_263
timestamp 1666464484
transform 1 0 25300 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_271
timestamp 1666464484
transform 1 0 26036 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1666464484
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_299
timestamp 1666464484
transform 1 0 28612 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_319
timestamp 1666464484
transform 1 0 30452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_331
timestamp 1666464484
transform 1 0 31556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1666464484
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1666464484
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1666464484
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1666464484
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1666464484
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1666464484
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1666464484
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1666464484
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1666464484
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_62
timestamp 1666464484
transform 1 0 6808 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_70
timestamp 1666464484
transform 1 0 7544 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1666464484
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_96
timestamp 1666464484
transform 1 0 9936 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_104
timestamp 1666464484
transform 1 0 10672 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_115
timestamp 1666464484
transform 1 0 11684 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_123
timestamp 1666464484
transform 1 0 12420 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_129
timestamp 1666464484
transform 1 0 12972 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1666464484
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_147
timestamp 1666464484
transform 1 0 14628 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_154
timestamp 1666464484
transform 1 0 15272 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_166
timestamp 1666464484
transform 1 0 16376 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_178
timestamp 1666464484
transform 1 0 17480 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_184
timestamp 1666464484
transform 1 0 18032 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_204
timestamp 1666464484
transform 1 0 19872 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_216
timestamp 1666464484
transform 1 0 20976 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_231
timestamp 1666464484
transform 1 0 22356 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_241
timestamp 1666464484
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1666464484
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_258
timestamp 1666464484
transform 1 0 24840 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_270
timestamp 1666464484
transform 1 0 25944 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_274
timestamp 1666464484
transform 1 0 26312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_291
timestamp 1666464484
transform 1 0 27876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1666464484
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1666464484
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1666464484
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1666464484
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1666464484
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1666464484
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1666464484
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1666464484
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1666464484
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1666464484
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_401
timestamp 1666464484
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_39
timestamp 1666464484
transform 1 0 4692 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_45
timestamp 1666464484
transform 1 0 5244 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1666464484
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666464484
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_99
timestamp 1666464484
transform 1 0 10212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_185
timestamp 1666464484
transform 1 0 18124 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_206
timestamp 1666464484
transform 1 0 20056 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_218
timestamp 1666464484
transform 1 0 21160 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_231
timestamp 1666464484
transform 1 0 22356 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_239
timestamp 1666464484
transform 1 0 23092 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_262
timestamp 1666464484
transform 1 0 25208 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp 1666464484
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1666464484
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_319
timestamp 1666464484
transform 1 0 30452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_331
timestamp 1666464484
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1666464484
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1666464484
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1666464484
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1666464484
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1666464484
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1666464484
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1666464484
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1666464484
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1666464484
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_37
timestamp 1666464484
transform 1 0 4508 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_62
timestamp 1666464484
transform 1 0 6808 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_74
timestamp 1666464484
transform 1 0 7912 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1666464484
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_103
timestamp 1666464484
transform 1 0 10580 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_115
timestamp 1666464484
transform 1 0 11684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_127
timestamp 1666464484
transform 1 0 12788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1666464484
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1666464484
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1666464484
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1666464484
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1666464484
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_289
timestamp 1666464484
transform 1 0 27692 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1666464484
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1666464484
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1666464484
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1666464484
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1666464484
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1666464484
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1666464484
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1666464484
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1666464484
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1666464484
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1666464484
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1666464484
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1666464484
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_124
timestamp 1666464484
transform 1 0 12512 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_136
timestamp 1666464484
transform 1 0 13616 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_148
timestamp 1666464484
transform 1 0 14720 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_160
timestamp 1666464484
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1666464484
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1666464484
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_261
timestamp 1666464484
transform 1 0 25116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1666464484
transform 1 0 25852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1666464484
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1666464484
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1666464484
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1666464484
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1666464484
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1666464484
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1666464484
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1666464484
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1666464484
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1666464484
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1666464484
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1666464484
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1666464484
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1666464484
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_57
timestamp 1666464484
transform 1 0 6348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_67
timestamp 1666464484
transform 1 0 7268 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 1666464484
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_101
timestamp 1666464484
transform 1 0 10396 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_111
timestamp 1666464484
transform 1 0 11316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_123
timestamp 1666464484
transform 1 0 12420 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1666464484
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_161
timestamp 1666464484
transform 1 0 15916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_173
timestamp 1666464484
transform 1 0 17020 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_185
timestamp 1666464484
transform 1 0 18124 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp 1666464484
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1666464484
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1666464484
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1666464484
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1666464484
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_271
timestamp 1666464484
transform 1 0 26036 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_283
timestamp 1666464484
transform 1 0 27140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_295
timestamp 1666464484
transform 1 0 28244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1666464484
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1666464484
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1666464484
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1666464484
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1666464484
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1666464484
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1666464484
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1666464484
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1666464484
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1666464484
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1666464484
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1666464484
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1666464484
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1666464484
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1666464484
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666464484
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_68
timestamp 1666464484
transform 1 0 7360 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_80
timestamp 1666464484
transform 1 0 8464 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_88
timestamp 1666464484
transform 1 0 9200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_119
timestamp 1666464484
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_123
timestamp 1666464484
transform 1 0 12420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_135
timestamp 1666464484
transform 1 0 13524 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_143
timestamp 1666464484
transform 1 0 14260 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_160
timestamp 1666464484
transform 1 0 15824 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_185
timestamp 1666464484
transform 1 0 18124 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_206
timestamp 1666464484
transform 1 0 20056 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_216
timestamp 1666464484
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_237
timestamp 1666464484
transform 1 0 22908 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_241
timestamp 1666464484
transform 1 0 23276 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_262
timestamp 1666464484
transform 1 0 25208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_272
timestamp 1666464484
transform 1 0 26128 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1666464484
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_319
timestamp 1666464484
transform 1 0 30452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_331
timestamp 1666464484
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1666464484
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1666464484
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1666464484
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1666464484
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1666464484
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1666464484
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1666464484
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1666464484
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1666464484
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1666464484
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_35
timestamp 1666464484
transform 1 0 4324 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_43
timestamp 1666464484
transform 1 0 5060 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_64
timestamp 1666464484
transform 1 0 6992 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1666464484
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_107
timestamp 1666464484
transform 1 0 10948 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_116
timestamp 1666464484
transform 1 0 11776 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_128
timestamp 1666464484
transform 1 0 12880 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_161
timestamp 1666464484
transform 1 0 15916 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_171
timestamp 1666464484
transform 1 0 16836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_183
timestamp 1666464484
transform 1 0 17940 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_187
timestamp 1666464484
transform 1 0 18308 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1666464484
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_215
timestamp 1666464484
transform 1 0 20884 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_227
timestamp 1666464484
transform 1 0 21988 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_235
timestamp 1666464484
transform 1 0 22724 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_242
timestamp 1666464484
transform 1 0 23368 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1666464484
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_257
timestamp 1666464484
transform 1 0 24748 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_274
timestamp 1666464484
transform 1 0 26312 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_286
timestamp 1666464484
transform 1 0 27416 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_298
timestamp 1666464484
transform 1 0 28520 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1666464484
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1666464484
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_317
timestamp 1666464484
transform 1 0 30268 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_329
timestamp 1666464484
transform 1 0 31372 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_341
timestamp 1666464484
transform 1 0 32476 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_353
timestamp 1666464484
transform 1 0 33580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp 1666464484
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1666464484
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1666464484
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1666464484
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1666464484
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_21
timestamp 1666464484
transform 1 0 3036 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_33
timestamp 1666464484
transform 1 0 4140 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_37
timestamp 1666464484
transform 1 0 4508 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1666464484
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_64
timestamp 1666464484
transform 1 0 6992 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_76
timestamp 1666464484
transform 1 0 8096 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_88
timestamp 1666464484
transform 1 0 9200 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1666464484
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_133
timestamp 1666464484
transform 1 0 13340 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_141
timestamp 1666464484
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 1666464484
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_177
timestamp 1666464484
transform 1 0 17388 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_185
timestamp 1666464484
transform 1 0 18124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_193
timestamp 1666464484
transform 1 0 18860 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_213
timestamp 1666464484
transform 1 0 20700 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1666464484
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_233
timestamp 1666464484
transform 1 0 22540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_252
timestamp 1666464484
transform 1 0 24288 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1666464484
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1666464484
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_299
timestamp 1666464484
transform 1 0 28612 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_316
timestamp 1666464484
transform 1 0 30176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_326
timestamp 1666464484
transform 1 0 31096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1666464484
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1666464484
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1666464484
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1666464484
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1666464484
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1666464484
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1666464484
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1666464484
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1666464484
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1666464484
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_159
timestamp 1666464484
transform 1 0 15732 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_169
timestamp 1666464484
transform 1 0 16652 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_181
timestamp 1666464484
transform 1 0 17756 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1666464484
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1666464484
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_229
timestamp 1666464484
transform 1 0 22172 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_241
timestamp 1666464484
transform 1 0 23276 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1666464484
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_271
timestamp 1666464484
transform 1 0 26036 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_283
timestamp 1666464484
transform 1 0 27140 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_289
timestamp 1666464484
transform 1 0 27692 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1666464484
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1666464484
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_327
timestamp 1666464484
transform 1 0 31188 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_339
timestamp 1666464484
transform 1 0 32292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_351
timestamp 1666464484
transform 1 0 33396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1666464484
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1666464484
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1666464484
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1666464484
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_401
timestamp 1666464484
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_15
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_20
timestamp 1666464484
transform 1 0 2944 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_32
timestamp 1666464484
transform 1 0 4048 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_44
timestamp 1666464484
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_159
timestamp 1666464484
transform 1 0 15732 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_189
timestamp 1666464484
transform 1 0 18492 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_207
timestamp 1666464484
transform 1 0 20148 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_218
timestamp 1666464484
transform 1 0 21160 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1666464484
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1666464484
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_261
timestamp 1666464484
transform 1 0 25116 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1666464484
transform 1 0 25852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1666464484
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_289
timestamp 1666464484
transform 1 0 27692 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_306
timestamp 1666464484
transform 1 0 29256 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_330
timestamp 1666464484
transform 1 0 31464 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1666464484
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1666464484
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1666464484
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1666464484
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1666464484
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1666464484
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1666464484
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1666464484
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1666464484
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666464484
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_47
timestamp 1666464484
transform 1 0 5428 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_59
timestamp 1666464484
transform 1 0 6532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_71
timestamp 1666464484
transform 1 0 7636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_103
timestamp 1666464484
transform 1 0 10580 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_115
timestamp 1666464484
transform 1 0 11684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_127
timestamp 1666464484
transform 1 0 12788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_205
timestamp 1666464484
transform 1 0 19964 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1666464484
transform 1 0 20700 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_234
timestamp 1666464484
transform 1 0 22632 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_246
timestamp 1666464484
transform 1 0 23736 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_257
timestamp 1666464484
transform 1 0 24748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_264
timestamp 1666464484
transform 1 0 25392 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_279
timestamp 1666464484
transform 1 0 26772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_287
timestamp 1666464484
transform 1 0 27508 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_296
timestamp 1666464484
transform 1 0 28336 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1666464484
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_317
timestamp 1666464484
transform 1 0 30268 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_327
timestamp 1666464484
transform 1 0 31188 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_339
timestamp 1666464484
transform 1 0 32292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_351
timestamp 1666464484
transform 1 0 33396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1666464484
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1666464484
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1666464484
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1666464484
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1666464484
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_46
timestamp 1666464484
transform 1 0 5336 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1666464484
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_89
timestamp 1666464484
transform 1 0 9292 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1666464484
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666464484
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_185
timestamp 1666464484
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_206
timestamp 1666464484
transform 1 0 20056 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1666464484
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1666464484
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1666464484
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1666464484
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1666464484
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666464484
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1666464484
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_319
timestamp 1666464484
transform 1 0 30452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_331
timestamp 1666464484
transform 1 0 31556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1666464484
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1666464484
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1666464484
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1666464484
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1666464484
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1666464484
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1666464484
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1666464484
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1666464484
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_41
timestamp 1666464484
transform 1 0 4876 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_63
timestamp 1666464484
transform 1 0 6900 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_75
timestamp 1666464484
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_103
timestamp 1666464484
transform 1 0 10580 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_115
timestamp 1666464484
transform 1 0 11684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_127
timestamp 1666464484
transform 1 0 12788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_159
timestamp 1666464484
transform 1 0 15732 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_171
timestamp 1666464484
transform 1 0 16836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_183
timestamp 1666464484
transform 1 0 17940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666464484
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666464484
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_221
timestamp 1666464484
transform 1 0 21436 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_243
timestamp 1666464484
transform 1 0 23460 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666464484
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1666464484
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1666464484
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1666464484
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1666464484
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1666464484
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1666464484
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_321
timestamp 1666464484
transform 1 0 30636 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_346
timestamp 1666464484
transform 1 0 32936 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_358
timestamp 1666464484
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1666464484
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1666464484
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1666464484
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1666464484
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1666464484
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1666464484
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1666464484
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1666464484
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1666464484
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_125
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666464484
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666464484
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666464484
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666464484
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666464484
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1666464484
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_254
timestamp 1666464484
transform 1 0 24472 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_266
timestamp 1666464484
transform 1 0 25576 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1666464484
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_293
timestamp 1666464484
transform 1 0 28060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_301
timestamp 1666464484
transform 1 0 28796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_324
timestamp 1666464484
transform 1 0 30912 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1666464484
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1666464484
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_345
timestamp 1666464484
transform 1 0 32844 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_357
timestamp 1666464484
transform 1 0 33948 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_369
timestamp 1666464484
transform 1 0 35052 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_381
timestamp 1666464484
transform 1 0 36156 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_389
timestamp 1666464484
transform 1 0 36892 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1666464484
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1666464484
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1666464484
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_37
timestamp 1666464484
transform 1 0 4508 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_45
timestamp 1666464484
transform 1 0 5244 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_63
timestamp 1666464484
transform 1 0 6900 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_75
timestamp 1666464484
transform 1 0 8004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_103
timestamp 1666464484
transform 1 0 10580 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_115
timestamp 1666464484
transform 1 0 11684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_127
timestamp 1666464484
transform 1 0 12788 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_131
timestamp 1666464484
transform 1 0 13156 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1666464484
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_159
timestamp 1666464484
transform 1 0 15732 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_171
timestamp 1666464484
transform 1 0 16836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_183
timestamp 1666464484
transform 1 0 17940 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1666464484
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_207
timestamp 1666464484
transform 1 0 20148 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_215
timestamp 1666464484
transform 1 0 20884 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_222
timestamp 1666464484
transform 1 0 21528 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_242
timestamp 1666464484
transform 1 0 23368 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1666464484
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_275
timestamp 1666464484
transform 1 0 26404 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_284
timestamp 1666464484
transform 1 0 27232 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_292
timestamp 1666464484
transform 1 0 27968 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1666464484
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1666464484
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1666464484
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_321
timestamp 1666464484
transform 1 0 30636 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_343
timestamp 1666464484
transform 1 0 32660 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_355
timestamp 1666464484
transform 1 0 33764 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1666464484
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1666464484
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1666464484
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1666464484
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1666464484
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_19
timestamp 1666464484
transform 1 0 2852 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_29
timestamp 1666464484
transform 1 0 3772 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_37
timestamp 1666464484
transform 1 0 4508 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1666464484
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_89
timestamp 1666464484
transform 1 0 9292 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1666464484
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_121
timestamp 1666464484
transform 1 0 12236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_129
timestamp 1666464484
transform 1 0 12972 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1666464484
transform 1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666464484
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_179
timestamp 1666464484
transform 1 0 17572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_191
timestamp 1666464484
transform 1 0 18676 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_203
timestamp 1666464484
transform 1 0 19780 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_215
timestamp 1666464484
transform 1 0 20884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666464484
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_237
timestamp 1666464484
transform 1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_241
timestamp 1666464484
transform 1 0 23276 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_262
timestamp 1666464484
transform 1 0 25208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_272
timestamp 1666464484
transform 1 0 26128 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_289
timestamp 1666464484
transform 1 0 27692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_297
timestamp 1666464484
transform 1 0 28428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_319
timestamp 1666464484
transform 1 0 30452 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_331
timestamp 1666464484
transform 1 0 31556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1666464484
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1666464484
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_358
timestamp 1666464484
transform 1 0 34040 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_370
timestamp 1666464484
transform 1 0 35144 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_382
timestamp 1666464484
transform 1 0 36248 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_390
timestamp 1666464484
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1666464484
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1666464484
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1666464484
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1666464484
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_37
timestamp 1666464484
transform 1 0 4508 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_49
timestamp 1666464484
transform 1 0 5612 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_61
timestamp 1666464484
transform 1 0 6716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1666464484
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666464484
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_163
timestamp 1666464484
transform 1 0 16100 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_171
timestamp 1666464484
transform 1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_185
timestamp 1666464484
transform 1 0 18124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1666464484
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_204
timestamp 1666464484
transform 1 0 19872 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1666464484
transform 1 0 20608 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_234
timestamp 1666464484
transform 1 0 22632 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_246
timestamp 1666464484
transform 1 0 23736 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_271
timestamp 1666464484
transform 1 0 26036 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_279
timestamp 1666464484
transform 1 0 26772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_291
timestamp 1666464484
transform 1 0 27876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1666464484
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1666464484
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1666464484
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_317
timestamp 1666464484
transform 1 0 30268 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_325
timestamp 1666464484
transform 1 0 31004 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_347
timestamp 1666464484
transform 1 0 33028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_359
timestamp 1666464484
transform 1 0 34132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1666464484
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1666464484
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1666464484
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1666464484
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1666464484
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_12
timestamp 1666464484
transform 1 0 2208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_25
timestamp 1666464484
transform 1 0 3404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_35
timestamp 1666464484
transform 1 0 4324 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_42
timestamp 1666464484
transform 1 0 4968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1666464484
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_99
timestamp 1666464484
transform 1 0 10212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_144
timestamp 1666464484
transform 1 0 14352 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_154
timestamp 1666464484
transform 1 0 15272 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1666464484
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_182
timestamp 1666464484
transform 1 0 17848 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_190
timestamp 1666464484
transform 1 0 18584 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_200
timestamp 1666464484
transform 1 0 19504 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_212
timestamp 1666464484
transform 1 0 20608 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_233
timestamp 1666464484
transform 1 0 22540 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_241
timestamp 1666464484
transform 1 0 23276 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_262
timestamp 1666464484
transform 1 0 25208 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_274
timestamp 1666464484
transform 1 0 26312 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1666464484
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1666464484
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1666464484
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1666464484
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1666464484
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1666464484
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_356
timestamp 1666464484
transform 1 0 33856 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_368
timestamp 1666464484
transform 1 0 34960 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_380
timestamp 1666464484
transform 1 0 36064 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1666464484
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1666464484
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_14
timestamp 1666464484
transform 1 0 2392 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1666464484
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666464484
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666464484
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_121
timestamp 1666464484
transform 1 0 12236 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_129
timestamp 1666464484
transform 1 0 12972 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1666464484
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_153
timestamp 1666464484
transform 1 0 15180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_166
timestamp 1666464484
transform 1 0 16376 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_177
timestamp 1666464484
transform 1 0 17388 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1666464484
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_205
timestamp 1666464484
transform 1 0 19964 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_213
timestamp 1666464484
transform 1 0 20700 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_225
timestamp 1666464484
transform 1 0 21804 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_243
timestamp 1666464484
transform 1 0 23460 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1666464484
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_265
timestamp 1666464484
transform 1 0 25484 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_281
timestamp 1666464484
transform 1 0 26956 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_293
timestamp 1666464484
transform 1 0 28060 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_305
timestamp 1666464484
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1666464484
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1666464484
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1666464484
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1666464484
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1666464484
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1666464484
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1666464484
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_373
timestamp 1666464484
transform 1 0 35420 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_377
timestamp 1666464484
transform 1 0 35788 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_382
timestamp 1666464484
transform 1 0 36248 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_394
timestamp 1666464484
transform 1 0 37352 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_406
timestamp 1666464484
transform 1 0 38456 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_24
timestamp 1666464484
transform 1 0 3312 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_31
timestamp 1666464484
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_43
timestamp 1666464484
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666464484
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_137
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_145
timestamp 1666464484
transform 1 0 14444 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_157
timestamp 1666464484
transform 1 0 15548 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1666464484
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_182
timestamp 1666464484
transform 1 0 17848 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_190
timestamp 1666464484
transform 1 0 18584 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_201
timestamp 1666464484
transform 1 0 19596 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_209
timestamp 1666464484
transform 1 0 20332 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1666464484
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1666464484
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1666464484
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_261
timestamp 1666464484
transform 1 0 25116 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_269
timestamp 1666464484
transform 1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1666464484
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_293
timestamp 1666464484
transform 1 0 28060 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_301
timestamp 1666464484
transform 1 0 28796 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_313
timestamp 1666464484
transform 1 0 29900 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_319
timestamp 1666464484
transform 1 0 30452 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_327
timestamp 1666464484
transform 1 0 31188 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1666464484
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_337
timestamp 1666464484
transform 1 0 32108 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_346
timestamp 1666464484
transform 1 0 32936 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_358
timestamp 1666464484
transform 1 0 34040 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_371
timestamp 1666464484
transform 1 0 35236 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_380
timestamp 1666464484
transform 1 0 36064 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_389
timestamp 1666464484
transform 1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1666464484
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1666464484
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1666464484
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_53
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_61
timestamp 1666464484
transform 1 0 6716 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_67
timestamp 1666464484
transform 1 0 7268 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1666464484
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666464484
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1666464484
transform 1 0 9476 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666464484
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_165
timestamp 1666464484
transform 1 0 16284 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_186
timestamp 1666464484
transform 1 0 18216 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1666464484
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_204
timestamp 1666464484
transform 1 0 19872 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_216
timestamp 1666464484
transform 1 0 20976 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_228
timestamp 1666464484
transform 1 0 22080 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_240
timestamp 1666464484
transform 1 0 23184 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_264
timestamp 1666464484
transform 1 0 25392 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_284
timestamp 1666464484
transform 1 0 27232 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_296
timestamp 1666464484
transform 1 0 28336 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1666464484
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_317
timestamp 1666464484
transform 1 0 30268 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_327
timestamp 1666464484
transform 1 0 31188 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_339
timestamp 1666464484
transform 1 0 32292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_351
timestamp 1666464484
transform 1 0 33396 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1666464484
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1666464484
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_372
timestamp 1666464484
transform 1 0 35328 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_380
timestamp 1666464484
transform 1 0 36064 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_390
timestamp 1666464484
transform 1 0 36984 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_397
timestamp 1666464484
transform 1 0 37628 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1666464484
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666464484
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_39
timestamp 1666464484
transform 1 0 4692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_47
timestamp 1666464484
transform 1 0 5428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1666464484
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_80
timestamp 1666464484
transform 1 0 8464 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1666464484
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_139
timestamp 1666464484
transform 1 0 13892 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_145
timestamp 1666464484
transform 1 0 14444 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_154
timestamp 1666464484
transform 1 0 15272 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1666464484
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_180
timestamp 1666464484
transform 1 0 17664 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666464484
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_205
timestamp 1666464484
transform 1 0 19964 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_213
timestamp 1666464484
transform 1 0 20700 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1666464484
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1666464484
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1666464484
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_261
timestamp 1666464484
transform 1 0 25116 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1666464484
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_293
timestamp 1666464484
transform 1 0 28060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_297
timestamp 1666464484
transform 1 0 28428 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_304
timestamp 1666464484
transform 1 0 29072 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_325
timestamp 1666464484
transform 1 0 31004 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1666464484
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1666464484
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1666464484
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1666464484
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_373
timestamp 1666464484
transform 1 0 35420 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_380
timestamp 1666464484
transform 1 0 36064 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_389
timestamp 1666464484
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1666464484
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_400
timestamp 1666464484
transform 1 0 37904 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_406
timestamp 1666464484
transform 1 0 38456 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1666464484
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_41
timestamp 1666464484
transform 1 0 4876 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_64
timestamp 1666464484
transform 1 0 6992 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_74
timestamp 1666464484
transform 1 0 7912 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1666464484
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_121
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_129
timestamp 1666464484
transform 1 0 12972 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1666464484
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_171
timestamp 1666464484
transform 1 0 16836 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_181
timestamp 1666464484
transform 1 0 17756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1666464484
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_209
timestamp 1666464484
transform 1 0 20332 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_215
timestamp 1666464484
transform 1 0 20884 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_232
timestamp 1666464484
transform 1 0 22448 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_240
timestamp 1666464484
transform 1 0 23184 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1666464484
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_265
timestamp 1666464484
transform 1 0 25484 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_274
timestamp 1666464484
transform 1 0 26312 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_286
timestamp 1666464484
transform 1 0 27416 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_298
timestamp 1666464484
transform 1 0 28520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1666464484
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1666464484
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_328
timestamp 1666464484
transform 1 0 31280 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_340
timestamp 1666464484
transform 1 0 32384 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_346
timestamp 1666464484
transform 1 0 32936 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_353
timestamp 1666464484
transform 1 0 33580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_361
timestamp 1666464484
transform 1 0 34316 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1666464484
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_377
timestamp 1666464484
transform 1 0 35788 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_383
timestamp 1666464484
transform 1 0 36340 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_393
timestamp 1666464484
transform 1 0 37260 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_405
timestamp 1666464484
transform 1 0 38364 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_39
timestamp 1666464484
transform 1 0 4692 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1666464484
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_71
timestamp 1666464484
transform 1 0 7636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_83
timestamp 1666464484
transform 1 0 8740 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_100
timestamp 1666464484
transform 1 0 10304 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1666464484
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_142
timestamp 1666464484
transform 1 0 14168 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_155
timestamp 1666464484
transform 1 0 15364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_182
timestamp 1666464484
transform 1 0 17848 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_194
timestamp 1666464484
transform 1 0 18952 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_206
timestamp 1666464484
transform 1 0 20056 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_214
timestamp 1666464484
transform 1 0 20792 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1666464484
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_243
timestamp 1666464484
transform 1 0 23460 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_263
timestamp 1666464484
transform 1 0 25300 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_275
timestamp 1666464484
transform 1 0 26404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1666464484
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1666464484
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1666464484
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1666464484
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1666464484
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1666464484
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_337
timestamp 1666464484
transform 1 0 32108 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_344
timestamp 1666464484
transform 1 0 32752 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_356
timestamp 1666464484
transform 1 0 33856 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_368
timestamp 1666464484
transform 1 0 34960 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_380
timestamp 1666464484
transform 1 0 36064 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1666464484
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1666464484
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_15
timestamp 1666464484
transform 1 0 2484 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_22
timestamp 1666464484
transform 1 0 3128 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1666464484
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_108
timestamp 1666464484
transform 1 0 11040 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_120
timestamp 1666464484
transform 1 0 12144 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1666464484
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_175
timestamp 1666464484
transform 1 0 17204 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_183
timestamp 1666464484
transform 1 0 17940 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1666464484
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1666464484
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1666464484
transform 1 0 20700 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_234
timestamp 1666464484
transform 1 0 22632 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_244
timestamp 1666464484
transform 1 0 23552 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_262
timestamp 1666464484
transform 1 0 25208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_286
timestamp 1666464484
transform 1 0 27416 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_294
timestamp 1666464484
transform 1 0 28152 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1666464484
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1666464484
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_331
timestamp 1666464484
transform 1 0 31556 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_344
timestamp 1666464484
transform 1 0 32752 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1666464484
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1666464484
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1666464484
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1666464484
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1666464484
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1666464484
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_28
timestamp 1666464484
transform 1 0 3680 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_38
timestamp 1666464484
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1666464484
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_93
timestamp 1666464484
transform 1 0 9660 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1666464484
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_144
timestamp 1666464484
transform 1 0 14352 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_156
timestamp 1666464484
transform 1 0 15456 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_173
timestamp 1666464484
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_183
timestamp 1666464484
transform 1 0 17940 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_194
timestamp 1666464484
transform 1 0 18952 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666464484
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666464484
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_253
timestamp 1666464484
transform 1 0 24380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_277
timestamp 1666464484
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp 1666464484
transform 1 0 28060 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_319
timestamp 1666464484
transform 1 0 30452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_326
timestamp 1666464484
transform 1 0 31096 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1666464484
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_337
timestamp 1666464484
transform 1 0 32108 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_358
timestamp 1666464484
transform 1 0 34040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_371
timestamp 1666464484
transform 1 0 35236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_382
timestamp 1666464484
transform 1 0 36248 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1666464484
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1666464484
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1666464484
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_14
timestamp 1666464484
transform 1 0 2392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1666464484
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666464484
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_52
timestamp 1666464484
transform 1 0 5888 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_60
timestamp 1666464484
transform 1 0 6624 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_67
timestamp 1666464484
transform 1 0 7268 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1666464484
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_100
timestamp 1666464484
transform 1 0 10304 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_112
timestamp 1666464484
transform 1 0 11408 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_124
timestamp 1666464484
transform 1 0 12512 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1666464484
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_172
timestamp 1666464484
transform 1 0 16928 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_181
timestamp 1666464484
transform 1 0 17756 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1666464484
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666464484
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_221
timestamp 1666464484
transform 1 0 21436 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_233
timestamp 1666464484
transform 1 0 22540 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_239
timestamp 1666464484
transform 1 0 23092 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1666464484
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_281
timestamp 1666464484
transform 1 0 26956 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_293
timestamp 1666464484
transform 1 0 28060 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1666464484
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1666464484
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_320
timestamp 1666464484
transform 1 0 30544 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_332
timestamp 1666464484
transform 1 0 31648 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_340
timestamp 1666464484
transform 1 0 32384 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_356
timestamp 1666464484
transform 1 0 33856 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_365
timestamp 1666464484
transform 1 0 34684 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_373
timestamp 1666464484
transform 1 0 35420 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_386
timestamp 1666464484
transform 1 0 36616 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_398
timestamp 1666464484
transform 1 0 37720 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 1666464484
transform 1 0 38456 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_39
timestamp 1666464484
transform 1 0 4692 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_45
timestamp 1666464484
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1666464484
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_65
timestamp 1666464484
transform 1 0 7084 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_75
timestamp 1666464484
transform 1 0 8004 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_87
timestamp 1666464484
transform 1 0 9108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_99
timestamp 1666464484
transform 1 0 10212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_146
timestamp 1666464484
transform 1 0 14536 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_158
timestamp 1666464484
transform 1 0 15640 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1666464484
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1666464484
transform 1 0 17756 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_189
timestamp 1666464484
transform 1 0 18492 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_201
timestamp 1666464484
transform 1 0 19596 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_213
timestamp 1666464484
transform 1 0 20700 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1666464484
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_231
timestamp 1666464484
transform 1 0 22356 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_248
timestamp 1666464484
transform 1 0 23920 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_260
timestamp 1666464484
transform 1 0 25024 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1666464484
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_289
timestamp 1666464484
transform 1 0 27692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_301
timestamp 1666464484
transform 1 0 28796 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_309
timestamp 1666464484
transform 1 0 29532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1666464484
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1666464484
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1666464484
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1666464484
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1666464484
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_373
timestamp 1666464484
transform 1 0 35420 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_377
timestamp 1666464484
transform 1 0 35788 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_390
timestamp 1666464484
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1666464484
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1666464484
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1666464484
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666464484
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1666464484
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_149
timestamp 1666464484
transform 1 0 14812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_157
timestamp 1666464484
transform 1 0 15548 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_176
timestamp 1666464484
transform 1 0 17296 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_188
timestamp 1666464484
transform 1 0 18400 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_215
timestamp 1666464484
transform 1 0 20884 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_227
timestamp 1666464484
transform 1 0 21988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_239
timestamp 1666464484
transform 1 0 23092 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_243
timestamp 1666464484
transform 1 0 23460 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1666464484
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_265
timestamp 1666464484
transform 1 0 25484 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_291
timestamp 1666464484
transform 1 0 27876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_300
timestamp 1666464484
transform 1 0 28704 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1666464484
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_330
timestamp 1666464484
transform 1 0 31464 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_340
timestamp 1666464484
transform 1 0 32384 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_352
timestamp 1666464484
transform 1 0 33488 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1666464484
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_372
timestamp 1666464484
transform 1 0 35328 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_381
timestamp 1666464484
transform 1 0 36156 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_390
timestamp 1666464484
transform 1 0 36984 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_402
timestamp 1666464484
transform 1 0 38088 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_406
timestamp 1666464484
transform 1 0 38456 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_15
timestamp 1666464484
transform 1 0 2484 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_20
timestamp 1666464484
transform 1 0 2944 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_32
timestamp 1666464484
transform 1 0 4048 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_44
timestamp 1666464484
transform 1 0 5152 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_67
timestamp 1666464484
transform 1 0 7268 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_74
timestamp 1666464484
transform 1 0 7912 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_95
timestamp 1666464484
transform 1 0 9844 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1666464484
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_123
timestamp 1666464484
transform 1 0 12420 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_149
timestamp 1666464484
transform 1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_159
timestamp 1666464484
transform 1 0 15732 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_177
timestamp 1666464484
transform 1 0 17388 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_185
timestamp 1666464484
transform 1 0 18124 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_206
timestamp 1666464484
transform 1 0 20056 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_218
timestamp 1666464484
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_237
timestamp 1666464484
transform 1 0 22908 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_245
timestamp 1666464484
transform 1 0 23644 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_252
timestamp 1666464484
transform 1 0 24288 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_264
timestamp 1666464484
transform 1 0 25392 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_268
timestamp 1666464484
transform 1 0 25760 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1666464484
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1666464484
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1666464484
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1666464484
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_317
timestamp 1666464484
transform 1 0 30268 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_324
timestamp 1666464484
transform 1 0 30912 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1666464484
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1666464484
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1666464484
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1666464484
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1666464484
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1666464484
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_393
timestamp 1666464484
transform 1 0 37260 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_401
timestamp 1666464484
transform 1 0 37996 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1666464484
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1666464484
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_45
timestamp 1666464484
transform 1 0 5244 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_51
timestamp 1666464484
transform 1 0 5796 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_63
timestamp 1666464484
transform 1 0 6900 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_67
timestamp 1666464484
transform 1 0 7268 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_71
timestamp 1666464484
transform 1 0 7636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_102
timestamp 1666464484
transform 1 0 10488 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_117
timestamp 1666464484
transform 1 0 11868 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_124
timestamp 1666464484
transform 1 0 12512 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1666464484
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_152
timestamp 1666464484
transform 1 0 15088 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_178
timestamp 1666464484
transform 1 0 17480 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_190
timestamp 1666464484
transform 1 0 18584 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_209
timestamp 1666464484
transform 1 0 20332 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1666464484
transform 1 0 20700 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_234
timestamp 1666464484
transform 1 0 22632 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_246
timestamp 1666464484
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_265
timestamp 1666464484
transform 1 0 25484 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_291
timestamp 1666464484
transform 1 0 27876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_303
timestamp 1666464484
transform 1 0 28980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1666464484
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1666464484
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_314
timestamp 1666464484
transform 1 0 29992 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_326
timestamp 1666464484
transform 1 0 31096 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_338
timestamp 1666464484
transform 1 0 32200 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_350
timestamp 1666464484
transform 1 0 33304 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1666464484
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1666464484
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_374
timestamp 1666464484
transform 1 0 35512 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_387
timestamp 1666464484
transform 1 0 36708 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_399
timestamp 1666464484
transform 1 0 37812 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_7
timestamp 1666464484
transform 1 0 1748 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_29
timestamp 1666464484
transform 1 0 3772 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_38
timestamp 1666464484
transform 1 0 4600 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_50
timestamp 1666464484
transform 1 0 5704 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_65
timestamp 1666464484
transform 1 0 7084 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_72
timestamp 1666464484
transform 1 0 7728 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_84
timestamp 1666464484
transform 1 0 8832 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_94
timestamp 1666464484
transform 1 0 9752 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_102
timestamp 1666464484
transform 1 0 10488 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1666464484
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_117
timestamp 1666464484
transform 1 0 11868 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_124
timestamp 1666464484
transform 1 0 12512 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_128
timestamp 1666464484
transform 1 0 12880 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_149
timestamp 1666464484
transform 1 0 14812 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_157
timestamp 1666464484
transform 1 0 15548 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1666464484
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_185
timestamp 1666464484
transform 1 0 18124 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_206
timestamp 1666464484
transform 1 0 20056 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_214
timestamp 1666464484
transform 1 0 20792 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1666464484
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_237
timestamp 1666464484
transform 1 0 22908 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_256
timestamp 1666464484
transform 1 0 24656 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_268
timestamp 1666464484
transform 1 0 25760 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_289
timestamp 1666464484
transform 1 0 27692 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_297
timestamp 1666464484
transform 1 0 28428 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_309
timestamp 1666464484
transform 1 0 29532 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_321
timestamp 1666464484
transform 1 0 30636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_333
timestamp 1666464484
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_337
timestamp 1666464484
transform 1 0 32108 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_345
timestamp 1666464484
transform 1 0 32844 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_354
timestamp 1666464484
transform 1 0 33672 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_369
timestamp 1666464484
transform 1 0 35052 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_390
timestamp 1666464484
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1666464484
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1666464484
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_11
timestamp 1666464484
transform 1 0 2116 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_17
timestamp 1666464484
transform 1 0 2668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1666464484
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_36
timestamp 1666464484
transform 1 0 4416 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_48
timestamp 1666464484
transform 1 0 5520 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_54
timestamp 1666464484
transform 1 0 6072 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_61
timestamp 1666464484
transform 1 0 6716 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_68
timestamp 1666464484
transform 1 0 7360 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_76
timestamp 1666464484
transform 1 0 8096 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1666464484
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_94
timestamp 1666464484
transform 1 0 9752 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_102
timestamp 1666464484
transform 1 0 10488 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_125
timestamp 1666464484
transform 1 0 12604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_137
timestamp 1666464484
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_152
timestamp 1666464484
transform 1 0 15088 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_167
timestamp 1666464484
transform 1 0 16468 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_187
timestamp 1666464484
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1666464484
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_215
timestamp 1666464484
transform 1 0 20884 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_227
timestamp 1666464484
transform 1 0 21988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_239
timestamp 1666464484
transform 1 0 23092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1666464484
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_260
timestamp 1666464484
transform 1 0 25024 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_272
timestamp 1666464484
transform 1 0 26128 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_278
timestamp 1666464484
transform 1 0 26680 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_286
timestamp 1666464484
transform 1 0 27416 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_294
timestamp 1666464484
transform 1 0 28152 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1666464484
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_309
timestamp 1666464484
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_318
timestamp 1666464484
transform 1 0 30360 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_325
timestamp 1666464484
transform 1 0 31004 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_337
timestamp 1666464484
transform 1 0 32108 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_356
timestamp 1666464484
transform 1 0 33856 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1666464484
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_371
timestamp 1666464484
transform 1 0 35236 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_384
timestamp 1666464484
transform 1 0 36432 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_395
timestamp 1666464484
transform 1 0 37444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_402
timestamp 1666464484
transform 1 0 38088 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_406
timestamp 1666464484
transform 1 0 38456 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_15
timestamp 1666464484
transform 1 0 2484 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_43
timestamp 1666464484
transform 1 0 5060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1666464484
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_71
timestamp 1666464484
transform 1 0 7636 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_84
timestamp 1666464484
transform 1 0 8832 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_92
timestamp 1666464484
transform 1 0 9568 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_96
timestamp 1666464484
transform 1 0 9936 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1666464484
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_120
timestamp 1666464484
transform 1 0 12144 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_128
timestamp 1666464484
transform 1 0 12880 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666464484
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666464484
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666464484
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_177
timestamp 1666464484
transform 1 0 17388 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_185
timestamp 1666464484
transform 1 0 18124 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_190
timestamp 1666464484
transform 1 0 18584 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_200
timestamp 1666464484
transform 1 0 19504 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_204
timestamp 1666464484
transform 1 0 19872 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_211
timestamp 1666464484
transform 1 0 20516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666464484
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_237
timestamp 1666464484
transform 1 0 22908 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_265
timestamp 1666464484
transform 1 0 25484 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1666464484
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1666464484
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_295
timestamp 1666464484
transform 1 0 28244 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_307
timestamp 1666464484
transform 1 0 29348 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_324
timestamp 1666464484
transform 1 0 30912 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1666464484
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_361
timestamp 1666464484
transform 1 0 34316 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_369
timestamp 1666464484
transform 1 0 35052 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_378
timestamp 1666464484
transform 1 0 35880 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1666464484
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1666464484
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1666464484
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1666464484
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1666464484
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666464484
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_38
timestamp 1666464484
transform 1 0 4600 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_50
timestamp 1666464484
transform 1 0 5704 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1666464484
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_66
timestamp 1666464484
transform 1 0 7176 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_76
timestamp 1666464484
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666464484
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666464484
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_121
timestamp 1666464484
transform 1 0 12236 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1666464484
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_148
timestamp 1666464484
transform 1 0 14720 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_160
timestamp 1666464484
transform 1 0 15824 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_172
timestamp 1666464484
transform 1 0 16928 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_184
timestamp 1666464484
transform 1 0 18032 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_207
timestamp 1666464484
transform 1 0 20148 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_218
timestamp 1666464484
transform 1 0 21160 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_230
timestamp 1666464484
transform 1 0 22264 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_238
timestamp 1666464484
transform 1 0 23000 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 1666464484
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_271
timestamp 1666464484
transform 1 0 26036 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_275
timestamp 1666464484
transform 1 0 26404 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_296
timestamp 1666464484
transform 1 0 28336 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1666464484
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_321
timestamp 1666464484
transform 1 0 30636 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_347
timestamp 1666464484
transform 1 0 33028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_359
timestamp 1666464484
transform 1 0 34132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1666464484
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_365
timestamp 1666464484
transform 1 0 34684 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_386
timestamp 1666464484
transform 1 0 36616 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_398
timestamp 1666464484
transform 1 0 37720 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_406
timestamp 1666464484
transform 1 0 38456 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1666464484
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1666464484
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1666464484
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1666464484
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1666464484
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666464484
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666464484
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666464484
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666464484
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666464484
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_125
timestamp 1666464484
transform 1 0 12604 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_147
timestamp 1666464484
transform 1 0 14628 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_159
timestamp 1666464484
transform 1 0 15732 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666464484
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1666464484
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_193
timestamp 1666464484
transform 1 0 18860 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_201
timestamp 1666464484
transform 1 0 19596 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_205
timestamp 1666464484
transform 1 0 19964 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_212
timestamp 1666464484
transform 1 0 20608 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_231
timestamp 1666464484
transform 1 0 22356 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_238
timestamp 1666464484
transform 1 0 23000 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_262
timestamp 1666464484
transform 1 0 25208 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1666464484
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1666464484
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_292
timestamp 1666464484
transform 1 0 27968 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_304
timestamp 1666464484
transform 1 0 29072 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_316
timestamp 1666464484
transform 1 0 30176 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_328
timestamp 1666464484
transform 1 0 31280 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1666464484
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1666464484
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_374
timestamp 1666464484
transform 1 0 35512 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_383
timestamp 1666464484
transform 1 0 36340 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1666464484
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1666464484
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1666464484
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1666464484
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1666464484
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1666464484
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1666464484
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666464484
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1666464484
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666464484
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1666464484
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1666464484
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1666464484
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666464484
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_153
timestamp 1666464484
transform 1 0 15180 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_172
timestamp 1666464484
transform 1 0 16928 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_184
timestamp 1666464484
transform 1 0 18032 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1666464484
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_221
timestamp 1666464484
transform 1 0 21436 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_230
timestamp 1666464484
transform 1 0 22264 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1666464484
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1666464484
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_277
timestamp 1666464484
transform 1 0 26588 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_283
timestamp 1666464484
transform 1 0 27140 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_290
timestamp 1666464484
transform 1 0 27784 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_302
timestamp 1666464484
transform 1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_309
timestamp 1666464484
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_313
timestamp 1666464484
transform 1 0 29900 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_330
timestamp 1666464484
transform 1 0 31464 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_342
timestamp 1666464484
transform 1 0 32568 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_354
timestamp 1666464484
transform 1 0 33672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1666464484
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1666464484
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1666464484
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1666464484
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1666464484
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666464484
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1666464484
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1666464484
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_69
timestamp 1666464484
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_90
timestamp 1666464484
transform 1 0 9384 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_97
timestamp 1666464484
transform 1 0 10028 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_104
timestamp 1666464484
transform 1 0 10672 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_124
timestamp 1666464484
transform 1 0 12512 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_133
timestamp 1666464484
transform 1 0 13340 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_145
timestamp 1666464484
transform 1 0 14444 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_157
timestamp 1666464484
transform 1 0 15548 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_165
timestamp 1666464484
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_177
timestamp 1666464484
transform 1 0 17388 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_189
timestamp 1666464484
transform 1 0 18492 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_201
timestamp 1666464484
transform 1 0 19596 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_213
timestamp 1666464484
transform 1 0 20700 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1666464484
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_231
timestamp 1666464484
transform 1 0 22356 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_238
timestamp 1666464484
transform 1 0 23000 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1666464484
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1666464484
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1666464484
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_287
timestamp 1666464484
transform 1 0 27508 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_307
timestamp 1666464484
transform 1 0 29348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_331
timestamp 1666464484
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1666464484
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1666464484
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_345
timestamp 1666464484
transform 1 0 32844 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_357
timestamp 1666464484
transform 1 0 33948 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_369
timestamp 1666464484
transform 1 0 35052 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_381
timestamp 1666464484
transform 1 0 36156 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1666464484
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1666464484
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1666464484
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_15
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1666464484
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_35
timestamp 1666464484
transform 1 0 4324 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_41
timestamp 1666464484
transform 1 0 4876 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_47
timestamp 1666464484
transform 1 0 5428 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_59
timestamp 1666464484
transform 1 0 6532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_67
timestamp 1666464484
transform 1 0 7268 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_74
timestamp 1666464484
transform 1 0 7912 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1666464484
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_95
timestamp 1666464484
transform 1 0 9844 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_99
timestamp 1666464484
transform 1 0 10212 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_107
timestamp 1666464484
transform 1 0 10948 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_118
timestamp 1666464484
transform 1 0 11960 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_127
timestamp 1666464484
transform 1 0 12788 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1666464484
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_153
timestamp 1666464484
transform 1 0 15180 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_157
timestamp 1666464484
transform 1 0 15548 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_178
timestamp 1666464484
transform 1 0 17480 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_188
timestamp 1666464484
transform 1 0 18400 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_202
timestamp 1666464484
transform 1 0 19688 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_211
timestamp 1666464484
transform 1 0 20516 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_223
timestamp 1666464484
transform 1 0 21620 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_235
timestamp 1666464484
transform 1 0 22724 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1666464484
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1666464484
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_277
timestamp 1666464484
transform 1 0 26588 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1666464484
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1666464484
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_309
timestamp 1666464484
transform 1 0 29532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_317
timestamp 1666464484
transform 1 0 30268 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_336
timestamp 1666464484
transform 1 0 32016 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_346
timestamp 1666464484
transform 1 0 32936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_358
timestamp 1666464484
transform 1 0 34040 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1666464484
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1666464484
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1666464484
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1666464484
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_11
timestamp 1666464484
transform 1 0 2116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_17
timestamp 1666464484
transform 1 0 2668 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_40
timestamp 1666464484
transform 1 0 4784 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1666464484
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666464484
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_81
timestamp 1666464484
transform 1 0 8556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_91
timestamp 1666464484
transform 1 0 9476 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_99
timestamp 1666464484
transform 1 0 10212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_106
timestamp 1666464484
transform 1 0 10856 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1666464484
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1666464484
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_149
timestamp 1666464484
transform 1 0 14812 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1666464484
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_190
timestamp 1666464484
transform 1 0 18584 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_202
timestamp 1666464484
transform 1 0 19688 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_214
timestamp 1666464484
transform 1 0 20792 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1666464484
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_237
timestamp 1666464484
transform 1 0 22908 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_257
timestamp 1666464484
transform 1 0 24748 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_269
timestamp 1666464484
transform 1 0 25852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1666464484
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp 1666464484
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_319
timestamp 1666464484
transform 1 0 30452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1666464484
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1666464484
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1666464484
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1666464484
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1666464484
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1666464484
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1666464484
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1666464484
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1666464484
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1666464484
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_11
timestamp 1666464484
transform 1 0 2116 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_25
timestamp 1666464484
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_39
timestamp 1666464484
transform 1 0 4692 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_47
timestamp 1666464484
transform 1 0 5428 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_59
timestamp 1666464484
transform 1 0 6532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_71
timestamp 1666464484
transform 1 0 7636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666464484
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_93
timestamp 1666464484
transform 1 0 9660 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_101
timestamp 1666464484
transform 1 0 10396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_113
timestamp 1666464484
transform 1 0 11500 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_127
timestamp 1666464484
transform 1 0 12788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1666464484
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_152
timestamp 1666464484
transform 1 0 15088 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_164
timestamp 1666464484
transform 1 0 16192 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_185
timestamp 1666464484
transform 1 0 18124 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 1666464484
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_205
timestamp 1666464484
transform 1 0 19964 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_213
timestamp 1666464484
transform 1 0 20700 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_219
timestamp 1666464484
transform 1 0 21252 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_223
timestamp 1666464484
transform 1 0 21620 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_227
timestamp 1666464484
transform 1 0 21988 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_236
timestamp 1666464484
transform 1 0 22816 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_240
timestamp 1666464484
transform 1 0 23184 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_247
timestamp 1666464484
transform 1 0 23828 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1666464484
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_272
timestamp 1666464484
transform 1 0 26128 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_284
timestamp 1666464484
transform 1 0 27232 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_296
timestamp 1666464484
transform 1 0 28336 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1666464484
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_321
timestamp 1666464484
transform 1 0 30636 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_327
timestamp 1666464484
transform 1 0 31188 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_334
timestamp 1666464484
transform 1 0 31832 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_338
timestamp 1666464484
transform 1 0 32200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_348
timestamp 1666464484
transform 1 0 33120 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_358
timestamp 1666464484
transform 1 0 34040 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1666464484
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1666464484
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1666464484
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1666464484
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_19
timestamp 1666464484
transform 1 0 2852 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_35
timestamp 1666464484
transform 1 0 4324 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_43
timestamp 1666464484
transform 1 0 5060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666464484
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1666464484
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1666464484
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1666464484
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1666464484
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1666464484
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_126
timestamp 1666464484
transform 1 0 12696 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_146
timestamp 1666464484
transform 1 0 14536 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_158
timestamp 1666464484
transform 1 0 15640 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1666464484
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_187
timestamp 1666464484
transform 1 0 18308 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_195
timestamp 1666464484
transform 1 0 19044 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_203
timestamp 1666464484
transform 1 0 19780 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_215
timestamp 1666464484
transform 1 0 20884 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1666464484
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_233
timestamp 1666464484
transform 1 0 22540 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_245
timestamp 1666464484
transform 1 0 23644 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_253
timestamp 1666464484
transform 1 0 24380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_262
timestamp 1666464484
transform 1 0 25208 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_274
timestamp 1666464484
transform 1 0 26312 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_287
timestamp 1666464484
transform 1 0 27508 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_296
timestamp 1666464484
transform 1 0 28336 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_308
timestamp 1666464484
transform 1 0 29440 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_320
timestamp 1666464484
transform 1 0 30544 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_328
timestamp 1666464484
transform 1 0 31280 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1666464484
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_337
timestamp 1666464484
transform 1 0 32108 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_341
timestamp 1666464484
transform 1 0 32476 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_355
timestamp 1666464484
transform 1 0 33764 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_367
timestamp 1666464484
transform 1 0 34868 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_379
timestamp 1666464484
transform 1 0 35972 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1666464484
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1666464484
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1666464484
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666464484
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_33
timestamp 1666464484
transform 1 0 4140 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_38
timestamp 1666464484
transform 1 0 4600 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_50
timestamp 1666464484
transform 1 0 5704 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_62
timestamp 1666464484
transform 1 0 6808 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_72
timestamp 1666464484
transform 1 0 7728 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1666464484
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1666464484
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1666464484
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1666464484
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666464484
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_150
timestamp 1666464484
transform 1 0 14904 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_158
timestamp 1666464484
transform 1 0 15640 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_180
timestamp 1666464484
transform 1 0 17664 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_190
timestamp 1666464484
transform 1 0 18584 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_204
timestamp 1666464484
transform 1 0 19872 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_216
timestamp 1666464484
transform 1 0 20976 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_228
timestamp 1666464484
transform 1 0 22080 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_240
timestamp 1666464484
transform 1 0 23184 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_258
timestamp 1666464484
transform 1 0 24840 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_262
timestamp 1666464484
transform 1 0 25208 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_266
timestamp 1666464484
transform 1 0 25576 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_278
timestamp 1666464484
transform 1 0 26680 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_290
timestamp 1666464484
transform 1 0 27784 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_300
timestamp 1666464484
transform 1 0 28704 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1666464484
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_321
timestamp 1666464484
transform 1 0 30636 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_332
timestamp 1666464484
transform 1 0 31648 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_353
timestamp 1666464484
transform 1 0 33580 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1666464484
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1666464484
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1666464484
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1666464484
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1666464484
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666464484
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1666464484
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_39
timestamp 1666464484
transform 1 0 4692 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_48
timestamp 1666464484
transform 1 0 5520 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_69
timestamp 1666464484
transform 1 0 7452 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_74
timestamp 1666464484
transform 1 0 7912 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_86
timestamp 1666464484
transform 1 0 9016 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_95
timestamp 1666464484
transform 1 0 9844 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_107
timestamp 1666464484
transform 1 0 10948 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1666464484
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1666464484
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1666464484
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_149
timestamp 1666464484
transform 1 0 14812 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_157
timestamp 1666464484
transform 1 0 15548 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1666464484
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_177
timestamp 1666464484
transform 1 0 17388 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_189
timestamp 1666464484
transform 1 0 18492 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_201
timestamp 1666464484
transform 1 0 19596 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_213
timestamp 1666464484
transform 1 0 20700 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1666464484
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_234
timestamp 1666464484
transform 1 0 22632 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_246
timestamp 1666464484
transform 1 0 23736 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_252
timestamp 1666464484
transform 1 0 24288 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_258
timestamp 1666464484
transform 1 0 24840 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_270
timestamp 1666464484
transform 1 0 25944 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1666464484
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_289
timestamp 1666464484
transform 1 0 27692 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_300
timestamp 1666464484
transform 1 0 28704 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_310
timestamp 1666464484
transform 1 0 29624 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_322
timestamp 1666464484
transform 1 0 30728 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_326
timestamp 1666464484
transform 1 0 31096 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_334
timestamp 1666464484
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1666464484
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_342
timestamp 1666464484
transform 1 0 32568 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_369
timestamp 1666464484
transform 1 0 35052 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_381
timestamp 1666464484
transform 1 0 36156 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_389
timestamp 1666464484
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1666464484
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1666464484
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1666464484
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1666464484
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_41
timestamp 1666464484
transform 1 0 4876 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_47
timestamp 1666464484
transform 1 0 5428 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_55
timestamp 1666464484
transform 1 0 6164 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_67
timestamp 1666464484
transform 1 0 7268 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_79
timestamp 1666464484
transform 1 0 8372 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666464484
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_96
timestamp 1666464484
transform 1 0 9936 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_107
timestamp 1666464484
transform 1 0 10948 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_119
timestamp 1666464484
transform 1 0 12052 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_131
timestamp 1666464484
transform 1 0 13156 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666464484
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_152
timestamp 1666464484
transform 1 0 15088 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_164
timestamp 1666464484
transform 1 0 16192 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_176
timestamp 1666464484
transform 1 0 17296 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_188
timestamp 1666464484
transform 1 0 18400 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1666464484
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_207
timestamp 1666464484
transform 1 0 20148 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_219
timestamp 1666464484
transform 1 0 21252 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_231
timestamp 1666464484
transform 1 0 22356 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_243
timestamp 1666464484
transform 1 0 23460 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1666464484
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_260
timestamp 1666464484
transform 1 0 25024 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_272
timestamp 1666464484
transform 1 0 26128 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_284
timestamp 1666464484
transform 1 0 27232 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_292
timestamp 1666464484
transform 1 0 27968 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_302
timestamp 1666464484
transform 1 0 28888 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1666464484
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_316
timestamp 1666464484
transform 1 0 30176 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_328
timestamp 1666464484
transform 1 0 31280 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_340
timestamp 1666464484
transform 1 0 32384 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_361
timestamp 1666464484
transform 1 0 34316 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1666464484
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1666464484
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1666464484
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1666464484
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_31
timestamp 1666464484
transform 1 0 3956 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1666464484
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_66
timestamp 1666464484
transform 1 0 7176 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_74
timestamp 1666464484
transform 1 0 7912 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_81
timestamp 1666464484
transform 1 0 8556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_104
timestamp 1666464484
transform 1 0 10672 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1666464484
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_137
timestamp 1666464484
transform 1 0 13708 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_146
timestamp 1666464484
transform 1 0 14536 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_158
timestamp 1666464484
transform 1 0 15640 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1666464484
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_181
timestamp 1666464484
transform 1 0 17756 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_189
timestamp 1666464484
transform 1 0 18492 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_199
timestamp 1666464484
transform 1 0 19412 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_214
timestamp 1666464484
transform 1 0 20792 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1666464484
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_231
timestamp 1666464484
transform 1 0 22356 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_238
timestamp 1666464484
transform 1 0 23000 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_250
timestamp 1666464484
transform 1 0 24104 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_262
timestamp 1666464484
transform 1 0 25208 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_270
timestamp 1666464484
transform 1 0 25944 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1666464484
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_287
timestamp 1666464484
transform 1 0 27508 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_295
timestamp 1666464484
transform 1 0 28244 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_308
timestamp 1666464484
transform 1 0 29440 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_320
timestamp 1666464484
transform 1 0 30544 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1666464484
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1666464484
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1666464484
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1666464484
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1666464484
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1666464484
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1666464484
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1666464484
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1666464484
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1666464484
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666464484
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_37
timestamp 1666464484
transform 1 0 4508 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_54
timestamp 1666464484
transform 1 0 6072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_65
timestamp 1666464484
transform 1 0 7084 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_72
timestamp 1666464484
transform 1 0 7728 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_76
timestamp 1666464484
transform 1 0 8096 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1666464484
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_91
timestamp 1666464484
transform 1 0 9476 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_117
timestamp 1666464484
transform 1 0 11868 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_129
timestamp 1666464484
transform 1 0 12972 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1666464484
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_160
timestamp 1666464484
transform 1 0 15824 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_172
timestamp 1666464484
transform 1 0 16928 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_178
timestamp 1666464484
transform 1 0 17480 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_184
timestamp 1666464484
transform 1 0 18032 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp 1666464484
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_206
timestamp 1666464484
transform 1 0 20056 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_216
timestamp 1666464484
transform 1 0 20976 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_223
timestamp 1666464484
transform 1 0 21620 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_235
timestamp 1666464484
transform 1 0 22724 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1666464484
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_260
timestamp 1666464484
transform 1 0 25024 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_275
timestamp 1666464484
transform 1 0 26404 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_287
timestamp 1666464484
transform 1 0 27508 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_299
timestamp 1666464484
transform 1 0 28612 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1666464484
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1666464484
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_315
timestamp 1666464484
transform 1 0 30084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_327
timestamp 1666464484
transform 1 0 31188 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_335
timestamp 1666464484
transform 1 0 31924 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_342
timestamp 1666464484
transform 1 0 32568 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_350
timestamp 1666464484
transform 1 0 33304 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 1666464484
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1666464484
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1666464484
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1666464484
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1666464484
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_39
timestamp 1666464484
transform 1 0 4692 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_48
timestamp 1666464484
transform 1 0 5520 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_63
timestamp 1666464484
transform 1 0 6900 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_75
timestamp 1666464484
transform 1 0 8004 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_86
timestamp 1666464484
transform 1 0 9016 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_103
timestamp 1666464484
transform 1 0 10580 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1666464484
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_125
timestamp 1666464484
transform 1 0 12604 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_148
timestamp 1666464484
transform 1 0 14720 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_155
timestamp 1666464484
transform 1 0 15364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1666464484
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_173
timestamp 1666464484
transform 1 0 17020 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_177
timestamp 1666464484
transform 1 0 17388 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_202
timestamp 1666464484
transform 1 0 19688 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1666464484
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1666464484
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_249
timestamp 1666464484
transform 1 0 24012 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_255
timestamp 1666464484
transform 1 0 24564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_267
timestamp 1666464484
transform 1 0 25668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1666464484
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_293
timestamp 1666464484
transform 1 0 28060 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_298
timestamp 1666464484
transform 1 0 28520 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_302
timestamp 1666464484
transform 1 0 28888 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_315
timestamp 1666464484
transform 1 0 30084 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_319
timestamp 1666464484
transform 1 0 30452 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_323
timestamp 1666464484
transform 1 0 30820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1666464484
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_337
timestamp 1666464484
transform 1 0 32108 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_347
timestamp 1666464484
transform 1 0 33028 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_357
timestamp 1666464484
transform 1 0 33948 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_369
timestamp 1666464484
transform 1 0 35052 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_381
timestamp 1666464484
transform 1 0 36156 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_389
timestamp 1666464484
transform 1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1666464484
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1666464484
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1666464484
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666464484
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_54
timestamp 1666464484
transform 1 0 6072 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_66
timestamp 1666464484
transform 1 0 7176 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_78
timestamp 1666464484
transform 1 0 8280 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_98
timestamp 1666464484
transform 1 0 10120 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_116
timestamp 1666464484
transform 1 0 11776 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_128
timestamp 1666464484
transform 1 0 12880 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_148
timestamp 1666464484
transform 1 0 14720 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_160
timestamp 1666464484
transform 1 0 15824 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_172
timestamp 1666464484
transform 1 0 16928 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_180
timestamp 1666464484
transform 1 0 17664 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1666464484
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1666464484
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_222
timestamp 1666464484
transform 1 0 21528 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_234
timestamp 1666464484
transform 1 0 22632 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_246
timestamp 1666464484
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1666464484
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1666464484
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_289
timestamp 1666464484
transform 1 0 27692 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_297
timestamp 1666464484
transform 1 0 28428 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1666464484
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1666464484
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_318
timestamp 1666464484
transform 1 0 30360 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_329
timestamp 1666464484
transform 1 0 31372 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_341
timestamp 1666464484
transform 1 0 32476 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_353
timestamp 1666464484
transform 1 0 33580 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_358
timestamp 1666464484
transform 1 0 34040 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_365
timestamp 1666464484
transform 1 0 34684 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_374
timestamp 1666464484
transform 1 0 35512 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_386
timestamp 1666464484
transform 1 0 36616 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_398
timestamp 1666464484
transform 1 0 37720 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_406
timestamp 1666464484
transform 1 0 38456 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1666464484
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1666464484
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_39
timestamp 1666464484
transform 1 0 4692 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_49
timestamp 1666464484
transform 1 0 5612 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1666464484
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666464484
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1666464484
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1666464484
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1666464484
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1666464484
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_146
timestamp 1666464484
transform 1 0 14536 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_155
timestamp 1666464484
transform 1 0 15364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1666464484
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_173
timestamp 1666464484
transform 1 0 17020 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_177
timestamp 1666464484
transform 1 0 17388 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_189
timestamp 1666464484
transform 1 0 18492 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_195
timestamp 1666464484
transform 1 0 19044 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_213
timestamp 1666464484
transform 1 0 20700 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_221
timestamp 1666464484
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_235
timestamp 1666464484
transform 1 0 22724 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_246
timestamp 1666464484
transform 1 0 23736 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_258
timestamp 1666464484
transform 1 0 24840 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_270
timestamp 1666464484
transform 1 0 25944 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1666464484
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1666464484
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_305
timestamp 1666464484
transform 1 0 29164 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_313
timestamp 1666464484
transform 1 0 29900 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_322
timestamp 1666464484
transform 1 0 30728 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_334
timestamp 1666464484
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1666464484
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_349
timestamp 1666464484
transform 1 0 33212 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_369
timestamp 1666464484
transform 1 0 35052 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_381
timestamp 1666464484
transform 1 0 36156 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_389
timestamp 1666464484
transform 1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1666464484
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1666464484
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1666464484
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666464484
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666464484
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666464484
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666464484
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666464484
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1666464484
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1666464484
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1666464484
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1666464484
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1666464484
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1666464484
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1666464484
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1666464484
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1666464484
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_152
timestamp 1666464484
transform 1 0 15088 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_164
timestamp 1666464484
transform 1 0 16192 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_176
timestamp 1666464484
transform 1 0 17296 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_182
timestamp 1666464484
transform 1 0 17848 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1666464484
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1666464484
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1666464484
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1666464484
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_233
timestamp 1666464484
transform 1 0 22540 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1666464484
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1666464484
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1666464484
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1666464484
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_277
timestamp 1666464484
transform 1 0 26588 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_285
timestamp 1666464484
transform 1 0 27324 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_291
timestamp 1666464484
transform 1 0 27876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_303
timestamp 1666464484
transform 1 0 28980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1666464484
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1666464484
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1666464484
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1666464484
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_345
timestamp 1666464484
transform 1 0 32844 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_351
timestamp 1666464484
transform 1 0 33396 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_355
timestamp 1666464484
transform 1 0 33764 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_362
timestamp 1666464484
transform 1 0 34408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_365
timestamp 1666464484
transform 1 0 34684 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_376
timestamp 1666464484
transform 1 0 35696 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_388
timestamp 1666464484
transform 1 0 36800 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_400
timestamp 1666464484
transform 1 0 37904 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_406
timestamp 1666464484
transform 1 0 38456 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666464484
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666464484
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1666464484
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1666464484
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1666464484
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666464484
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1666464484
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1666464484
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1666464484
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666464484
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666464484
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1666464484
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1666464484
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1666464484
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1666464484
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1666464484
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666464484
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_169
timestamp 1666464484
transform 1 0 16652 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_175
timestamp 1666464484
transform 1 0 17204 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_183
timestamp 1666464484
transform 1 0 17940 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_192
timestamp 1666464484
transform 1 0 18768 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_204
timestamp 1666464484
transform 1 0 19872 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_212
timestamp 1666464484
transform 1 0 20608 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_218
timestamp 1666464484
transform 1 0 21160 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_225
timestamp 1666464484
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_233
timestamp 1666464484
transform 1 0 22540 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_258
timestamp 1666464484
transform 1 0 24840 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_270
timestamp 1666464484
transform 1 0 25944 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1666464484
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1666464484
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_288
timestamp 1666464484
transform 1 0 27600 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_297
timestamp 1666464484
transform 1 0 28428 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_304
timestamp 1666464484
transform 1 0 29072 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_316
timestamp 1666464484
transform 1 0 30176 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_328
timestamp 1666464484
transform 1 0 31280 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1666464484
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_349
timestamp 1666464484
transform 1 0 33212 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_355
timestamp 1666464484
transform 1 0 33764 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_360
timestamp 1666464484
transform 1 0 34224 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_367
timestamp 1666464484
transform 1 0 34868 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_374
timestamp 1666464484
transform 1 0 35512 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_386
timestamp 1666464484
transform 1 0 36616 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1666464484
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1666464484
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1666464484
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1666464484
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1666464484
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1666464484
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1666464484
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1666464484
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666464484
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1666464484
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666464484
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1666464484
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1666464484
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1666464484
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1666464484
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1666464484
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1666464484
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1666464484
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1666464484
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_165
timestamp 1666464484
transform 1 0 16284 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_174
timestamp 1666464484
transform 1 0 17112 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_187
timestamp 1666464484
transform 1 0 18308 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1666464484
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1666464484
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1666464484
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1666464484
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_233
timestamp 1666464484
transform 1 0 22540 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1666464484
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1666464484
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1666464484
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_264
timestamp 1666464484
transform 1 0 25392 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_275
timestamp 1666464484
transform 1 0 26404 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_279
timestamp 1666464484
transform 1 0 26772 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_288
timestamp 1666464484
transform 1 0 27600 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_292
timestamp 1666464484
transform 1 0 27968 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1666464484
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1666464484
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1666464484
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1666464484
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1666464484
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1666464484
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1666464484
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1666464484
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1666464484
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1666464484
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1666464484
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1666464484
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1666464484
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1666464484
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1666464484
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1666464484
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1666464484
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1666464484
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1666464484
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1666464484
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1666464484
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1666464484
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1666464484
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1666464484
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1666464484
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1666464484
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1666464484
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 1666464484
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_169
timestamp 1666464484
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_181
timestamp 1666464484
transform 1 0 17756 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_201
timestamp 1666464484
transform 1 0 19596 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_213
timestamp 1666464484
transform 1 0 20700 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 1666464484
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1666464484
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1666464484
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_249
timestamp 1666464484
transform 1 0 24012 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_257
timestamp 1666464484
transform 1 0 24748 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_265
timestamp 1666464484
transform 1 0 25484 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_273
timestamp 1666464484
transform 1 0 26220 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1666464484
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_281
timestamp 1666464484
transform 1 0 26956 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_306
timestamp 1666464484
transform 1 0 29256 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1666464484
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_57_337
timestamp 1666464484
transform 1 0 32108 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_346
timestamp 1666464484
transform 1 0 32936 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_358
timestamp 1666464484
transform 1 0 34040 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_370
timestamp 1666464484
transform 1 0 35144 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_382
timestamp 1666464484
transform 1 0 36248 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_390
timestamp 1666464484
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1666464484
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1666464484
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1666464484
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1666464484
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1666464484
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1666464484
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1666464484
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1666464484
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1666464484
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1666464484
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1666464484
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1666464484
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1666464484
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1666464484
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1666464484
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1666464484
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1666464484
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1666464484
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1666464484
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_165
timestamp 1666464484
transform 1 0 16284 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_179
timestamp 1666464484
transform 1 0 17572 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1666464484
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1666464484
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_209
timestamp 1666464484
transform 1 0 20332 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_230
timestamp 1666464484
transform 1 0 22264 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_242
timestamp 1666464484
transform 1 0 23368 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1666464484
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_253
timestamp 1666464484
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_261
timestamp 1666464484
transform 1 0 25116 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_280
timestamp 1666464484
transform 1 0 26864 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_292
timestamp 1666464484
transform 1 0 27968 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_304
timestamp 1666464484
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1666464484
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1666464484
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_333
timestamp 1666464484
transform 1 0 31740 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_348
timestamp 1666464484
transform 1 0 33120 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1666464484
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1666464484
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1666464484
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1666464484
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1666464484
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1666464484
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1666464484
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1666464484
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1666464484
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1666464484
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1666464484
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1666464484
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1666464484
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1666464484
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1666464484
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1666464484
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1666464484
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1666464484
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1666464484
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1666464484
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1666464484
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1666464484
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1666464484
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_169
timestamp 1666464484
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_194
timestamp 1666464484
transform 1 0 18952 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_202
timestamp 1666464484
transform 1 0 19688 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1666464484
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1666464484
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_233
timestamp 1666464484
transform 1 0 22540 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_241
timestamp 1666464484
transform 1 0 23276 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_260
timestamp 1666464484
transform 1 0 25024 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_269
timestamp 1666464484
transform 1 0 25852 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_277
timestamp 1666464484
transform 1 0 26588 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1666464484
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1666464484
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_305
timestamp 1666464484
transform 1 0 29164 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_311
timestamp 1666464484
transform 1 0 29716 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_315
timestamp 1666464484
transform 1 0 30084 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_327
timestamp 1666464484
transform 1 0 31188 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1666464484
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_337
timestamp 1666464484
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_343
timestamp 1666464484
transform 1 0 32660 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_369
timestamp 1666464484
transform 1 0 35052 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_381
timestamp 1666464484
transform 1 0 36156 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_389
timestamp 1666464484
transform 1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1666464484
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1666464484
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1666464484
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1666464484
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1666464484
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1666464484
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1666464484
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1666464484
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1666464484
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1666464484
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1666464484
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1666464484
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1666464484
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1666464484
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1666464484
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1666464484
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1666464484
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1666464484
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1666464484
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1666464484
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_177
timestamp 1666464484
transform 1 0 17388 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1666464484
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_197
timestamp 1666464484
transform 1 0 19228 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_214
timestamp 1666464484
transform 1 0 20792 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_225
timestamp 1666464484
transform 1 0 21804 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_229
timestamp 1666464484
transform 1 0 22172 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_236
timestamp 1666464484
transform 1 0 22816 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1666464484
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1666464484
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 1666464484
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_261
timestamp 1666464484
transform 1 0 25116 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_269
timestamp 1666464484
transform 1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_285
timestamp 1666464484
transform 1 0 27324 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_297
timestamp 1666464484
transform 1 0 28428 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_305
timestamp 1666464484
transform 1 0 29164 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_309
timestamp 1666464484
transform 1 0 29532 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_320
timestamp 1666464484
transform 1 0 30544 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_332
timestamp 1666464484
transform 1 0 31648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_355
timestamp 1666464484
transform 1 0 33764 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1666464484
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_365
timestamp 1666464484
transform 1 0 34684 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_380
timestamp 1666464484
transform 1 0 36064 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_392
timestamp 1666464484
transform 1 0 37168 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_404
timestamp 1666464484
transform 1 0 38272 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1666464484
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1666464484
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1666464484
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1666464484
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1666464484
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1666464484
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1666464484
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1666464484
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1666464484
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1666464484
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1666464484
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1666464484
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1666464484
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1666464484
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_137
timestamp 1666464484
transform 1 0 13708 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_147
timestamp 1666464484
transform 1 0 14628 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_159
timestamp 1666464484
transform 1 0 15732 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1666464484
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1666464484
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_181
timestamp 1666464484
transform 1 0 17756 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_209
timestamp 1666464484
transform 1 0 20332 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_217
timestamp 1666464484
transform 1 0 21068 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1666464484
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1666464484
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_236
timestamp 1666464484
transform 1 0 22816 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_245
timestamp 1666464484
transform 1 0 23644 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_257
timestamp 1666464484
transform 1 0 24748 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_271
timestamp 1666464484
transform 1 0 26036 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1666464484
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1666464484
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_293
timestamp 1666464484
transform 1 0 28060 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_301
timestamp 1666464484
transform 1 0 28796 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_305
timestamp 1666464484
transform 1 0 29164 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_323
timestamp 1666464484
transform 1 0 30820 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_331
timestamp 1666464484
transform 1 0 31556 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1666464484
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_337
timestamp 1666464484
transform 1 0 32108 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_361
timestamp 1666464484
transform 1 0 34316 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_370
timestamp 1666464484
transform 1 0 35144 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_382
timestamp 1666464484
transform 1 0 36248 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1666464484
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1666464484
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1666464484
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1666464484
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1666464484
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1666464484
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1666464484
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1666464484
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1666464484
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1666464484
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1666464484
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1666464484
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1666464484
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1666464484
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1666464484
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1666464484
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1666464484
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1666464484
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 1666464484
transform 1 0 14076 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_154
timestamp 1666464484
transform 1 0 15272 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_166
timestamp 1666464484
transform 1 0 16376 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_184
timestamp 1666464484
transform 1 0 18032 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1666464484
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1666464484
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1666464484
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1666464484
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1666464484
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1666464484
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_253
timestamp 1666464484
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_260
timestamp 1666464484
transform 1 0 25024 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_273
timestamp 1666464484
transform 1 0 26220 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_285
timestamp 1666464484
transform 1 0 27324 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_297
timestamp 1666464484
transform 1 0 28428 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1666464484
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_309
timestamp 1666464484
transform 1 0 29532 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_317
timestamp 1666464484
transform 1 0 30268 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_326
timestamp 1666464484
transform 1 0 31096 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_338
timestamp 1666464484
transform 1 0 32200 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_346
timestamp 1666464484
transform 1 0 32936 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_355
timestamp 1666464484
transform 1 0 33764 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_362
timestamp 1666464484
transform 1 0 34408 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1666464484
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1666464484
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_389
timestamp 1666464484
transform 1 0 36892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_394
timestamp 1666464484
transform 1 0 37352 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_406
timestamp 1666464484
transform 1 0 38456 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1666464484
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1666464484
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1666464484
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1666464484
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1666464484
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1666464484
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1666464484
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1666464484
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1666464484
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1666464484
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1666464484
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1666464484
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1666464484
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1666464484
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_137
timestamp 1666464484
transform 1 0 13708 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_147
timestamp 1666464484
transform 1 0 14628 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_159
timestamp 1666464484
transform 1 0 15732 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1666464484
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1666464484
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_181
timestamp 1666464484
transform 1 0 17756 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_207
timestamp 1666464484
transform 1 0 20148 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_219
timestamp 1666464484
transform 1 0 21252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1666464484
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1666464484
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1666464484
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_249
timestamp 1666464484
transform 1 0 24012 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_257
timestamp 1666464484
transform 1 0 24748 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_266
timestamp 1666464484
transform 1 0 25576 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1666464484
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1666464484
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1666464484
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1666464484
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_305
timestamp 1666464484
transform 1 0 29164 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_313
timestamp 1666464484
transform 1 0 29900 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_318
timestamp 1666464484
transform 1 0 30360 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_330
timestamp 1666464484
transform 1 0 31464 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1666464484
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1666464484
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1666464484
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1666464484
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1666464484
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1666464484
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1666464484
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1666464484
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1666464484
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1666464484
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1666464484
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1666464484
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_41
timestamp 1666464484
transform 1 0 4876 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_48
timestamp 1666464484
transform 1 0 5520 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_57
timestamp 1666464484
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_69
timestamp 1666464484
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1666464484
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1666464484
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_91
timestamp 1666464484
transform 1 0 9476 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_103
timestamp 1666464484
transform 1 0 10580 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1666464484
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_113
timestamp 1666464484
transform 1 0 11500 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_120
timestamp 1666464484
transform 1 0 12144 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_132
timestamp 1666464484
transform 1 0 13248 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_141
timestamp 1666464484
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_149
timestamp 1666464484
transform 1 0 14812 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_156
timestamp 1666464484
transform 1 0 15456 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_169
timestamp 1666464484
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_181
timestamp 1666464484
transform 1 0 17756 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_187
timestamp 1666464484
transform 1 0 18308 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1666464484
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1666464484
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1666464484
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 1666464484
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1666464484
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_231
timestamp 1666464484
transform 1 0 22356 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_243
timestamp 1666464484
transform 1 0 23460 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1666464484
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_253
timestamp 1666464484
transform 1 0 24380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_259
timestamp 1666464484
transform 1 0 24932 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_264
timestamp 1666464484
transform 1 0 25392 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_276
timestamp 1666464484
transform 1 0 26496 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_281
timestamp 1666464484
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_293
timestamp 1666464484
transform 1 0 28060 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_300
timestamp 1666464484
transform 1 0 28704 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1666464484
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1666464484
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_333
timestamp 1666464484
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1666464484
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_343
timestamp 1666464484
transform 1 0 32660 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_355
timestamp 1666464484
transform 1 0 33764 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1666464484
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_365
timestamp 1666464484
transform 1 0 34684 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_372
timestamp 1666464484
transform 1 0 35328 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_384
timestamp 1666464484
transform 1 0 36432 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_393
timestamp 1666464484
transform 1 0 37260 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1666464484
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666464484
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666464484
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666464484
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666464484
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666464484
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666464484
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666464484
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666464484
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666464484
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666464484
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666464484
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666464484
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666464484
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666464484
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666464484
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666464484
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666464484
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666464484
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666464484
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666464484
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666464484
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666464484
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666464484
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666464484
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666464484
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666464484
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666464484
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666464484
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666464484
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666464484
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666464484
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666464484
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666464484
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666464484
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666464484
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666464484
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666464484
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666464484
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666464484
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666464484
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666464484
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666464484
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666464484
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666464484
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666464484
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666464484
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666464484
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666464484
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666464484
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666464484
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666464484
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666464484
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666464484
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666464484
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666464484
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666464484
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666464484
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666464484
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666464484
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666464484
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666464484
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666464484
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666464484
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666464484
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666464484
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666464484
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666464484
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666464484
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666464484
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666464484
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666464484
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666464484
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666464484
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666464484
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666464484
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666464484
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666464484
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666464484
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666464484
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666464484
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666464484
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666464484
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666464484
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666464484
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666464484
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666464484
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666464484
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666464484
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666464484
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666464484
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666464484
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666464484
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666464484
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666464484
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666464484
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666464484
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666464484
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666464484
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666464484
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666464484
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666464484
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666464484
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666464484
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666464484
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666464484
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666464484
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666464484
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666464484
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666464484
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666464484
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666464484
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666464484
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666464484
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666464484
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666464484
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666464484
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666464484
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666464484
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666464484
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666464484
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666464484
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666464484
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666464484
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666464484
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666464484
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666464484
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0465_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1666464484
transform 1 0 2668 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_6  _0467_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7084 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_4  _0468_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10120 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0469_
timestamp 1666464484
transform 1 0 11684 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0470_
timestamp 1666464484
transform 1 0 10396 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0471_
timestamp 1666464484
transform 1 0 10856 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1666464484
transform 1 0 12236 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_6  _0473_
timestamp 1666464484
transform 1 0 23092 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__inv_4  _0474_
timestamp 1666464484
transform 1 0 34684 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _0475_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22356 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _0476_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20056 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0477_
timestamp 1666464484
transform 1 0 20332 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1666464484
transform 1 0 18676 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1666464484
transform 1 0 17112 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0480_
timestamp 1666464484
transform 1 0 36984 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0481_
timestamp 1666464484
transform 1 0 34132 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0482__1
timestamp 1666464484
transform 1 0 12696 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0483_
timestamp 1666464484
transform 1 0 2576 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1666464484
transform 1 0 4692 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1666464484
transform 1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _0486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27232 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0487_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8280 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0488_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0489_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9200 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9108 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_4  _0491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9108 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__mux2_1  _0492_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7820 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0493_
timestamp 1666464484
transform 1 0 9108 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0494_
timestamp 1666464484
transform 1 0 24564 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0495_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11040 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0496_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10304 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0497_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14260 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0498_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22724 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0499_
timestamp 1666464484
transform 1 0 10488 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0500_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_4  _0501_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9936 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _0502_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16836 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0503_
timestamp 1666464484
transform 1 0 18032 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0504_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16468 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1666464484
transform 1 0 14812 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0506_
timestamp 1666464484
transform 1 0 14444 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0507_
timestamp 1666464484
transform 1 0 7360 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _0508_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9016 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0509_
timestamp 1666464484
transform 1 0 12144 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0510_
timestamp 1666464484
transform 1 0 11684 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0511_
timestamp 1666464484
transform 1 0 21528 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0512_
timestamp 1666464484
transform 1 0 6532 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0513_
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1666464484
transform 1 0 7636 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0515_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0516_
timestamp 1666464484
transform 1 0 6440 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0517_
timestamp 1666464484
transform 1 0 19780 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0518_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5244 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0519_
timestamp 1666464484
transform 1 0 18400 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0520_
timestamp 1666464484
transform 1 0 9568 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0521_
timestamp 1666464484
transform 1 0 16836 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0522_
timestamp 1666464484
transform 1 0 9568 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0523_
timestamp 1666464484
transform 1 0 14812 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0524_
timestamp 1666464484
transform 1 0 6992 0 1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0525_
timestamp 1666464484
transform 1 0 14076 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0526_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4140 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _0527_
timestamp 1666464484
transform 1 0 28244 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _0528_
timestamp 1666464484
transform 1 0 13800 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0529_
timestamp 1666464484
transform 1 0 13800 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0530_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14444 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0531_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16928 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _0532_
timestamp 1666464484
transform 1 0 2668 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1666464484
transform 1 0 9660 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0534_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0535_
timestamp 1666464484
transform 1 0 3680 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0536_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2760 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0537_
timestamp 1666464484
transform 1 0 3772 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0538_
timestamp 1666464484
transform 1 0 1656 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0539_
timestamp 1666464484
transform 1 0 2576 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_2  _0540_
timestamp 1666464484
transform 1 0 2484 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _0541_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2576 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0542_
timestamp 1666464484
transform 1 0 2760 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0543_
timestamp 1666464484
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0544_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8004 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0545_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4968 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0546_
timestamp 1666464484
transform 1 0 32292 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0547_
timestamp 1666464484
transform 1 0 33488 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0548_
timestamp 1666464484
transform 1 0 33948 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0549_
timestamp 1666464484
transform 1 0 20056 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0550_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0551_
timestamp 1666464484
transform 1 0 19228 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0552_
timestamp 1666464484
transform 1 0 18768 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0553_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0554_
timestamp 1666464484
transform 1 0 17112 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0555_
timestamp 1666464484
transform 1 0 17572 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0556_
timestamp 1666464484
transform 1 0 21344 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0557_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20424 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0558_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19504 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0559_
timestamp 1666464484
transform 1 0 18400 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_2  _0560_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19964 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_4  _0561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20056 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__a32o_4  _0562_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19136 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _0563_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18308 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0564_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17296 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0565_
timestamp 1666464484
transform 1 0 15916 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a311oi_4  _0566_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19596 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_2  _0567_
timestamp 1666464484
transform 1 0 21988 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0568_
timestamp 1666464484
transform 1 0 21252 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0569_
timestamp 1666464484
transform 1 0 20700 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0570_
timestamp 1666464484
transform 1 0 17940 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_8  _0571_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17756 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_4  _0572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18124 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0573_
timestamp 1666464484
transform 1 0 17388 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0574_
timestamp 1666464484
transform 1 0 17480 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _0575_
timestamp 1666464484
transform 1 0 16560 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0576_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17020 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_4  _0577_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18124 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__o31ai_4  _0578_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19964 0 -1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__o31a_2  _0579_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16836 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_4  _0580_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17388 0 -1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__o311a_4  _0581_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20700 0 1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__and2b_1  _0582_
timestamp 1666464484
transform 1 0 23092 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0583_
timestamp 1666464484
transform 1 0 23184 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0584_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17940 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_2  _0585_
timestamp 1666464484
transform 1 0 19964 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _0586_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18124 0 -1 36992
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0587_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18308 0 -1 35904
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1666464484
transform 1 0 24748 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0589_
timestamp 1666464484
transform 1 0 28796 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0590_
timestamp 1666464484
transform 1 0 27140 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1666464484
transform 1 0 26404 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0592_
timestamp 1666464484
transform 1 0 27968 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0593_
timestamp 1666464484
transform 1 0 23092 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_4  _0594_
timestamp 1666464484
transform 1 0 22816 0 -1 32640
box -38 -48 2062 592
use sky130_fd_sc_hd__a21oi_2  _0595_
timestamp 1666464484
transform 1 0 24840 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_2  _0596_
timestamp 1666464484
transform 1 0 24564 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0597_
timestamp 1666464484
transform 1 0 25392 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0598_
timestamp 1666464484
transform 1 0 25760 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0599_
timestamp 1666464484
transform 1 0 24748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23184 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0601_
timestamp 1666464484
transform 1 0 22264 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_4  _0602_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23460 0 -1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__or3b_1  _0603_
timestamp 1666464484
transform 1 0 21160 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _0604_
timestamp 1666464484
transform 1 0 21988 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _0605_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24932 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _0606_
timestamp 1666464484
transform 1 0 27600 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_4  _0607_
timestamp 1666464484
transform 1 0 25392 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__xnor2_2  _0608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26128 0 1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0609_
timestamp 1666464484
transform 1 0 28888 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0610_
timestamp 1666464484
transform 1 0 31372 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0611_
timestamp 1666464484
transform 1 0 32384 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0612_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32476 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _0613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28060 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _0614_
timestamp 1666464484
transform 1 0 29624 0 -1 33728
box -38 -48 2062 592
use sky130_fd_sc_hd__o21ai_1  _0615_
timestamp 1666464484
transform 1 0 32292 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _0616_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26864 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _0617_
timestamp 1666464484
transform 1 0 27232 0 -1 33728
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0618_
timestamp 1666464484
transform 1 0 29808 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_4  _0619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31832 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _0620_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24932 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0621_
timestamp 1666464484
transform 1 0 25944 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0622_
timestamp 1666464484
transform 1 0 25392 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_1  _0623_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29716 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_4  _0624_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29532 0 -1 35904
box -38 -48 1326 592
use sky130_fd_sc_hd__a21boi_2  _0625_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _0626_
timestamp 1666464484
transform 1 0 32568 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_4  _0627_
timestamp 1666464484
transform 1 0 31004 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0628_
timestamp 1666464484
transform 1 0 33120 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0629_
timestamp 1666464484
transform 1 0 34132 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0630_
timestamp 1666464484
transform 1 0 34868 0 1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1666464484
transform 1 0 35236 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0632_
timestamp 1666464484
transform 1 0 33488 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_4  _0633_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32844 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__xnor2_4  _0634_
timestamp 1666464484
transform 1 0 33028 0 -1 34816
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0635_
timestamp 1666464484
transform 1 0 33764 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_4  _0636_
timestamp 1666464484
transform 1 0 33120 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _0637_
timestamp 1666464484
transform 1 0 34132 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0638_
timestamp 1666464484
transform 1 0 30636 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0639_
timestamp 1666464484
transform 1 0 31188 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0640_
timestamp 1666464484
transform 1 0 30084 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0641_
timestamp 1666464484
transform 1 0 28980 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0642_
timestamp 1666464484
transform 1 0 29716 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0643_
timestamp 1666464484
transform 1 0 33856 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_4  _0644_
timestamp 1666464484
transform 1 0 33764 0 -1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__o211ai_4  _0645_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32752 0 1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__a21o_1  _0646_
timestamp 1666464484
transform 1 0 33396 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0647_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32936 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_2  _0648_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0649_
timestamp 1666464484
transform 1 0 32016 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0650_
timestamp 1666464484
transform 1 0 30544 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0651_
timestamp 1666464484
transform 1 0 30176 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0652_
timestamp 1666464484
transform 1 0 31188 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_4  _0653_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32016 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _0654_
timestamp 1666464484
transform 1 0 29716 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0655_
timestamp 1666464484
transform 1 0 25300 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0656_
timestamp 1666464484
transform 1 0 24564 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1666464484
transform 1 0 23828 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0658_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24380 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0659_
timestamp 1666464484
transform 1 0 24564 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0660_
timestamp 1666464484
transform 1 0 25576 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0661_
timestamp 1666464484
transform 1 0 24288 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0662_
timestamp 1666464484
transform 1 0 24472 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0663_
timestamp 1666464484
transform 1 0 29072 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0664_
timestamp 1666464484
transform 1 0 27600 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0665_
timestamp 1666464484
transform 1 0 34592 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0666_
timestamp 1666464484
transform 1 0 34868 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0667_
timestamp 1666464484
transform 1 0 34868 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0668_
timestamp 1666464484
transform 1 0 30728 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _0669_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28980 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_1  _0670_
timestamp 1666464484
transform 1 0 28704 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0671_
timestamp 1666464484
transform 1 0 29716 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0672_
timestamp 1666464484
transform 1 0 29716 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0673_
timestamp 1666464484
transform 1 0 16744 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0674_
timestamp 1666464484
transform 1 0 19320 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0675_
timestamp 1666464484
transform 1 0 28152 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0676_
timestamp 1666464484
transform 1 0 28060 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _0677_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16376 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _0678_
timestamp 1666464484
transform 1 0 17112 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_4  _0679_
timestamp 1666464484
transform 1 0 16836 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__or2_4  _0680_
timestamp 1666464484
transform 1 0 18308 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0681_
timestamp 1666464484
transform 1 0 35696 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0682_
timestamp 1666464484
transform 1 0 36432 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0683_
timestamp 1666464484
transform 1 0 35604 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0684_
timestamp 1666464484
transform 1 0 36432 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0685_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 33304 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1666464484
transform 1 0 32660 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _0687_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 34592 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _0688_
timestamp 1666464484
transform 1 0 36340 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_2  _0689_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 35696 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0690_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 35604 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0691_
timestamp 1666464484
transform 1 0 35512 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _0692_
timestamp 1666464484
transform 1 0 36156 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0693_
timestamp 1666464484
transform 1 0 34868 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0694_
timestamp 1666464484
transform 1 0 34868 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _0695_
timestamp 1666464484
transform 1 0 34408 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0696_
timestamp 1666464484
transform 1 0 36524 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0697_
timestamp 1666464484
transform 1 0 36248 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _0698_
timestamp 1666464484
transform 1 0 34408 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_2  _0699_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 35788 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _0700_
timestamp 1666464484
transform 1 0 35880 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0701_
timestamp 1666464484
transform 1 0 37352 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0702_
timestamp 1666464484
transform 1 0 37444 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0703_
timestamp 1666464484
transform 1 0 36708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0704_
timestamp 1666464484
transform 1 0 35972 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_2  _0705_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 35880 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0706_
timestamp 1666464484
transform 1 0 35420 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0707_
timestamp 1666464484
transform 1 0 37812 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0708_
timestamp 1666464484
transform 1 0 36800 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0709_
timestamp 1666464484
transform 1 0 32292 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_4  _0710_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32476 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ba_1  _0711_
timestamp 1666464484
transform 1 0 33120 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0712_
timestamp 1666464484
transform 1 0 35788 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 35880 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_4  _0714_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 33120 0 1 17408
box -38 -48 1326 592
use sky130_fd_sc_hd__xor2_2  _0715_
timestamp 1666464484
transform 1 0 32660 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__a22oi_1  _0716_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 34868 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0717_
timestamp 1666464484
transform 1 0 34132 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0718_
timestamp 1666464484
transform 1 0 34868 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0719_
timestamp 1666464484
transform 1 0 33028 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0720_
timestamp 1666464484
transform 1 0 29900 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _0721_
timestamp 1666464484
transform 1 0 32292 0 -1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0722_
timestamp 1666464484
transform 1 0 30728 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_4  _0723_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32476 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__and2_1  _0724_
timestamp 1666464484
transform 1 0 35880 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0725_
timestamp 1666464484
transform 1 0 35236 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0726_
timestamp 1666464484
transform 1 0 34868 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0727_
timestamp 1666464484
transform 1 0 30820 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_4  _0728_
timestamp 1666464484
transform 1 0 16836 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _0729_
timestamp 1666464484
transform 1 0 18124 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_4  _0730_
timestamp 1666464484
transform 1 0 17112 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _0731_
timestamp 1666464484
transform 1 0 17756 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _0732_
timestamp 1666464484
transform 1 0 17204 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0733_
timestamp 1666464484
transform 1 0 18124 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0734_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18124 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0735_
timestamp 1666464484
transform 1 0 18492 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0736_
timestamp 1666464484
transform 1 0 15916 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0737_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0738_
timestamp 1666464484
transform 1 0 18676 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0739_
timestamp 1666464484
transform 1 0 19412 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0740_
timestamp 1666464484
transform 1 0 18768 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0741_
timestamp 1666464484
transform 1 0 19412 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0742_
timestamp 1666464484
transform 1 0 24748 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0743_
timestamp 1666464484
transform 1 0 25852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0744_
timestamp 1666464484
transform 1 0 17296 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0745_
timestamp 1666464484
transform 1 0 16928 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0746_
timestamp 1666464484
transform 1 0 15824 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0747_
timestamp 1666464484
transform 1 0 18308 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1666464484
transform 1 0 19688 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0749_
timestamp 1666464484
transform 1 0 19412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0750_
timestamp 1666464484
transform 1 0 19412 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0751_
timestamp 1666464484
transform 1 0 26772 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0752_
timestamp 1666464484
transform 1 0 28244 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0753_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27508 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _0754_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27600 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_4  _0755_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12512 0 1 22848
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_1  _0756_
timestamp 1666464484
transform 1 0 3220 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0757_
timestamp 1666464484
transform 1 0 2208 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0758_
timestamp 1666464484
transform 1 0 2392 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0759_
timestamp 1666464484
transform 1 0 25760 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0760_
timestamp 1666464484
transform 1 0 28244 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _0761_
timestamp 1666464484
transform 1 0 28152 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0762_
timestamp 1666464484
transform 1 0 27968 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0763_
timestamp 1666464484
transform 1 0 33028 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0764_
timestamp 1666464484
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0765_
timestamp 1666464484
transform 1 0 32384 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0766_
timestamp 1666464484
transform 1 0 18124 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0767_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18952 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0768_
timestamp 1666464484
transform 1 0 25208 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0769_
timestamp 1666464484
transform 1 0 20424 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0770_
timestamp 1666464484
transform 1 0 20516 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0771_
timestamp 1666464484
transform 1 0 24748 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0772_
timestamp 1666464484
transform 1 0 28428 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0773_
timestamp 1666464484
transform 1 0 28244 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_2  _0774_
timestamp 1666464484
transform 1 0 27600 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0775_
timestamp 1666464484
transform 1 0 13248 0 -1 27200
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1666464484
transform 1 0 7452 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _0777_
timestamp 1666464484
transform 1 0 4048 0 -1 29376
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_2  _0778_
timestamp 1666464484
transform 1 0 4048 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0779_
timestamp 1666464484
transform 1 0 5060 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0780_
timestamp 1666464484
transform 1 0 23460 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0781_
timestamp 1666464484
transform 1 0 23368 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0782_
timestamp 1666464484
transform 1 0 24564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0783_
timestamp 1666464484
transform 1 0 22448 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0784_
timestamp 1666464484
transform 1 0 34316 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _0785_
timestamp 1666464484
transform 1 0 30544 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0786_
timestamp 1666464484
transform 1 0 26128 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0787_
timestamp 1666464484
transform 1 0 20056 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0788_
timestamp 1666464484
transform 1 0 26220 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0789_
timestamp 1666464484
transform 1 0 14536 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0790_
timestamp 1666464484
transform 1 0 28152 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0791_
timestamp 1666464484
transform 1 0 18216 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _0792_
timestamp 1666464484
transform 1 0 18768 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _0793_
timestamp 1666464484
transform 1 0 17940 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0794_
timestamp 1666464484
transform 1 0 21988 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _0795_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21988 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0796_
timestamp 1666464484
transform 1 0 15088 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_4  _0797_
timestamp 1666464484
transform 1 0 14260 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1666464484
transform 1 0 10948 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _0799_
timestamp 1666464484
transform 1 0 9844 0 1 29376
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_2  _0800_
timestamp 1666464484
transform 1 0 8004 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0801_
timestamp 1666464484
transform 1 0 8740 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25576 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _0803_
timestamp 1666464484
transform 1 0 24564 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0804_
timestamp 1666464484
transform 1 0 21344 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0805_
timestamp 1666464484
transform 1 0 29900 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _0806_
timestamp 1666464484
transform 1 0 29716 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__a32o_1  _0807_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28060 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0808_
timestamp 1666464484
transform 1 0 16836 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0809_
timestamp 1666464484
transform 1 0 20516 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0810_
timestamp 1666464484
transform 1 0 20608 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0811_
timestamp 1666464484
transform 1 0 20792 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0812_
timestamp 1666464484
transform 1 0 21252 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _0813_
timestamp 1666464484
transform 1 0 22080 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_4  _0814_
timestamp 1666464484
transform 1 0 24564 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _0815_
timestamp 1666464484
transform 1 0 13524 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0816_
timestamp 1666464484
transform 1 0 13800 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0817_
timestamp 1666464484
transform 1 0 12236 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0819_
timestamp 1666464484
transform 1 0 12052 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _0820_
timestamp 1666464484
transform 1 0 12052 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0821_
timestamp 1666464484
transform 1 0 9752 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0822_
timestamp 1666464484
transform 1 0 10028 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0823_
timestamp 1666464484
transform 1 0 9844 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0824_
timestamp 1666464484
transform 1 0 8924 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0825_
timestamp 1666464484
transform 1 0 6164 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1666464484
transform 1 0 7084 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0827_
timestamp 1666464484
transform 1 0 7268 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0828_
timestamp 1666464484
transform 1 0 9108 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0829_
timestamp 1666464484
transform 1 0 9384 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _0830_
timestamp 1666464484
transform 1 0 8188 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _0831_
timestamp 1666464484
transform 1 0 4876 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _0832_
timestamp 1666464484
transform 1 0 5520 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0833_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2944 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0834_
timestamp 1666464484
transform 1 0 4232 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _0835_
timestamp 1666464484
transform 1 0 6532 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _0836_
timestamp 1666464484
transform 1 0 7544 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0837_
timestamp 1666464484
transform 1 0 3956 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0838_
timestamp 1666464484
transform 1 0 8280 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0839_
timestamp 1666464484
transform 1 0 7544 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0840_
timestamp 1666464484
transform 1 0 10580 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0841_
timestamp 1666464484
transform 1 0 10304 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0842_
timestamp 1666464484
transform 1 0 9108 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0843_
timestamp 1666464484
transform 1 0 9292 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0844_
timestamp 1666464484
transform 1 0 10304 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0845_
timestamp 1666464484
transform 1 0 9108 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0846_
timestamp 1666464484
transform 1 0 9660 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0847_
timestamp 1666464484
transform 1 0 9200 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0848_
timestamp 1666464484
transform 1 0 6532 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0849_
timestamp 1666464484
transform 1 0 5244 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0850_
timestamp 1666464484
transform 1 0 6440 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0851_
timestamp 1666464484
transform 1 0 6532 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _0852_
timestamp 1666464484
transform 1 0 4784 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0853_
timestamp 1666464484
transform 1 0 5060 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5152 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0855_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4416 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0856_
timestamp 1666464484
transform 1 0 3956 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0857_
timestamp 1666464484
transform 1 0 5336 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0858_
timestamp 1666464484
transform 1 0 4048 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0859_
timestamp 1666464484
transform 1 0 3036 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0860_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0861_
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _0862_
timestamp 1666464484
transform 1 0 3956 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0863_
timestamp 1666464484
transform 1 0 3220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0864_
timestamp 1666464484
transform 1 0 6716 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _0865_
timestamp 1666464484
transform 1 0 4968 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0866_
timestamp 1666464484
transform 1 0 10028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _0867_
timestamp 1666464484
transform 1 0 9476 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0868_
timestamp 1666464484
transform 1 0 7820 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0869_
timestamp 1666464484
transform 1 0 3036 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _0870_
timestamp 1666464484
transform 1 0 3956 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0871_
timestamp 1666464484
transform 1 0 26220 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0872_
timestamp 1666464484
transform 1 0 16836 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0873_
timestamp 1666464484
transform 1 0 21988 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0874_
timestamp 1666464484
transform 1 0 24656 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0875_
timestamp 1666464484
transform 1 0 28244 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0876_
timestamp 1666464484
transform 1 0 27968 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0877_
timestamp 1666464484
transform 1 0 27508 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0878_
timestamp 1666464484
transform 1 0 15824 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0879_
timestamp 1666464484
transform 1 0 24564 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0880_
timestamp 1666464484
transform 1 0 18308 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0881_
timestamp 1666464484
transform 1 0 12420 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0882_
timestamp 1666464484
transform 1 0 23368 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0883_
timestamp 1666464484
transform 1 0 23920 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0884_
timestamp 1666464484
transform 1 0 27784 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0885_
timestamp 1666464484
transform 1 0 13064 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0886_
timestamp 1666464484
transform 1 0 17572 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0887_
timestamp 1666464484
transform 1 0 13156 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0888_
timestamp 1666464484
transform 1 0 18400 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0889_
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0890_
timestamp 1666464484
transform 1 0 19412 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0891_
timestamp 1666464484
transform 1 0 12328 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0892_
timestamp 1666464484
transform 1 0 14720 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0893_
timestamp 1666464484
transform 1 0 12880 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0894_
timestamp 1666464484
transform 1 0 13248 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0895_
timestamp 1666464484
transform 1 0 15180 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0896_
timestamp 1666464484
transform 1 0 13248 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0897_
timestamp 1666464484
transform 1 0 22816 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0898_
timestamp 1666464484
transform 1 0 25300 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0899_
timestamp 1666464484
transform 1 0 25576 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0900_
timestamp 1666464484
transform 1 0 24840 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0901_
timestamp 1666464484
transform 1 0 21988 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0902_
timestamp 1666464484
transform 1 0 27140 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0903_
timestamp 1666464484
transform 1 0 25576 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0904_
timestamp 1666464484
transform 1 0 20976 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0905_
timestamp 1666464484
transform 1 0 30636 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0906_
timestamp 1666464484
transform 1 0 29716 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0907_
timestamp 1666464484
transform 1 0 30544 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0908_
timestamp 1666464484
transform 1 0 29716 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0909_
timestamp 1666464484
transform 1 0 16100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0910_
timestamp 1666464484
transform 1 0 13524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0911_
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0912_
timestamp 1666464484
transform 1 0 15180 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0913_
timestamp 1666464484
transform 1 0 13340 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0914_
timestamp 1666464484
transform 1 0 13248 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0915_
timestamp 1666464484
transform 1 0 14260 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0916_
timestamp 1666464484
transform 1 0 15180 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0917_
timestamp 1666464484
transform 1 0 19964 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0918_
timestamp 1666464484
transform 1 0 16836 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0919_
timestamp 1666464484
transform 1 0 20884 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0920_
timestamp 1666464484
transform 1 0 15824 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0921_
timestamp 1666464484
transform 1 0 26404 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0922_
timestamp 1666464484
transform 1 0 26128 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0923_
timestamp 1666464484
transform 1 0 27508 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0924_
timestamp 1666464484
transform 1 0 28612 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0925_
timestamp 1666464484
transform 1 0 23000 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0926_
timestamp 1666464484
transform 1 0 20976 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0927_
timestamp 1666464484
transform 1 0 23184 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0928_
timestamp 1666464484
transform 1 0 23368 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0929_
timestamp 1666464484
transform 1 0 25852 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0930_
timestamp 1666464484
transform 1 0 26128 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0931_
timestamp 1666464484
transform 1 0 27140 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0932_
timestamp 1666464484
transform 1 0 25760 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0933_
timestamp 1666464484
transform 1 0 29716 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0934_
timestamp 1666464484
transform 1 0 31280 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0935_
timestamp 1666464484
transform 1 0 32292 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0936_
timestamp 1666464484
transform 1 0 31004 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0937_
timestamp 1666464484
transform 1 0 28520 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0938_
timestamp 1666464484
transform 1 0 30636 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0939_
timestamp 1666464484
transform 1 0 31832 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0940_
timestamp 1666464484
transform 1 0 30360 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0941_
timestamp 1666464484
transform 1 0 27232 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0942_
timestamp 1666464484
transform 1 0 30820 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0943_
timestamp 1666464484
transform 1 0 31280 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0944_
timestamp 1666464484
transform 1 0 32292 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0945_
timestamp 1666464484
transform 1 0 16836 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0946_
timestamp 1666464484
transform 1 0 15640 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0947_
timestamp 1666464484
transform 1 0 18032 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0948_
timestamp 1666464484
transform 1 0 17848 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0949_
timestamp 1666464484
transform 1 0 22448 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0950_
timestamp 1666464484
transform 1 0 25852 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0951_
timestamp 1666464484
transform 1 0 22448 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0952_
timestamp 1666464484
transform 1 0 23184 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0953_
timestamp 1666464484
transform 1 0 20424 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0954_
timestamp 1666464484
transform 1 0 21620 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0955_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0956_
timestamp 1666464484
transform 1 0 5336 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0957_
timestamp 1666464484
transform 1 0 2576 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1666464484
transform 1 0 2392 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0959_
timestamp 1666464484
transform 1 0 14904 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0960_
timestamp 1666464484
transform 1 0 14260 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0961_
timestamp 1666464484
transform 1 0 14260 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0962_
timestamp 1666464484
transform 1 0 11684 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0963_
timestamp 1666464484
transform 1 0 2668 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0964_
timestamp 1666464484
transform 1 0 6348 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0965_
timestamp 1666464484
transform 1 0 9844 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0966_
timestamp 1666464484
transform 1 0 11316 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0967_
timestamp 1666464484
transform 1 0 6532 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0968_
timestamp 1666464484
transform 1 0 5612 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0969_
timestamp 1666464484
transform 1 0 10672 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0970_
timestamp 1666464484
transform 1 0 9568 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0971_
timestamp 1666464484
transform 1 0 6808 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0972_
timestamp 1666464484
transform 1 0 3956 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0973_
timestamp 1666464484
transform 1 0 4784 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0974__2
timestamp 1666464484
transform 1 0 14996 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975__3
timestamp 1666464484
transform 1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976__4
timestamp 1666464484
transform 1 0 17756 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977__5
timestamp 1666464484
transform 1 0 19596 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978__6
timestamp 1666464484
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979__7
timestamp 1666464484
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980__8
timestamp 1666464484
transform 1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0981_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18492 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1666464484
transform 1 0 18676 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1666464484
transform 1 0 13340 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1666464484
transform 1 0 12880 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1666464484
transform 1 0 14260 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1666464484
transform 1 0 14260 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1666464484
transform 1 0 22816 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1666464484
transform 1 0 24564 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1666464484
transform 1 0 24840 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1666464484
transform 1 0 24564 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1666464484
transform 1 0 21896 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1666464484
transform 1 0 24564 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1666464484
transform 1 0 22080 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1666464484
transform 1 0 21988 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1666464484
transform 1 0 28704 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1666464484
transform 1 0 29716 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1666464484
transform 1 0 27784 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1666464484
transform 1 0 27784 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1666464484
transform 1 0 14260 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1666464484
transform 1 0 14352 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1666464484
transform 1 0 14444 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1666464484
transform 1 0 14444 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1666464484
transform 1 0 12328 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1666464484
transform 1 0 12696 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1666464484
transform 1 0 12328 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1666464484
transform 1 0 12880 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_4  _1007_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4600 0 1 5440
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_2  _1008_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1564 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1009_
timestamp 1666464484
transform 1 0 1840 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1010_
timestamp 1666464484
transform 1 0 12604 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1011_
timestamp 1666464484
transform 1 0 12788 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1012_
timestamp 1666464484
transform 1 0 12696 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1013_
timestamp 1666464484
transform 1 0 10672 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1014_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1840 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1666464484
transform 1 0 3956 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1666464484
transform 1 0 9108 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1666464484
transform 1 0 8740 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1666464484
transform 1 0 4600 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1666464484
transform 1 0 6532 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1666464484
transform 1 0 9476 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1666464484
transform 1 0 9292 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1666464484
transform 1 0 4600 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1666464484
transform 1 0 3864 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1666464484
transform 1 0 9108 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1666464484
transform 1 0 9108 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1666464484
transform 1 0 5428 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1027_
timestamp 1666464484
transform 1 0 5612 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1028_
timestamp 1666464484
transform 1 0 8924 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1029_
timestamp 1666464484
transform 1 0 9108 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1030_
timestamp 1666464484
transform 1 0 5152 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1031_
timestamp 1666464484
transform 1 0 5060 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1032_
timestamp 1666464484
transform 1 0 9108 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1033_
timestamp 1666464484
transform 1 0 9200 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1034_
timestamp 1666464484
transform 1 0 6532 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_4  _1035_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4324 0 1 30464
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1036_
timestamp 1666464484
transform 1 0 8924 0 -1 29376
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1037_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7820 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_1  _1038_
timestamp 1666464484
transform 1 0 3220 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_4  _1039_
timestamp 1666464484
transform 1 0 3036 0 -1 26112
box -38 -48 1786 592
use sky130_fd_sc_hd__dfrtp_2  _1040_
timestamp 1666464484
transform 1 0 3956 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1666464484
transform 1 0 14444 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1666464484
transform 1 0 16560 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1666464484
transform 1 0 17664 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1666464484
transform 1 0 19504 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1666464484
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1666464484
transform 1 0 22540 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1666464484
transform 1 0 23828 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1666464484
transform 1 0 19412 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1666464484
transform 1 0 16836 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1666464484
transform 1 0 19412 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1666464484
transform 1 0 15824 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1666464484
transform 1 0 26404 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1666464484
transform 1 0 27140 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1666464484
transform 1 0 27784 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1666464484
transform 1 0 28980 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1666464484
transform 1 0 21988 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1666464484
transform 1 0 20976 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1666464484
transform 1 0 22448 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1666464484
transform 1 0 23828 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1666464484
transform 1 0 25208 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1666464484
transform 1 0 25760 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1666464484
transform 1 0 25484 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1666464484
transform 1 0 25208 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1065_
timestamp 1666464484
transform 1 0 29164 0 -1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1066_
timestamp 1666464484
transform 1 0 31188 0 1 10880
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1067_
timestamp 1666464484
transform 1 0 32292 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1068_
timestamp 1666464484
transform 1 0 32292 0 -1 13056
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1069_
timestamp 1666464484
transform 1 0 29716 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1070_
timestamp 1666464484
transform 1 0 29440 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1071_
timestamp 1666464484
transform 1 0 29624 0 -1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1072_
timestamp 1666464484
transform 1 0 29716 0 1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1666464484
transform 1 0 27324 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1666464484
transform 1 0 29992 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1666464484
transform 1 0 30544 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1076_
timestamp 1666464484
transform 1 0 27600 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1077_
timestamp 1666464484
transform 1 0 15916 0 1 27200
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1666464484
transform 1 0 15456 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1666464484
transform 1 0 16836 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1080_
timestamp 1666464484
transform 1 0 17020 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1666464484
transform 1 0 22632 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1666464484
transform 1 0 24564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1083_
timestamp 1666464484
transform 1 0 23092 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1084_
timestamp 1666464484
transform 1 0 23368 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1666464484
transform 1 0 19412 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1666464484
transform 1 0 19228 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_21.result $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14444 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_22.result
timestamp 1666464484
transform 1 0 22540 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_23.result
timestamp 1666464484
transform 1 0 25576 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_24.result
timestamp 1666464484
transform 1 0 30820 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_25.result
timestamp 1666464484
transform 1 0 29716 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_26.result
timestamp 1666464484
transform 1 0 29716 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_27.result
timestamp 1666464484
transform 1 0 16284 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_28.result
timestamp 1666464484
transform 1 0 23644 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_29.result
timestamp 1666464484
transform 1 0 19412 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_30.result
timestamp 1666464484
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_31.result
timestamp 1666464484
transform 1 0 24656 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_32.result
timestamp 1666464484
transform 1 0 24564 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_33.result
timestamp 1666464484
transform 1 0 29624 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_50.result
timestamp 1666464484
transform 1 0 12696 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_53.result
timestamp 1666464484
transform 1 0 18216 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0460_
timestamp 1666464484
transform 1 0 26496 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1666464484
transform 1 0 15364 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_21.result
timestamp 1666464484
transform 1 0 12972 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_22.result
timestamp 1666464484
transform 1 0 20792 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_23.result
timestamp 1666464484
transform 1 0 23368 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_24.result
timestamp 1666464484
transform 1 0 28612 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_25.result
timestamp 1666464484
transform 1 0 28612 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_26.result
timestamp 1666464484
transform 1 0 28612 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_27.result
timestamp 1666464484
transform 1 0 12972 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_28.result
timestamp 1666464484
transform 1 0 20792 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_29.result
timestamp 1666464484
transform 1 0 18216 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_30.result
timestamp 1666464484
transform 1 0 12972 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_31.result
timestamp 1666464484
transform 1 0 23368 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_32.result
timestamp 1666464484
transform 1 0 20792 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_33.result
timestamp 1666464484
transform 1 0 28612 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_50.result
timestamp 1666464484
transform 1 0 10396 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_53.result
timestamp 1666464484
transform 1 0 12972 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0460_
timestamp 1666464484
transform 1 0 23368 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_21.result
timestamp 1666464484
transform 1 0 12972 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_22.result
timestamp 1666464484
transform 1 0 20792 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_23.result
timestamp 1666464484
transform 1 0 24748 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_24.result
timestamp 1666464484
transform 1 0 31188 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_25.result
timestamp 1666464484
transform 1 0 28612 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_26.result
timestamp 1666464484
transform 1 0 31188 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_27.result
timestamp 1666464484
transform 1 0 15640 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_28.result
timestamp 1666464484
transform 1 0 26036 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_29.result
timestamp 1666464484
transform 1 0 18216 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_30.result
timestamp 1666464484
transform 1 0 10396 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_31.result
timestamp 1666464484
transform 1 0 23368 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_32.result
timestamp 1666464484
transform 1 0 23368 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_33.result
timestamp 1666464484
transform 1 0 28612 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_50.result
timestamp 1666464484
transform 1 0 12972 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_53.result
timestamp 1666464484
transform 1 0 18216 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0460_
timestamp 1666464484
transform 1 0 26036 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1666464484
transform 1 0 12972 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1666464484
transform 1 0 18216 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1666464484
transform 1 0 7820 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1666464484
transform 1 0 15640 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  fanout28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23644 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout30
timestamp 1666464484
transform 1 0 28612 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout31
timestamp 1666464484
transform 1 0 25576 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout32
timestamp 1666464484
transform 1 0 25760 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout33
timestamp 1666464484
transform 1 0 23092 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23276 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout35
timestamp 1666464484
transform 1 0 15548 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26404 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout37
timestamp 1666464484
transform 1 0 14536 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout38
timestamp 1666464484
transform 1 0 16836 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout39
timestamp 1666464484
transform 1 0 14260 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout40
timestamp 1666464484
transform 1 0 21712 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout41
timestamp 1666464484
transform 1 0 14260 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1666464484
transform 1 0 32384 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout43
timestamp 1666464484
transform 1 0 22632 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout44
timestamp 1666464484
transform 1 0 14260 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13892 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout46
timestamp 1666464484
transform 1 0 11868 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout47
timestamp 1666464484
transform 1 0 11960 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout48
timestamp 1666464484
transform 1 0 11960 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout49
timestamp 1666464484
transform 1 0 22908 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout50
timestamp 1666464484
transform 1 0 29716 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout51
timestamp 1666464484
transform 1 0 23736 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout52
timestamp 1666464484
transform 1 0 23552 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout53
timestamp 1666464484
transform 1 0 10672 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout54
timestamp 1666464484
transform 1 0 6532 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout55
timestamp 1666464484
transform 1 0 7360 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout56
timestamp 1666464484
transform 1 0 14260 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1666464484
transform 1 0 9108 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1666464484
transform 1 0 11776 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1666464484
transform 1 0 15088 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1666464484
transform 1 0 18400 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1666464484
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1666464484
transform 1 0 25024 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1666464484
transform 1 0 28336 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1666464484
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1666464484
transform 1 0 34960 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1666464484
transform 1 0 37996 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1666464484
transform 1 0 5152 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1666464484
transform 1 0 1564 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output13
timestamp 1666464484
transform 1 0 15640 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output14
timestamp 1666464484
transform 1 0 17112 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output15
timestamp 1666464484
transform 1 0 18400 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output16
timestamp 1666464484
transform 1 0 20056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output17
timestamp 1666464484
transform 1 0 21988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output18
timestamp 1666464484
transform 1 0 23000 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output19
timestamp 1666464484
transform 1 0 24564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output20
timestamp 1666464484
transform 1 0 25944 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output21
timestamp 1666464484
transform 1 0 27416 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output22
timestamp 1666464484
transform 1 0 29716 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output23
timestamp 1666464484
transform 1 0 2392 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output24
timestamp 1666464484
transform 1 0 30636 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output25
timestamp 1666464484
transform 1 0 32292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output26
timestamp 1666464484
transform 1 0 3956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output27
timestamp 1666464484
transform 1 0 5336 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_58
timestamp 1666464484
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_59
timestamp 1666464484
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_60
timestamp 1666464484
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_61
timestamp 1666464484
transform 1 0 12696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_62
timestamp 1666464484
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_63
timestamp 1666464484
transform 1 0 33304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_64
timestamp 1666464484
transform 1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_65
timestamp 1666464484
transform 1 0 36248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_66
timestamp 1666464484
transform 1 0 37720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_67
timestamp 1666464484
transform 1 0 38088 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_68
timestamp 1666464484
transform 1 0 38088 0 -1 3264
box -38 -48 314 592
<< labels >>
flabel metal2 s 1766 39200 1822 40000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 8390 39200 8446 40000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 11702 39200 11758 40000 0 FreeSans 224 90 0 0 io_in[1]
port 2 nsew signal input
flabel metal2 s 15014 39200 15070 40000 0 FreeSans 224 90 0 0 io_in[2]
port 3 nsew signal input
flabel metal2 s 18326 39200 18382 40000 0 FreeSans 224 90 0 0 io_in[3]
port 4 nsew signal input
flabel metal2 s 21638 39200 21694 40000 0 FreeSans 224 90 0 0 io_in[4]
port 5 nsew signal input
flabel metal2 s 24950 39200 25006 40000 0 FreeSans 224 90 0 0 io_in[5]
port 6 nsew signal input
flabel metal2 s 28262 39200 28318 40000 0 FreeSans 224 90 0 0 io_in[6]
port 7 nsew signal input
flabel metal2 s 31574 39200 31630 40000 0 FreeSans 224 90 0 0 io_in[7]
port 8 nsew signal input
flabel metal2 s 34886 39200 34942 40000 0 FreeSans 224 90 0 0 io_in[8]
port 9 nsew signal input
flabel metal2 s 38198 39200 38254 40000 0 FreeSans 224 90 0 0 io_in[9]
port 10 nsew signal input
flabel metal3 s 39200 19864 40000 19984 0 FreeSans 480 0 0 0 io_oeb
port 11 nsew signal tristate
flabel metal2 s 846 0 902 800 0 FreeSans 224 90 0 0 io_out[0]
port 12 nsew signal tristate
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 io_out[10]
port 13 nsew signal tristate
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 io_out[11]
port 14 nsew signal tristate
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 io_out[12]
port 15 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 io_out[13]
port 16 nsew signal tristate
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 io_out[14]
port 17 nsew signal tristate
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 io_out[15]
port 18 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 io_out[16]
port 19 nsew signal tristate
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 io_out[17]
port 20 nsew signal tristate
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 io_out[18]
port 21 nsew signal tristate
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 io_out[19]
port 22 nsew signal tristate
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 io_out[1]
port 23 nsew signal tristate
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 io_out[20]
port 24 nsew signal tristate
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 io_out[21]
port 25 nsew signal tristate
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 io_out[22]
port 26 nsew signal tristate
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 io_out[23]
port 27 nsew signal tristate
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 io_out[24]
port 28 nsew signal tristate
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 io_out[25]
port 29 nsew signal tristate
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 io_out[26]
port 30 nsew signal tristate
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 io_out[2]
port 31 nsew signal tristate
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 io_out[3]
port 32 nsew signal tristate
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 io_out[4]
port 33 nsew signal tristate
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 io_out[5]
port 34 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 io_out[6]
port 35 nsew signal tristate
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 io_out[7]
port 36 nsew signal tristate
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 io_out[8]
port 37 nsew signal tristate
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 io_out[9]
port 38 nsew signal tristate
flabel metal2 s 5078 39200 5134 40000 0 FreeSans 224 90 0 0 rst
port 39 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
