magic
tech sky130B
magscale 1 2
timestamp 1681463275
<< obsli1 >>
rect 1104 2159 58880 61489
<< obsm1 >>
rect 842 76 59602 63300
<< metal2 >>
rect 846 63200 902 64000
rect 1582 63200 1638 64000
rect 2318 63200 2374 64000
rect 3054 63200 3110 64000
rect 3790 63200 3846 64000
rect 4526 63200 4582 64000
rect 5262 63200 5318 64000
rect 5998 63200 6054 64000
rect 6734 63200 6790 64000
rect 7470 63200 7526 64000
rect 8206 63200 8262 64000
rect 8942 63200 8998 64000
rect 9678 63200 9734 64000
rect 10414 63200 10470 64000
rect 11150 63200 11206 64000
rect 11886 63200 11942 64000
rect 12622 63200 12678 64000
rect 13358 63200 13414 64000
rect 14094 63200 14150 64000
rect 14830 63200 14886 64000
rect 15566 63200 15622 64000
rect 16302 63200 16358 64000
rect 17038 63200 17094 64000
rect 17774 63200 17830 64000
rect 18510 63200 18566 64000
rect 19246 63200 19302 64000
rect 19982 63200 20038 64000
rect 20718 63200 20774 64000
rect 21454 63200 21510 64000
rect 22190 63200 22246 64000
rect 22926 63200 22982 64000
rect 23662 63200 23718 64000
rect 24398 63200 24454 64000
rect 25134 63200 25190 64000
rect 25870 63200 25926 64000
rect 26606 63200 26662 64000
rect 27342 63200 27398 64000
rect 28078 63200 28134 64000
rect 28814 63200 28870 64000
rect 29550 63200 29606 64000
rect 30286 63200 30342 64000
rect 31022 63200 31078 64000
rect 31758 63200 31814 64000
rect 32494 63200 32550 64000
rect 33230 63200 33286 64000
rect 33966 63200 34022 64000
rect 34702 63200 34758 64000
rect 35438 63200 35494 64000
rect 36174 63200 36230 64000
rect 36910 63200 36966 64000
rect 37646 63200 37702 64000
rect 38382 63200 38438 64000
rect 39118 63200 39174 64000
rect 39854 63200 39910 64000
rect 40590 63200 40646 64000
rect 41326 63200 41382 64000
rect 42062 63200 42118 64000
rect 42798 63200 42854 64000
rect 43534 63200 43590 64000
rect 44270 63200 44326 64000
rect 45006 63200 45062 64000
rect 45742 63200 45798 64000
rect 46478 63200 46534 64000
rect 47214 63200 47270 64000
rect 47950 63200 48006 64000
rect 48686 63200 48742 64000
rect 49422 63200 49478 64000
rect 50158 63200 50214 64000
rect 50894 63200 50950 64000
rect 51630 63200 51686 64000
rect 52366 63200 52422 64000
rect 53102 63200 53158 64000
rect 53838 63200 53894 64000
rect 54574 63200 54630 64000
rect 55310 63200 55366 64000
rect 56046 63200 56102 64000
rect 56782 63200 56838 64000
rect 57518 63200 57574 64000
rect 58254 63200 58310 64000
rect 58990 63200 59046 64000
rect 4526 0 4582 800
rect 4802 0 4858 800
rect 5078 0 5134 800
rect 5354 0 5410 800
rect 5630 0 5686 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16394 0 16450 800
rect 16670 0 16726 800
rect 16946 0 17002 800
rect 17222 0 17278 800
rect 17498 0 17554 800
rect 17774 0 17830 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18878 0 18934 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19706 0 19762 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20534 0 20590 800
rect 20810 0 20866 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23846 0 23902 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34058 0 34114 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35438 0 35494 800
rect 35714 0 35770 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39854 0 39910 800
rect 40130 0 40186 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41510 0 41566 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43166 0 43222 800
rect 43442 0 43498 800
rect 43718 0 43774 800
rect 43994 0 44050 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45098 0 45154 800
rect 45374 0 45430 800
rect 45650 0 45706 800
rect 45926 0 45982 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48962 0 49018 800
rect 49238 0 49294 800
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50894 0 50950 800
rect 51170 0 51226 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52826 0 52882 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53654 0 53710 800
rect 53930 0 53986 800
rect 54206 0 54262 800
rect 54482 0 54538 800
rect 54758 0 54814 800
rect 55034 0 55090 800
rect 55310 0 55366 800
<< obsm2 >>
rect 958 63144 1526 63322
rect 1694 63144 2262 63322
rect 2430 63144 2998 63322
rect 3166 63144 3734 63322
rect 3902 63144 4470 63322
rect 4638 63144 5206 63322
rect 5374 63144 5942 63322
rect 6110 63144 6678 63322
rect 6846 63144 7414 63322
rect 7582 63144 8150 63322
rect 8318 63144 8886 63322
rect 9054 63144 9622 63322
rect 9790 63144 10358 63322
rect 10526 63144 11094 63322
rect 11262 63144 11830 63322
rect 11998 63144 12566 63322
rect 12734 63144 13302 63322
rect 13470 63144 14038 63322
rect 14206 63144 14774 63322
rect 14942 63144 15510 63322
rect 15678 63144 16246 63322
rect 16414 63144 16982 63322
rect 17150 63144 17718 63322
rect 17886 63144 18454 63322
rect 18622 63144 19190 63322
rect 19358 63144 19926 63322
rect 20094 63144 20662 63322
rect 20830 63144 21398 63322
rect 21566 63144 22134 63322
rect 22302 63144 22870 63322
rect 23038 63144 23606 63322
rect 23774 63144 24342 63322
rect 24510 63144 25078 63322
rect 25246 63144 25814 63322
rect 25982 63144 26550 63322
rect 26718 63144 27286 63322
rect 27454 63144 28022 63322
rect 28190 63144 28758 63322
rect 28926 63144 29494 63322
rect 29662 63144 30230 63322
rect 30398 63144 30966 63322
rect 31134 63144 31702 63322
rect 31870 63144 32438 63322
rect 32606 63144 33174 63322
rect 33342 63144 33910 63322
rect 34078 63144 34646 63322
rect 34814 63144 35382 63322
rect 35550 63144 36118 63322
rect 36286 63144 36854 63322
rect 37022 63144 37590 63322
rect 37758 63144 38326 63322
rect 38494 63144 39062 63322
rect 39230 63144 39798 63322
rect 39966 63144 40534 63322
rect 40702 63144 41270 63322
rect 41438 63144 42006 63322
rect 42174 63144 42742 63322
rect 42910 63144 43478 63322
rect 43646 63144 44214 63322
rect 44382 63144 44950 63322
rect 45118 63144 45686 63322
rect 45854 63144 46422 63322
rect 46590 63144 47158 63322
rect 47326 63144 47894 63322
rect 48062 63144 48630 63322
rect 48798 63144 49366 63322
rect 49534 63144 50102 63322
rect 50270 63144 50838 63322
rect 51006 63144 51574 63322
rect 51742 63144 52310 63322
rect 52478 63144 53046 63322
rect 53214 63144 53782 63322
rect 53950 63144 54518 63322
rect 54686 63144 55254 63322
rect 55422 63144 55990 63322
rect 56158 63144 56726 63322
rect 56894 63144 57462 63322
rect 57630 63144 58198 63322
rect 58366 63144 58934 63322
rect 59102 63144 59596 63322
rect 848 856 59596 63144
rect 848 70 4470 856
rect 4638 70 4746 856
rect 4914 70 5022 856
rect 5190 70 5298 856
rect 5466 70 5574 856
rect 5742 70 5850 856
rect 6018 70 6126 856
rect 6294 70 6402 856
rect 6570 70 6678 856
rect 6846 70 6954 856
rect 7122 70 7230 856
rect 7398 70 7506 856
rect 7674 70 7782 856
rect 7950 70 8058 856
rect 8226 70 8334 856
rect 8502 70 8610 856
rect 8778 70 8886 856
rect 9054 70 9162 856
rect 9330 70 9438 856
rect 9606 70 9714 856
rect 9882 70 9990 856
rect 10158 70 10266 856
rect 10434 70 10542 856
rect 10710 70 10818 856
rect 10986 70 11094 856
rect 11262 70 11370 856
rect 11538 70 11646 856
rect 11814 70 11922 856
rect 12090 70 12198 856
rect 12366 70 12474 856
rect 12642 70 12750 856
rect 12918 70 13026 856
rect 13194 70 13302 856
rect 13470 70 13578 856
rect 13746 70 13854 856
rect 14022 70 14130 856
rect 14298 70 14406 856
rect 14574 70 14682 856
rect 14850 70 14958 856
rect 15126 70 15234 856
rect 15402 70 15510 856
rect 15678 70 15786 856
rect 15954 70 16062 856
rect 16230 70 16338 856
rect 16506 70 16614 856
rect 16782 70 16890 856
rect 17058 70 17166 856
rect 17334 70 17442 856
rect 17610 70 17718 856
rect 17886 70 17994 856
rect 18162 70 18270 856
rect 18438 70 18546 856
rect 18714 70 18822 856
rect 18990 70 19098 856
rect 19266 70 19374 856
rect 19542 70 19650 856
rect 19818 70 19926 856
rect 20094 70 20202 856
rect 20370 70 20478 856
rect 20646 70 20754 856
rect 20922 70 21030 856
rect 21198 70 21306 856
rect 21474 70 21582 856
rect 21750 70 21858 856
rect 22026 70 22134 856
rect 22302 70 22410 856
rect 22578 70 22686 856
rect 22854 70 22962 856
rect 23130 70 23238 856
rect 23406 70 23514 856
rect 23682 70 23790 856
rect 23958 70 24066 856
rect 24234 70 24342 856
rect 24510 70 24618 856
rect 24786 70 24894 856
rect 25062 70 25170 856
rect 25338 70 25446 856
rect 25614 70 25722 856
rect 25890 70 25998 856
rect 26166 70 26274 856
rect 26442 70 26550 856
rect 26718 70 26826 856
rect 26994 70 27102 856
rect 27270 70 27378 856
rect 27546 70 27654 856
rect 27822 70 27930 856
rect 28098 70 28206 856
rect 28374 70 28482 856
rect 28650 70 28758 856
rect 28926 70 29034 856
rect 29202 70 29310 856
rect 29478 70 29586 856
rect 29754 70 29862 856
rect 30030 70 30138 856
rect 30306 70 30414 856
rect 30582 70 30690 856
rect 30858 70 30966 856
rect 31134 70 31242 856
rect 31410 70 31518 856
rect 31686 70 31794 856
rect 31962 70 32070 856
rect 32238 70 32346 856
rect 32514 70 32622 856
rect 32790 70 32898 856
rect 33066 70 33174 856
rect 33342 70 33450 856
rect 33618 70 33726 856
rect 33894 70 34002 856
rect 34170 70 34278 856
rect 34446 70 34554 856
rect 34722 70 34830 856
rect 34998 70 35106 856
rect 35274 70 35382 856
rect 35550 70 35658 856
rect 35826 70 35934 856
rect 36102 70 36210 856
rect 36378 70 36486 856
rect 36654 70 36762 856
rect 36930 70 37038 856
rect 37206 70 37314 856
rect 37482 70 37590 856
rect 37758 70 37866 856
rect 38034 70 38142 856
rect 38310 70 38418 856
rect 38586 70 38694 856
rect 38862 70 38970 856
rect 39138 70 39246 856
rect 39414 70 39522 856
rect 39690 70 39798 856
rect 39966 70 40074 856
rect 40242 70 40350 856
rect 40518 70 40626 856
rect 40794 70 40902 856
rect 41070 70 41178 856
rect 41346 70 41454 856
rect 41622 70 41730 856
rect 41898 70 42006 856
rect 42174 70 42282 856
rect 42450 70 42558 856
rect 42726 70 42834 856
rect 43002 70 43110 856
rect 43278 70 43386 856
rect 43554 70 43662 856
rect 43830 70 43938 856
rect 44106 70 44214 856
rect 44382 70 44490 856
rect 44658 70 44766 856
rect 44934 70 45042 856
rect 45210 70 45318 856
rect 45486 70 45594 856
rect 45762 70 45870 856
rect 46038 70 46146 856
rect 46314 70 46422 856
rect 46590 70 46698 856
rect 46866 70 46974 856
rect 47142 70 47250 856
rect 47418 70 47526 856
rect 47694 70 47802 856
rect 47970 70 48078 856
rect 48246 70 48354 856
rect 48522 70 48630 856
rect 48798 70 48906 856
rect 49074 70 49182 856
rect 49350 70 49458 856
rect 49626 70 49734 856
rect 49902 70 50010 856
rect 50178 70 50286 856
rect 50454 70 50562 856
rect 50730 70 50838 856
rect 51006 70 51114 856
rect 51282 70 51390 856
rect 51558 70 51666 856
rect 51834 70 51942 856
rect 52110 70 52218 856
rect 52386 70 52494 856
rect 52662 70 52770 856
rect 52938 70 53046 856
rect 53214 70 53322 856
rect 53490 70 53598 856
rect 53766 70 53874 856
rect 54042 70 54150 856
rect 54318 70 54426 856
rect 54594 70 54702 856
rect 54870 70 54978 856
rect 55146 70 55254 856
rect 55422 70 59596 856
<< metal3 >>
rect 59200 62568 60000 62688
rect 59200 62024 60000 62144
rect 0 61752 800 61872
rect 59200 61480 60000 61600
rect 0 61072 800 61192
rect 59200 60936 60000 61056
rect 0 60392 800 60512
rect 59200 60392 60000 60512
rect 0 59712 800 59832
rect 59200 59848 60000 59968
rect 59200 59304 60000 59424
rect 0 59032 800 59152
rect 59200 58760 60000 58880
rect 0 58352 800 58472
rect 59200 58216 60000 58336
rect 0 57672 800 57792
rect 59200 57672 60000 57792
rect 0 56992 800 57112
rect 59200 57128 60000 57248
rect 59200 56584 60000 56704
rect 0 56312 800 56432
rect 59200 56040 60000 56160
rect 0 55632 800 55752
rect 59200 55496 60000 55616
rect 0 54952 800 55072
rect 59200 54952 60000 55072
rect 0 54272 800 54392
rect 59200 54408 60000 54528
rect 59200 53864 60000 53984
rect 0 53592 800 53712
rect 59200 53320 60000 53440
rect 0 52912 800 53032
rect 59200 52776 60000 52896
rect 0 52232 800 52352
rect 59200 52232 60000 52352
rect 0 51552 800 51672
rect 59200 51688 60000 51808
rect 59200 51144 60000 51264
rect 0 50872 800 50992
rect 59200 50600 60000 50720
rect 0 50192 800 50312
rect 59200 50056 60000 50176
rect 0 49512 800 49632
rect 59200 49512 60000 49632
rect 0 48832 800 48952
rect 59200 48968 60000 49088
rect 59200 48424 60000 48544
rect 0 48152 800 48272
rect 59200 47880 60000 48000
rect 0 47472 800 47592
rect 59200 47336 60000 47456
rect 0 46792 800 46912
rect 59200 46792 60000 46912
rect 0 46112 800 46232
rect 59200 46248 60000 46368
rect 59200 45704 60000 45824
rect 0 45432 800 45552
rect 59200 45160 60000 45280
rect 0 44752 800 44872
rect 59200 44616 60000 44736
rect 0 44072 800 44192
rect 59200 44072 60000 44192
rect 0 43392 800 43512
rect 59200 43528 60000 43648
rect 59200 42984 60000 43104
rect 0 42712 800 42832
rect 59200 42440 60000 42560
rect 0 42032 800 42152
rect 59200 41896 60000 42016
rect 0 41352 800 41472
rect 59200 41352 60000 41472
rect 0 40672 800 40792
rect 59200 40808 60000 40928
rect 59200 40264 60000 40384
rect 0 39992 800 40112
rect 59200 39720 60000 39840
rect 0 39312 800 39432
rect 59200 39176 60000 39296
rect 0 38632 800 38752
rect 59200 38632 60000 38752
rect 0 37952 800 38072
rect 59200 38088 60000 38208
rect 59200 37544 60000 37664
rect 0 37272 800 37392
rect 59200 37000 60000 37120
rect 0 36592 800 36712
rect 59200 36456 60000 36576
rect 0 35912 800 36032
rect 59200 35912 60000 36032
rect 0 35232 800 35352
rect 59200 35368 60000 35488
rect 59200 34824 60000 34944
rect 0 34552 800 34672
rect 59200 34280 60000 34400
rect 0 33872 800 33992
rect 59200 33736 60000 33856
rect 0 33192 800 33312
rect 59200 33192 60000 33312
rect 0 32512 800 32632
rect 59200 32648 60000 32768
rect 59200 32104 60000 32224
rect 0 31832 800 31952
rect 59200 31560 60000 31680
rect 0 31152 800 31272
rect 59200 31016 60000 31136
rect 0 30472 800 30592
rect 59200 30472 60000 30592
rect 0 29792 800 29912
rect 59200 29928 60000 30048
rect 59200 29384 60000 29504
rect 0 29112 800 29232
rect 59200 28840 60000 28960
rect 0 28432 800 28552
rect 59200 28296 60000 28416
rect 0 27752 800 27872
rect 59200 27752 60000 27872
rect 0 27072 800 27192
rect 59200 27208 60000 27328
rect 59200 26664 60000 26784
rect 0 26392 800 26512
rect 59200 26120 60000 26240
rect 0 25712 800 25832
rect 59200 25576 60000 25696
rect 0 25032 800 25152
rect 59200 25032 60000 25152
rect 0 24352 800 24472
rect 59200 24488 60000 24608
rect 59200 23944 60000 24064
rect 0 23672 800 23792
rect 59200 23400 60000 23520
rect 0 22992 800 23112
rect 59200 22856 60000 22976
rect 0 22312 800 22432
rect 59200 22312 60000 22432
rect 0 21632 800 21752
rect 59200 21768 60000 21888
rect 59200 21224 60000 21344
rect 0 20952 800 21072
rect 59200 20680 60000 20800
rect 0 20272 800 20392
rect 59200 20136 60000 20256
rect 0 19592 800 19712
rect 59200 19592 60000 19712
rect 0 18912 800 19032
rect 59200 19048 60000 19168
rect 59200 18504 60000 18624
rect 0 18232 800 18352
rect 59200 17960 60000 18080
rect 0 17552 800 17672
rect 59200 17416 60000 17536
rect 0 16872 800 16992
rect 59200 16872 60000 16992
rect 0 16192 800 16312
rect 59200 16328 60000 16448
rect 59200 15784 60000 15904
rect 0 15512 800 15632
rect 59200 15240 60000 15360
rect 0 14832 800 14952
rect 59200 14696 60000 14816
rect 0 14152 800 14272
rect 59200 14152 60000 14272
rect 0 13472 800 13592
rect 59200 13608 60000 13728
rect 59200 13064 60000 13184
rect 0 12792 800 12912
rect 59200 12520 60000 12640
rect 0 12112 800 12232
rect 59200 11976 60000 12096
rect 0 11432 800 11552
rect 59200 11432 60000 11552
rect 0 10752 800 10872
rect 59200 10888 60000 11008
rect 59200 10344 60000 10464
rect 0 10072 800 10192
rect 59200 9800 60000 9920
rect 0 9392 800 9512
rect 59200 9256 60000 9376
rect 0 8712 800 8832
rect 59200 8712 60000 8832
rect 0 8032 800 8152
rect 59200 8168 60000 8288
rect 59200 7624 60000 7744
rect 0 7352 800 7472
rect 59200 7080 60000 7200
rect 0 6672 800 6792
rect 59200 6536 60000 6656
rect 0 5992 800 6112
rect 59200 5992 60000 6112
rect 0 5312 800 5432
rect 59200 5448 60000 5568
rect 59200 4904 60000 5024
rect 0 4632 800 4752
rect 59200 4360 60000 4480
rect 0 3952 800 4072
rect 59200 3816 60000 3936
rect 0 3272 800 3392
rect 59200 3272 60000 3392
rect 0 2592 800 2712
rect 59200 2728 60000 2848
rect 59200 2184 60000 2304
rect 0 1912 800 2032
rect 59200 1640 60000 1760
rect 59200 1096 60000 1216
<< obsm3 >>
rect 800 62488 59120 62661
rect 800 62224 59200 62488
rect 800 61952 59120 62224
rect 880 61944 59120 61952
rect 880 61680 59200 61944
rect 880 61672 59120 61680
rect 800 61400 59120 61672
rect 800 61272 59200 61400
rect 880 61136 59200 61272
rect 880 60992 59120 61136
rect 800 60856 59120 60992
rect 800 60592 59200 60856
rect 880 60312 59120 60592
rect 800 60048 59200 60312
rect 800 59912 59120 60048
rect 880 59768 59120 59912
rect 880 59632 59200 59768
rect 800 59504 59200 59632
rect 800 59232 59120 59504
rect 880 59224 59120 59232
rect 880 58960 59200 59224
rect 880 58952 59120 58960
rect 800 58680 59120 58952
rect 800 58552 59200 58680
rect 880 58416 59200 58552
rect 880 58272 59120 58416
rect 800 58136 59120 58272
rect 800 57872 59200 58136
rect 880 57592 59120 57872
rect 800 57328 59200 57592
rect 800 57192 59120 57328
rect 880 57048 59120 57192
rect 880 56912 59200 57048
rect 800 56784 59200 56912
rect 800 56512 59120 56784
rect 880 56504 59120 56512
rect 880 56240 59200 56504
rect 880 56232 59120 56240
rect 800 55960 59120 56232
rect 800 55832 59200 55960
rect 880 55696 59200 55832
rect 880 55552 59120 55696
rect 800 55416 59120 55552
rect 800 55152 59200 55416
rect 880 54872 59120 55152
rect 800 54608 59200 54872
rect 800 54472 59120 54608
rect 880 54328 59120 54472
rect 880 54192 59200 54328
rect 800 54064 59200 54192
rect 800 53792 59120 54064
rect 880 53784 59120 53792
rect 880 53520 59200 53784
rect 880 53512 59120 53520
rect 800 53240 59120 53512
rect 800 53112 59200 53240
rect 880 52976 59200 53112
rect 880 52832 59120 52976
rect 800 52696 59120 52832
rect 800 52432 59200 52696
rect 880 52152 59120 52432
rect 800 51888 59200 52152
rect 800 51752 59120 51888
rect 880 51608 59120 51752
rect 880 51472 59200 51608
rect 800 51344 59200 51472
rect 800 51072 59120 51344
rect 880 51064 59120 51072
rect 880 50800 59200 51064
rect 880 50792 59120 50800
rect 800 50520 59120 50792
rect 800 50392 59200 50520
rect 880 50256 59200 50392
rect 880 50112 59120 50256
rect 800 49976 59120 50112
rect 800 49712 59200 49976
rect 880 49432 59120 49712
rect 800 49168 59200 49432
rect 800 49032 59120 49168
rect 880 48888 59120 49032
rect 880 48752 59200 48888
rect 800 48624 59200 48752
rect 800 48352 59120 48624
rect 880 48344 59120 48352
rect 880 48080 59200 48344
rect 880 48072 59120 48080
rect 800 47800 59120 48072
rect 800 47672 59200 47800
rect 880 47536 59200 47672
rect 880 47392 59120 47536
rect 800 47256 59120 47392
rect 800 46992 59200 47256
rect 880 46712 59120 46992
rect 800 46448 59200 46712
rect 800 46312 59120 46448
rect 880 46168 59120 46312
rect 880 46032 59200 46168
rect 800 45904 59200 46032
rect 800 45632 59120 45904
rect 880 45624 59120 45632
rect 880 45360 59200 45624
rect 880 45352 59120 45360
rect 800 45080 59120 45352
rect 800 44952 59200 45080
rect 880 44816 59200 44952
rect 880 44672 59120 44816
rect 800 44536 59120 44672
rect 800 44272 59200 44536
rect 880 43992 59120 44272
rect 800 43728 59200 43992
rect 800 43592 59120 43728
rect 880 43448 59120 43592
rect 880 43312 59200 43448
rect 800 43184 59200 43312
rect 800 42912 59120 43184
rect 880 42904 59120 42912
rect 880 42640 59200 42904
rect 880 42632 59120 42640
rect 800 42360 59120 42632
rect 800 42232 59200 42360
rect 880 42096 59200 42232
rect 880 41952 59120 42096
rect 800 41816 59120 41952
rect 800 41552 59200 41816
rect 880 41272 59120 41552
rect 800 41008 59200 41272
rect 800 40872 59120 41008
rect 880 40728 59120 40872
rect 880 40592 59200 40728
rect 800 40464 59200 40592
rect 800 40192 59120 40464
rect 880 40184 59120 40192
rect 880 39920 59200 40184
rect 880 39912 59120 39920
rect 800 39640 59120 39912
rect 800 39512 59200 39640
rect 880 39376 59200 39512
rect 880 39232 59120 39376
rect 800 39096 59120 39232
rect 800 38832 59200 39096
rect 880 38552 59120 38832
rect 800 38288 59200 38552
rect 800 38152 59120 38288
rect 880 38008 59120 38152
rect 880 37872 59200 38008
rect 800 37744 59200 37872
rect 800 37472 59120 37744
rect 880 37464 59120 37472
rect 880 37200 59200 37464
rect 880 37192 59120 37200
rect 800 36920 59120 37192
rect 800 36792 59200 36920
rect 880 36656 59200 36792
rect 880 36512 59120 36656
rect 800 36376 59120 36512
rect 800 36112 59200 36376
rect 880 35832 59120 36112
rect 800 35568 59200 35832
rect 800 35432 59120 35568
rect 880 35288 59120 35432
rect 880 35152 59200 35288
rect 800 35024 59200 35152
rect 800 34752 59120 35024
rect 880 34744 59120 34752
rect 880 34480 59200 34744
rect 880 34472 59120 34480
rect 800 34200 59120 34472
rect 800 34072 59200 34200
rect 880 33936 59200 34072
rect 880 33792 59120 33936
rect 800 33656 59120 33792
rect 800 33392 59200 33656
rect 880 33112 59120 33392
rect 800 32848 59200 33112
rect 800 32712 59120 32848
rect 880 32568 59120 32712
rect 880 32432 59200 32568
rect 800 32304 59200 32432
rect 800 32032 59120 32304
rect 880 32024 59120 32032
rect 880 31760 59200 32024
rect 880 31752 59120 31760
rect 800 31480 59120 31752
rect 800 31352 59200 31480
rect 880 31216 59200 31352
rect 880 31072 59120 31216
rect 800 30936 59120 31072
rect 800 30672 59200 30936
rect 880 30392 59120 30672
rect 800 30128 59200 30392
rect 800 29992 59120 30128
rect 880 29848 59120 29992
rect 880 29712 59200 29848
rect 800 29584 59200 29712
rect 800 29312 59120 29584
rect 880 29304 59120 29312
rect 880 29040 59200 29304
rect 880 29032 59120 29040
rect 800 28760 59120 29032
rect 800 28632 59200 28760
rect 880 28496 59200 28632
rect 880 28352 59120 28496
rect 800 28216 59120 28352
rect 800 27952 59200 28216
rect 880 27672 59120 27952
rect 800 27408 59200 27672
rect 800 27272 59120 27408
rect 880 27128 59120 27272
rect 880 26992 59200 27128
rect 800 26864 59200 26992
rect 800 26592 59120 26864
rect 880 26584 59120 26592
rect 880 26320 59200 26584
rect 880 26312 59120 26320
rect 800 26040 59120 26312
rect 800 25912 59200 26040
rect 880 25776 59200 25912
rect 880 25632 59120 25776
rect 800 25496 59120 25632
rect 800 25232 59200 25496
rect 880 24952 59120 25232
rect 800 24688 59200 24952
rect 800 24552 59120 24688
rect 880 24408 59120 24552
rect 880 24272 59200 24408
rect 800 24144 59200 24272
rect 800 23872 59120 24144
rect 880 23864 59120 23872
rect 880 23600 59200 23864
rect 880 23592 59120 23600
rect 800 23320 59120 23592
rect 800 23192 59200 23320
rect 880 23056 59200 23192
rect 880 22912 59120 23056
rect 800 22776 59120 22912
rect 800 22512 59200 22776
rect 880 22232 59120 22512
rect 800 21968 59200 22232
rect 800 21832 59120 21968
rect 880 21688 59120 21832
rect 880 21552 59200 21688
rect 800 21424 59200 21552
rect 800 21152 59120 21424
rect 880 21144 59120 21152
rect 880 20880 59200 21144
rect 880 20872 59120 20880
rect 800 20600 59120 20872
rect 800 20472 59200 20600
rect 880 20336 59200 20472
rect 880 20192 59120 20336
rect 800 20056 59120 20192
rect 800 19792 59200 20056
rect 880 19512 59120 19792
rect 800 19248 59200 19512
rect 800 19112 59120 19248
rect 880 18968 59120 19112
rect 880 18832 59200 18968
rect 800 18704 59200 18832
rect 800 18432 59120 18704
rect 880 18424 59120 18432
rect 880 18160 59200 18424
rect 880 18152 59120 18160
rect 800 17880 59120 18152
rect 800 17752 59200 17880
rect 880 17616 59200 17752
rect 880 17472 59120 17616
rect 800 17336 59120 17472
rect 800 17072 59200 17336
rect 880 16792 59120 17072
rect 800 16528 59200 16792
rect 800 16392 59120 16528
rect 880 16248 59120 16392
rect 880 16112 59200 16248
rect 800 15984 59200 16112
rect 800 15712 59120 15984
rect 880 15704 59120 15712
rect 880 15440 59200 15704
rect 880 15432 59120 15440
rect 800 15160 59120 15432
rect 800 15032 59200 15160
rect 880 14896 59200 15032
rect 880 14752 59120 14896
rect 800 14616 59120 14752
rect 800 14352 59200 14616
rect 880 14072 59120 14352
rect 800 13808 59200 14072
rect 800 13672 59120 13808
rect 880 13528 59120 13672
rect 880 13392 59200 13528
rect 800 13264 59200 13392
rect 800 12992 59120 13264
rect 880 12984 59120 12992
rect 880 12720 59200 12984
rect 880 12712 59120 12720
rect 800 12440 59120 12712
rect 800 12312 59200 12440
rect 880 12176 59200 12312
rect 880 12032 59120 12176
rect 800 11896 59120 12032
rect 800 11632 59200 11896
rect 880 11352 59120 11632
rect 800 11088 59200 11352
rect 800 10952 59120 11088
rect 880 10808 59120 10952
rect 880 10672 59200 10808
rect 800 10544 59200 10672
rect 800 10272 59120 10544
rect 880 10264 59120 10272
rect 880 10000 59200 10264
rect 880 9992 59120 10000
rect 800 9720 59120 9992
rect 800 9592 59200 9720
rect 880 9456 59200 9592
rect 880 9312 59120 9456
rect 800 9176 59120 9312
rect 800 8912 59200 9176
rect 880 8632 59120 8912
rect 800 8368 59200 8632
rect 800 8232 59120 8368
rect 880 8088 59120 8232
rect 880 7952 59200 8088
rect 800 7824 59200 7952
rect 800 7552 59120 7824
rect 880 7544 59120 7552
rect 880 7280 59200 7544
rect 880 7272 59120 7280
rect 800 7000 59120 7272
rect 800 6872 59200 7000
rect 880 6736 59200 6872
rect 880 6592 59120 6736
rect 800 6456 59120 6592
rect 800 6192 59200 6456
rect 880 5912 59120 6192
rect 800 5648 59200 5912
rect 800 5512 59120 5648
rect 880 5368 59120 5512
rect 880 5232 59200 5368
rect 800 5104 59200 5232
rect 800 4832 59120 5104
rect 880 4824 59120 4832
rect 880 4560 59200 4824
rect 880 4552 59120 4560
rect 800 4280 59120 4552
rect 800 4152 59200 4280
rect 880 4016 59200 4152
rect 880 3872 59120 4016
rect 800 3736 59120 3872
rect 800 3472 59200 3736
rect 880 3192 59120 3472
rect 800 2928 59200 3192
rect 800 2792 59120 2928
rect 880 2648 59120 2792
rect 880 2512 59200 2648
rect 800 2384 59200 2512
rect 800 2112 59120 2384
rect 880 2104 59120 2112
rect 880 1840 59200 2104
rect 880 1832 59120 1840
rect 800 1560 59120 1832
rect 800 1296 59200 1560
rect 800 1123 59120 1296
<< metal4 >>
rect 4208 2128 4528 61520
rect 19568 2128 19888 61520
rect 34928 2128 35248 61520
rect 50288 2128 50608 61520
<< obsm4 >>
rect 15883 2347 19488 60757
rect 19968 2347 34848 60757
rect 35328 2347 43917 60757
<< labels >>
rlabel metal3 s 0 20952 800 21072 6 design_clk_o
port 1 nsew signal output
rlabel metal3 s 0 1912 800 2032 6 dsi_all[0]
port 2 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 dsi_all[10]
port 3 nsew signal output
rlabel metal3 s 0 9392 800 9512 6 dsi_all[11]
port 4 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 dsi_all[12]
port 5 nsew signal output
rlabel metal3 s 0 10752 800 10872 6 dsi_all[13]
port 6 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 dsi_all[14]
port 7 nsew signal output
rlabel metal3 s 0 12112 800 12232 6 dsi_all[15]
port 8 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 dsi_all[16]
port 9 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 dsi_all[17]
port 10 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 dsi_all[18]
port 11 nsew signal output
rlabel metal3 s 0 14832 800 14952 6 dsi_all[19]
port 12 nsew signal output
rlabel metal3 s 0 2592 800 2712 6 dsi_all[1]
port 13 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 dsi_all[20]
port 14 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 dsi_all[21]
port 15 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 dsi_all[22]
port 16 nsew signal output
rlabel metal3 s 0 17552 800 17672 6 dsi_all[23]
port 17 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 dsi_all[24]
port 18 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 dsi_all[25]
port 19 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 dsi_all[26]
port 20 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 dsi_all[27]
port 21 nsew signal output
rlabel metal3 s 0 3272 800 3392 6 dsi_all[2]
port 22 nsew signal output
rlabel metal3 s 0 3952 800 4072 6 dsi_all[3]
port 23 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 dsi_all[4]
port 24 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 dsi_all[5]
port 25 nsew signal output
rlabel metal3 s 0 5992 800 6112 6 dsi_all[6]
port 26 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 dsi_all[7]
port 27 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 dsi_all[8]
port 28 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 dsi_all[9]
port 29 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 dso_6502[0]
port 30 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 dso_6502[10]
port 31 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 dso_6502[11]
port 32 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 dso_6502[12]
port 33 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 dso_6502[13]
port 34 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 dso_6502[14]
port 35 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 dso_6502[15]
port 36 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 dso_6502[16]
port 37 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 dso_6502[17]
port 38 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 dso_6502[18]
port 39 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 dso_6502[19]
port 40 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 dso_6502[1]
port 41 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 dso_6502[20]
port 42 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 dso_6502[21]
port 43 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 dso_6502[22]
port 44 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 dso_6502[23]
port 45 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 dso_6502[24]
port 46 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 dso_6502[25]
port 47 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 dso_6502[26]
port 48 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 dso_6502[2]
port 49 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 dso_6502[3]
port 50 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 dso_6502[4]
port 51 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 dso_6502[5]
port 52 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 dso_6502[6]
port 53 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 dso_6502[7]
port 54 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 dso_6502[8]
port 55 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 dso_6502[9]
port 56 nsew signal input
rlabel metal2 s 53838 63200 53894 64000 6 dso_LCD[0]
port 57 nsew signal input
rlabel metal2 s 54574 63200 54630 64000 6 dso_LCD[1]
port 58 nsew signal input
rlabel metal2 s 55310 63200 55366 64000 6 dso_LCD[2]
port 59 nsew signal input
rlabel metal2 s 56046 63200 56102 64000 6 dso_LCD[3]
port 60 nsew signal input
rlabel metal2 s 56782 63200 56838 64000 6 dso_LCD[4]
port 61 nsew signal input
rlabel metal2 s 57518 63200 57574 64000 6 dso_LCD[5]
port 62 nsew signal input
rlabel metal2 s 58254 63200 58310 64000 6 dso_LCD[6]
port 63 nsew signal input
rlabel metal2 s 58990 63200 59046 64000 6 dso_LCD[7]
port 64 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 dso_as1802[0]
port 65 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 dso_as1802[10]
port 66 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 dso_as1802[11]
port 67 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 dso_as1802[12]
port 68 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 dso_as1802[13]
port 69 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 dso_as1802[14]
port 70 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 dso_as1802[15]
port 71 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 dso_as1802[16]
port 72 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 dso_as1802[17]
port 73 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 dso_as1802[18]
port 74 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 dso_as1802[19]
port 75 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 dso_as1802[1]
port 76 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 dso_as1802[20]
port 77 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 dso_as1802[21]
port 78 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 dso_as1802[22]
port 79 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 dso_as1802[23]
port 80 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 dso_as1802[24]
port 81 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 dso_as1802[25]
port 82 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 dso_as1802[26]
port 83 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 dso_as1802[2]
port 84 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 dso_as1802[3]
port 85 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 dso_as1802[4]
port 86 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 dso_as1802[5]
port 87 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 dso_as1802[6]
port 88 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 dso_as1802[7]
port 89 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 dso_as1802[8]
port 90 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 dso_as1802[9]
port 91 nsew signal input
rlabel metal2 s 13358 63200 13414 64000 6 dso_as2650[0]
port 92 nsew signal input
rlabel metal2 s 20718 63200 20774 64000 6 dso_as2650[10]
port 93 nsew signal input
rlabel metal2 s 21454 63200 21510 64000 6 dso_as2650[11]
port 94 nsew signal input
rlabel metal2 s 22190 63200 22246 64000 6 dso_as2650[12]
port 95 nsew signal input
rlabel metal2 s 22926 63200 22982 64000 6 dso_as2650[13]
port 96 nsew signal input
rlabel metal2 s 23662 63200 23718 64000 6 dso_as2650[14]
port 97 nsew signal input
rlabel metal2 s 24398 63200 24454 64000 6 dso_as2650[15]
port 98 nsew signal input
rlabel metal2 s 25134 63200 25190 64000 6 dso_as2650[16]
port 99 nsew signal input
rlabel metal2 s 25870 63200 25926 64000 6 dso_as2650[17]
port 100 nsew signal input
rlabel metal2 s 26606 63200 26662 64000 6 dso_as2650[18]
port 101 nsew signal input
rlabel metal2 s 27342 63200 27398 64000 6 dso_as2650[19]
port 102 nsew signal input
rlabel metal2 s 14094 63200 14150 64000 6 dso_as2650[1]
port 103 nsew signal input
rlabel metal2 s 28078 63200 28134 64000 6 dso_as2650[20]
port 104 nsew signal input
rlabel metal2 s 28814 63200 28870 64000 6 dso_as2650[21]
port 105 nsew signal input
rlabel metal2 s 29550 63200 29606 64000 6 dso_as2650[22]
port 106 nsew signal input
rlabel metal2 s 30286 63200 30342 64000 6 dso_as2650[23]
port 107 nsew signal input
rlabel metal2 s 31022 63200 31078 64000 6 dso_as2650[24]
port 108 nsew signal input
rlabel metal2 s 31758 63200 31814 64000 6 dso_as2650[25]
port 109 nsew signal input
rlabel metal2 s 32494 63200 32550 64000 6 dso_as2650[26]
port 110 nsew signal input
rlabel metal2 s 14830 63200 14886 64000 6 dso_as2650[2]
port 111 nsew signal input
rlabel metal2 s 15566 63200 15622 64000 6 dso_as2650[3]
port 112 nsew signal input
rlabel metal2 s 16302 63200 16358 64000 6 dso_as2650[4]
port 113 nsew signal input
rlabel metal2 s 17038 63200 17094 64000 6 dso_as2650[5]
port 114 nsew signal input
rlabel metal2 s 17774 63200 17830 64000 6 dso_as2650[6]
port 115 nsew signal input
rlabel metal2 s 18510 63200 18566 64000 6 dso_as2650[7]
port 116 nsew signal input
rlabel metal2 s 19246 63200 19302 64000 6 dso_as2650[8]
port 117 nsew signal input
rlabel metal2 s 19982 63200 20038 64000 6 dso_as2650[9]
port 118 nsew signal input
rlabel metal3 s 0 42712 800 42832 6 dso_as512512512[0]
port 119 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 dso_as512512512[10]
port 120 nsew signal input
rlabel metal3 s 0 50192 800 50312 6 dso_as512512512[11]
port 121 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 dso_as512512512[12]
port 122 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 dso_as512512512[13]
port 123 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 dso_as512512512[14]
port 124 nsew signal input
rlabel metal3 s 0 52912 800 53032 6 dso_as512512512[15]
port 125 nsew signal input
rlabel metal3 s 0 53592 800 53712 6 dso_as512512512[16]
port 126 nsew signal input
rlabel metal3 s 0 54272 800 54392 6 dso_as512512512[17]
port 127 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 dso_as512512512[18]
port 128 nsew signal input
rlabel metal3 s 0 55632 800 55752 6 dso_as512512512[19]
port 129 nsew signal input
rlabel metal3 s 0 43392 800 43512 6 dso_as512512512[1]
port 130 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 dso_as512512512[20]
port 131 nsew signal input
rlabel metal3 s 0 56992 800 57112 6 dso_as512512512[21]
port 132 nsew signal input
rlabel metal3 s 0 57672 800 57792 6 dso_as512512512[22]
port 133 nsew signal input
rlabel metal3 s 0 58352 800 58472 6 dso_as512512512[23]
port 134 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 dso_as512512512[24]
port 135 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 dso_as512512512[25]
port 136 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 dso_as512512512[26]
port 137 nsew signal input
rlabel metal3 s 0 61072 800 61192 6 dso_as512512512[27]
port 138 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 dso_as512512512[2]
port 139 nsew signal input
rlabel metal3 s 0 44752 800 44872 6 dso_as512512512[3]
port 140 nsew signal input
rlabel metal3 s 0 45432 800 45552 6 dso_as512512512[4]
port 141 nsew signal input
rlabel metal3 s 0 46112 800 46232 6 dso_as512512512[5]
port 142 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 dso_as512512512[6]
port 143 nsew signal input
rlabel metal3 s 0 47472 800 47592 6 dso_as512512512[7]
port 144 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 dso_as512512512[8]
port 145 nsew signal input
rlabel metal3 s 0 48832 800 48952 6 dso_as512512512[9]
port 146 nsew signal input
rlabel metal2 s 33230 63200 33286 64000 6 dso_as5401[0]
port 147 nsew signal input
rlabel metal2 s 40590 63200 40646 64000 6 dso_as5401[10]
port 148 nsew signal input
rlabel metal2 s 41326 63200 41382 64000 6 dso_as5401[11]
port 149 nsew signal input
rlabel metal2 s 42062 63200 42118 64000 6 dso_as5401[12]
port 150 nsew signal input
rlabel metal2 s 42798 63200 42854 64000 6 dso_as5401[13]
port 151 nsew signal input
rlabel metal2 s 43534 63200 43590 64000 6 dso_as5401[14]
port 152 nsew signal input
rlabel metal2 s 44270 63200 44326 64000 6 dso_as5401[15]
port 153 nsew signal input
rlabel metal2 s 45006 63200 45062 64000 6 dso_as5401[16]
port 154 nsew signal input
rlabel metal2 s 45742 63200 45798 64000 6 dso_as5401[17]
port 155 nsew signal input
rlabel metal2 s 46478 63200 46534 64000 6 dso_as5401[18]
port 156 nsew signal input
rlabel metal2 s 47214 63200 47270 64000 6 dso_as5401[19]
port 157 nsew signal input
rlabel metal2 s 33966 63200 34022 64000 6 dso_as5401[1]
port 158 nsew signal input
rlabel metal2 s 47950 63200 48006 64000 6 dso_as5401[20]
port 159 nsew signal input
rlabel metal2 s 48686 63200 48742 64000 6 dso_as5401[21]
port 160 nsew signal input
rlabel metal2 s 49422 63200 49478 64000 6 dso_as5401[22]
port 161 nsew signal input
rlabel metal2 s 50158 63200 50214 64000 6 dso_as5401[23]
port 162 nsew signal input
rlabel metal2 s 50894 63200 50950 64000 6 dso_as5401[24]
port 163 nsew signal input
rlabel metal2 s 51630 63200 51686 64000 6 dso_as5401[25]
port 164 nsew signal input
rlabel metal2 s 52366 63200 52422 64000 6 dso_as5401[26]
port 165 nsew signal input
rlabel metal2 s 34702 63200 34758 64000 6 dso_as5401[2]
port 166 nsew signal input
rlabel metal2 s 35438 63200 35494 64000 6 dso_as5401[3]
port 167 nsew signal input
rlabel metal2 s 36174 63200 36230 64000 6 dso_as5401[4]
port 168 nsew signal input
rlabel metal2 s 36910 63200 36966 64000 6 dso_as5401[5]
port 169 nsew signal input
rlabel metal2 s 37646 63200 37702 64000 6 dso_as5401[6]
port 170 nsew signal input
rlabel metal2 s 38382 63200 38438 64000 6 dso_as5401[7]
port 171 nsew signal input
rlabel metal2 s 39118 63200 39174 64000 6 dso_as5401[8]
port 172 nsew signal input
rlabel metal2 s 39854 63200 39910 64000 6 dso_as5401[9]
port 173 nsew signal input
rlabel metal3 s 59200 56584 60000 56704 6 dso_counter[0]
port 174 nsew signal input
rlabel metal3 s 59200 62024 60000 62144 6 dso_counter[10]
port 175 nsew signal input
rlabel metal3 s 59200 62568 60000 62688 6 dso_counter[11]
port 176 nsew signal input
rlabel metal3 s 59200 57128 60000 57248 6 dso_counter[1]
port 177 nsew signal input
rlabel metal3 s 59200 57672 60000 57792 6 dso_counter[2]
port 178 nsew signal input
rlabel metal3 s 59200 58216 60000 58336 6 dso_counter[3]
port 179 nsew signal input
rlabel metal3 s 59200 58760 60000 58880 6 dso_counter[4]
port 180 nsew signal input
rlabel metal3 s 59200 59304 60000 59424 6 dso_counter[5]
port 181 nsew signal input
rlabel metal3 s 59200 59848 60000 59968 6 dso_counter[6]
port 182 nsew signal input
rlabel metal3 s 59200 60392 60000 60512 6 dso_counter[7]
port 183 nsew signal input
rlabel metal3 s 59200 60936 60000 61056 6 dso_counter[8]
port 184 nsew signal input
rlabel metal3 s 59200 61480 60000 61600 6 dso_counter[9]
port 185 nsew signal input
rlabel metal2 s 6734 63200 6790 64000 6 dso_diceroll[0]
port 186 nsew signal input
rlabel metal2 s 7470 63200 7526 64000 6 dso_diceroll[1]
port 187 nsew signal input
rlabel metal2 s 8206 63200 8262 64000 6 dso_diceroll[2]
port 188 nsew signal input
rlabel metal2 s 8942 63200 8998 64000 6 dso_diceroll[3]
port 189 nsew signal input
rlabel metal2 s 9678 63200 9734 64000 6 dso_diceroll[4]
port 190 nsew signal input
rlabel metal2 s 10414 63200 10470 64000 6 dso_diceroll[5]
port 191 nsew signal input
rlabel metal2 s 11150 63200 11206 64000 6 dso_diceroll[6]
port 192 nsew signal input
rlabel metal2 s 11886 63200 11942 64000 6 dso_diceroll[7]
port 193 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 dso_mc14500[0]
port 194 nsew signal input
rlabel metal3 s 0 31152 800 31272 6 dso_mc14500[1]
port 195 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 dso_mc14500[2]
port 196 nsew signal input
rlabel metal3 s 0 32512 800 32632 6 dso_mc14500[3]
port 197 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 dso_mc14500[4]
port 198 nsew signal input
rlabel metal3 s 0 33872 800 33992 6 dso_mc14500[5]
port 199 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 dso_mc14500[6]
port 200 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 dso_mc14500[7]
port 201 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 dso_mc14500[8]
port 202 nsew signal input
rlabel metal2 s 846 63200 902 64000 6 dso_multiplier[0]
port 203 nsew signal input
rlabel metal2 s 1582 63200 1638 64000 6 dso_multiplier[1]
port 204 nsew signal input
rlabel metal2 s 2318 63200 2374 64000 6 dso_multiplier[2]
port 205 nsew signal input
rlabel metal2 s 3054 63200 3110 64000 6 dso_multiplier[3]
port 206 nsew signal input
rlabel metal2 s 3790 63200 3846 64000 6 dso_multiplier[4]
port 207 nsew signal input
rlabel metal2 s 4526 63200 4582 64000 6 dso_multiplier[5]
port 208 nsew signal input
rlabel metal2 s 5262 63200 5318 64000 6 dso_multiplier[6]
port 209 nsew signal input
rlabel metal2 s 5998 63200 6054 64000 6 dso_multiplier[7]
port 210 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 dso_posit[0]
port 211 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 dso_posit[1]
port 212 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 dso_posit[2]
port 213 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 dso_posit[3]
port 214 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 dso_tbb1143[0]
port 215 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 dso_tbb1143[1]
port 216 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 dso_tbb1143[2]
port 217 nsew signal input
rlabel metal3 s 0 39312 800 39432 6 dso_tbb1143[3]
port 218 nsew signal input
rlabel metal3 s 0 39992 800 40112 6 dso_tbb1143[4]
port 219 nsew signal input
rlabel metal3 s 0 40672 800 40792 6 dso_tbb1143[5]
port 220 nsew signal input
rlabel metal3 s 0 41352 800 41472 6 dso_tbb1143[6]
port 221 nsew signal input
rlabel metal3 s 0 42032 800 42152 6 dso_tbb1143[7]
port 222 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 dso_tune
port 223 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 dso_vgatest[0]
port 224 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 dso_vgatest[1]
port 225 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 dso_vgatest[2]
port 226 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 dso_vgatest[3]
port 227 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 dso_vgatest[4]
port 228 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 dso_vgatest[5]
port 229 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 dso_vgatest[6]
port 230 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 dso_vgatest[7]
port 231 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 dso_vgatest[8]
port 232 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 dso_vgatest[9]
port 233 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 io_in[0]
port 234 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 io_in[10]
port 235 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 io_in[11]
port 236 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 io_in[12]
port 237 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 io_in[13]
port 238 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 io_in[14]
port 239 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 io_in[15]
port 240 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 io_in[16]
port 241 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 io_in[17]
port 242 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 io_in[18]
port 243 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 io_in[19]
port 244 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 io_in[1]
port 245 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 io_in[20]
port 246 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 io_in[21]
port 247 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 io_in[22]
port 248 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 io_in[23]
port 249 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 io_in[24]
port 250 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 io_in[25]
port 251 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 io_in[26]
port 252 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 io_in[27]
port 253 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 io_in[28]
port 254 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 io_in[29]
port 255 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 io_in[2]
port 256 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 io_in[30]
port 257 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 io_in[31]
port 258 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 io_in[32]
port 259 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 io_in[33]
port 260 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 io_in[34]
port 261 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 io_in[35]
port 262 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 io_in[36]
port 263 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 io_in[37]
port 264 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 io_in[3]
port 265 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 io_in[4]
port 266 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 io_in[5]
port 267 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 io_in[6]
port 268 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 io_in[7]
port 269 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 io_in[8]
port 270 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 io_in[9]
port 271 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 io_oeb[0]
port 272 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 io_oeb[10]
port 273 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 io_oeb[11]
port 274 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 io_oeb[12]
port 275 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 io_oeb[13]
port 276 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 io_oeb[14]
port 277 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 io_oeb[15]
port 278 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 io_oeb[16]
port 279 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 io_oeb[17]
port 280 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 io_oeb[18]
port 281 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 io_oeb[19]
port 282 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 io_oeb[1]
port 283 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 io_oeb[20]
port 284 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 io_oeb[21]
port 285 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 io_oeb[22]
port 286 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 io_oeb[23]
port 287 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 io_oeb[24]
port 288 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 io_oeb[25]
port 289 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 io_oeb[26]
port 290 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 io_oeb[27]
port 291 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 io_oeb[28]
port 292 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 io_oeb[29]
port 293 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 io_oeb[2]
port 294 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 io_oeb[30]
port 295 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 io_oeb[31]
port 296 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 io_oeb[32]
port 297 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 io_oeb[33]
port 298 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 io_oeb[34]
port 299 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 io_oeb[35]
port 300 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 io_oeb[36]
port 301 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 io_oeb[37]
port 302 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 io_oeb[3]
port 303 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 io_oeb[4]
port 304 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 io_oeb[5]
port 305 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 io_oeb[6]
port 306 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 io_oeb[7]
port 307 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 io_oeb[8]
port 308 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 io_oeb[9]
port 309 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 io_out[0]
port 310 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 io_out[10]
port 311 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 io_out[11]
port 312 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 io_out[12]
port 313 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 io_out[13]
port 314 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 io_out[14]
port 315 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 io_out[15]
port 316 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 io_out[16]
port 317 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 io_out[17]
port 318 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 io_out[18]
port 319 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 io_out[19]
port 320 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 io_out[1]
port 321 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 io_out[20]
port 322 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 io_out[21]
port 323 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 io_out[22]
port 324 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 io_out[23]
port 325 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 io_out[24]
port 326 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 io_out[25]
port 327 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 io_out[26]
port 328 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 io_out[27]
port 329 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 io_out[28]
port 330 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 io_out[29]
port 331 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 io_out[2]
port 332 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 io_out[30]
port 333 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 io_out[31]
port 334 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 io_out[32]
port 335 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 io_out[33]
port 336 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 io_out[34]
port 337 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 io_out[35]
port 338 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 io_out[36]
port 339 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 io_out[37]
port 340 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 io_out[3]
port 341 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 io_out[4]
port 342 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 io_out[5]
port 343 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 io_out[6]
port 344 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 io_out[7]
port 345 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 io_out[8]
port 346 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 io_out[9]
port 347 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 oeb_6502
port 348 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 oeb_as1802
port 349 nsew signal input
rlabel metal2 s 12622 63200 12678 64000 6 oeb_as2650
port 350 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 oeb_as512512512
port 351 nsew signal input
rlabel metal2 s 53102 63200 53158 64000 6 oeb_as5401
port 352 nsew signal input
rlabel metal3 s 0 36592 800 36712 6 oeb_mc14500
port 353 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 rst_6502
port 354 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 rst_LCD
port 355 nsew signal output
rlabel metal3 s 0 22992 800 23112 6 rst_as1802
port 356 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 rst_as2650
port 357 nsew signal output
rlabel metal3 s 0 25032 800 25152 6 rst_as512512512
port 358 nsew signal output
rlabel metal3 s 0 24352 800 24472 6 rst_as5401
port 359 nsew signal output
rlabel metal3 s 0 25712 800 25832 6 rst_counter
port 360 nsew signal output
rlabel metal3 s 0 26392 800 26512 6 rst_diceroll
port 361 nsew signal output
rlabel metal3 s 0 27072 800 27192 6 rst_mc14500
port 362 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 rst_posit
port 363 nsew signal output
rlabel metal3 s 0 28432 800 28552 6 rst_tbb1143
port 364 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 rst_tune
port 365 nsew signal output
rlabel metal3 s 0 29792 800 29912 6 rst_vgatest
port 366 nsew signal output
rlabel metal4 s 4208 2128 4528 61520 6 vccd1
port 367 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 61520 6 vccd1
port 367 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 61520 6 vssd1
port 368 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 61520 6 vssd1
port 368 nsew ground bidirectional
rlabel metal3 s 59200 1096 60000 1216 6 wb_clk_i
port 369 nsew signal input
rlabel metal3 s 59200 1640 60000 1760 6 wb_rst_i
port 370 nsew signal input
rlabel metal3 s 59200 2184 60000 2304 6 wbs_ack_o
port 371 nsew signal output
rlabel metal3 s 59200 4360 60000 4480 6 wbs_adr_i[0]
port 372 nsew signal input
rlabel metal3 s 59200 20680 60000 20800 6 wbs_adr_i[10]
port 373 nsew signal input
rlabel metal3 s 59200 22312 60000 22432 6 wbs_adr_i[11]
port 374 nsew signal input
rlabel metal3 s 59200 23944 60000 24064 6 wbs_adr_i[12]
port 375 nsew signal input
rlabel metal3 s 59200 25576 60000 25696 6 wbs_adr_i[13]
port 376 nsew signal input
rlabel metal3 s 59200 27208 60000 27328 6 wbs_adr_i[14]
port 377 nsew signal input
rlabel metal3 s 59200 28840 60000 28960 6 wbs_adr_i[15]
port 378 nsew signal input
rlabel metal3 s 59200 30472 60000 30592 6 wbs_adr_i[16]
port 379 nsew signal input
rlabel metal3 s 59200 32104 60000 32224 6 wbs_adr_i[17]
port 380 nsew signal input
rlabel metal3 s 59200 33736 60000 33856 6 wbs_adr_i[18]
port 381 nsew signal input
rlabel metal3 s 59200 35368 60000 35488 6 wbs_adr_i[19]
port 382 nsew signal input
rlabel metal3 s 59200 5992 60000 6112 6 wbs_adr_i[1]
port 383 nsew signal input
rlabel metal3 s 59200 37000 60000 37120 6 wbs_adr_i[20]
port 384 nsew signal input
rlabel metal3 s 59200 38632 60000 38752 6 wbs_adr_i[21]
port 385 nsew signal input
rlabel metal3 s 59200 40264 60000 40384 6 wbs_adr_i[22]
port 386 nsew signal input
rlabel metal3 s 59200 41896 60000 42016 6 wbs_adr_i[23]
port 387 nsew signal input
rlabel metal3 s 59200 43528 60000 43648 6 wbs_adr_i[24]
port 388 nsew signal input
rlabel metal3 s 59200 45160 60000 45280 6 wbs_adr_i[25]
port 389 nsew signal input
rlabel metal3 s 59200 46792 60000 46912 6 wbs_adr_i[26]
port 390 nsew signal input
rlabel metal3 s 59200 48424 60000 48544 6 wbs_adr_i[27]
port 391 nsew signal input
rlabel metal3 s 59200 50056 60000 50176 6 wbs_adr_i[28]
port 392 nsew signal input
rlabel metal3 s 59200 51688 60000 51808 6 wbs_adr_i[29]
port 393 nsew signal input
rlabel metal3 s 59200 7624 60000 7744 6 wbs_adr_i[2]
port 394 nsew signal input
rlabel metal3 s 59200 53320 60000 53440 6 wbs_adr_i[30]
port 395 nsew signal input
rlabel metal3 s 59200 54952 60000 55072 6 wbs_adr_i[31]
port 396 nsew signal input
rlabel metal3 s 59200 9256 60000 9376 6 wbs_adr_i[3]
port 397 nsew signal input
rlabel metal3 s 59200 10888 60000 11008 6 wbs_adr_i[4]
port 398 nsew signal input
rlabel metal3 s 59200 12520 60000 12640 6 wbs_adr_i[5]
port 399 nsew signal input
rlabel metal3 s 59200 14152 60000 14272 6 wbs_adr_i[6]
port 400 nsew signal input
rlabel metal3 s 59200 15784 60000 15904 6 wbs_adr_i[7]
port 401 nsew signal input
rlabel metal3 s 59200 17416 60000 17536 6 wbs_adr_i[8]
port 402 nsew signal input
rlabel metal3 s 59200 19048 60000 19168 6 wbs_adr_i[9]
port 403 nsew signal input
rlabel metal3 s 59200 2728 60000 2848 6 wbs_cyc_i
port 404 nsew signal input
rlabel metal3 s 59200 4904 60000 5024 6 wbs_dat_i[0]
port 405 nsew signal input
rlabel metal3 s 59200 21224 60000 21344 6 wbs_dat_i[10]
port 406 nsew signal input
rlabel metal3 s 59200 22856 60000 22976 6 wbs_dat_i[11]
port 407 nsew signal input
rlabel metal3 s 59200 24488 60000 24608 6 wbs_dat_i[12]
port 408 nsew signal input
rlabel metal3 s 59200 26120 60000 26240 6 wbs_dat_i[13]
port 409 nsew signal input
rlabel metal3 s 59200 27752 60000 27872 6 wbs_dat_i[14]
port 410 nsew signal input
rlabel metal3 s 59200 29384 60000 29504 6 wbs_dat_i[15]
port 411 nsew signal input
rlabel metal3 s 59200 31016 60000 31136 6 wbs_dat_i[16]
port 412 nsew signal input
rlabel metal3 s 59200 32648 60000 32768 6 wbs_dat_i[17]
port 413 nsew signal input
rlabel metal3 s 59200 34280 60000 34400 6 wbs_dat_i[18]
port 414 nsew signal input
rlabel metal3 s 59200 35912 60000 36032 6 wbs_dat_i[19]
port 415 nsew signal input
rlabel metal3 s 59200 6536 60000 6656 6 wbs_dat_i[1]
port 416 nsew signal input
rlabel metal3 s 59200 37544 60000 37664 6 wbs_dat_i[20]
port 417 nsew signal input
rlabel metal3 s 59200 39176 60000 39296 6 wbs_dat_i[21]
port 418 nsew signal input
rlabel metal3 s 59200 40808 60000 40928 6 wbs_dat_i[22]
port 419 nsew signal input
rlabel metal3 s 59200 42440 60000 42560 6 wbs_dat_i[23]
port 420 nsew signal input
rlabel metal3 s 59200 44072 60000 44192 6 wbs_dat_i[24]
port 421 nsew signal input
rlabel metal3 s 59200 45704 60000 45824 6 wbs_dat_i[25]
port 422 nsew signal input
rlabel metal3 s 59200 47336 60000 47456 6 wbs_dat_i[26]
port 423 nsew signal input
rlabel metal3 s 59200 48968 60000 49088 6 wbs_dat_i[27]
port 424 nsew signal input
rlabel metal3 s 59200 50600 60000 50720 6 wbs_dat_i[28]
port 425 nsew signal input
rlabel metal3 s 59200 52232 60000 52352 6 wbs_dat_i[29]
port 426 nsew signal input
rlabel metal3 s 59200 8168 60000 8288 6 wbs_dat_i[2]
port 427 nsew signal input
rlabel metal3 s 59200 53864 60000 53984 6 wbs_dat_i[30]
port 428 nsew signal input
rlabel metal3 s 59200 55496 60000 55616 6 wbs_dat_i[31]
port 429 nsew signal input
rlabel metal3 s 59200 9800 60000 9920 6 wbs_dat_i[3]
port 430 nsew signal input
rlabel metal3 s 59200 11432 60000 11552 6 wbs_dat_i[4]
port 431 nsew signal input
rlabel metal3 s 59200 13064 60000 13184 6 wbs_dat_i[5]
port 432 nsew signal input
rlabel metal3 s 59200 14696 60000 14816 6 wbs_dat_i[6]
port 433 nsew signal input
rlabel metal3 s 59200 16328 60000 16448 6 wbs_dat_i[7]
port 434 nsew signal input
rlabel metal3 s 59200 17960 60000 18080 6 wbs_dat_i[8]
port 435 nsew signal input
rlabel metal3 s 59200 19592 60000 19712 6 wbs_dat_i[9]
port 436 nsew signal input
rlabel metal3 s 59200 5448 60000 5568 6 wbs_dat_o[0]
port 437 nsew signal output
rlabel metal3 s 59200 21768 60000 21888 6 wbs_dat_o[10]
port 438 nsew signal output
rlabel metal3 s 59200 23400 60000 23520 6 wbs_dat_o[11]
port 439 nsew signal output
rlabel metal3 s 59200 25032 60000 25152 6 wbs_dat_o[12]
port 440 nsew signal output
rlabel metal3 s 59200 26664 60000 26784 6 wbs_dat_o[13]
port 441 nsew signal output
rlabel metal3 s 59200 28296 60000 28416 6 wbs_dat_o[14]
port 442 nsew signal output
rlabel metal3 s 59200 29928 60000 30048 6 wbs_dat_o[15]
port 443 nsew signal output
rlabel metal3 s 59200 31560 60000 31680 6 wbs_dat_o[16]
port 444 nsew signal output
rlabel metal3 s 59200 33192 60000 33312 6 wbs_dat_o[17]
port 445 nsew signal output
rlabel metal3 s 59200 34824 60000 34944 6 wbs_dat_o[18]
port 446 nsew signal output
rlabel metal3 s 59200 36456 60000 36576 6 wbs_dat_o[19]
port 447 nsew signal output
rlabel metal3 s 59200 7080 60000 7200 6 wbs_dat_o[1]
port 448 nsew signal output
rlabel metal3 s 59200 38088 60000 38208 6 wbs_dat_o[20]
port 449 nsew signal output
rlabel metal3 s 59200 39720 60000 39840 6 wbs_dat_o[21]
port 450 nsew signal output
rlabel metal3 s 59200 41352 60000 41472 6 wbs_dat_o[22]
port 451 nsew signal output
rlabel metal3 s 59200 42984 60000 43104 6 wbs_dat_o[23]
port 452 nsew signal output
rlabel metal3 s 59200 44616 60000 44736 6 wbs_dat_o[24]
port 453 nsew signal output
rlabel metal3 s 59200 46248 60000 46368 6 wbs_dat_o[25]
port 454 nsew signal output
rlabel metal3 s 59200 47880 60000 48000 6 wbs_dat_o[26]
port 455 nsew signal output
rlabel metal3 s 59200 49512 60000 49632 6 wbs_dat_o[27]
port 456 nsew signal output
rlabel metal3 s 59200 51144 60000 51264 6 wbs_dat_o[28]
port 457 nsew signal output
rlabel metal3 s 59200 52776 60000 52896 6 wbs_dat_o[29]
port 458 nsew signal output
rlabel metal3 s 59200 8712 60000 8832 6 wbs_dat_o[2]
port 459 nsew signal output
rlabel metal3 s 59200 54408 60000 54528 6 wbs_dat_o[30]
port 460 nsew signal output
rlabel metal3 s 59200 56040 60000 56160 6 wbs_dat_o[31]
port 461 nsew signal output
rlabel metal3 s 59200 10344 60000 10464 6 wbs_dat_o[3]
port 462 nsew signal output
rlabel metal3 s 59200 11976 60000 12096 6 wbs_dat_o[4]
port 463 nsew signal output
rlabel metal3 s 59200 13608 60000 13728 6 wbs_dat_o[5]
port 464 nsew signal output
rlabel metal3 s 59200 15240 60000 15360 6 wbs_dat_o[6]
port 465 nsew signal output
rlabel metal3 s 59200 16872 60000 16992 6 wbs_dat_o[7]
port 466 nsew signal output
rlabel metal3 s 59200 18504 60000 18624 6 wbs_dat_o[8]
port 467 nsew signal output
rlabel metal3 s 59200 20136 60000 20256 6 wbs_dat_o[9]
port 468 nsew signal output
rlabel metal3 s 59200 3272 60000 3392 6 wbs_stb_i
port 469 nsew signal input
rlabel metal3 s 59200 3816 60000 3936 6 wbs_we_i
port 470 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 64000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4585948
string GDS_FILE /media/lucah/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/Multiplexer/runs/23_04_14_11_03/results/signoff/multiplexer.magic.gds
string GDS_START 642702
<< end >>

