magic
tech sky130B
magscale 1 2
timestamp 1674825085
<< viali >>
rect 2789 15657 2823 15691
rect 5089 15657 5123 15691
rect 2053 15589 2087 15623
rect 4261 15589 4295 15623
rect 4445 15589 4479 15623
rect 2237 15521 2271 15555
rect 14289 15521 14323 15555
rect 15577 15521 15611 15555
rect 2973 15453 3007 15487
rect 4905 15453 4939 15487
rect 5917 15453 5951 15487
rect 9137 15453 9171 15487
rect 10333 15453 10367 15487
rect 11069 15453 11103 15487
rect 11897 15453 11931 15487
rect 12541 15453 12575 15487
rect 13001 15453 13035 15487
rect 14565 15453 14599 15487
rect 1777 15385 1811 15419
rect 3985 15385 4019 15419
rect 6009 15385 6043 15419
rect 6561 15385 6595 15419
rect 12449 15385 12483 15419
rect 7849 15317 7883 15351
rect 9321 15317 9355 15351
rect 10241 15317 10275 15351
rect 10977 15317 11011 15351
rect 11713 15317 11747 15351
rect 13093 15317 13127 15351
rect 13737 15317 13771 15351
rect 2053 15113 2087 15147
rect 2421 15113 2455 15147
rect 14381 15113 14415 15147
rect 4741 14977 4775 15011
rect 4997 14977 5031 15011
rect 6009 14977 6043 15011
rect 6561 14977 6595 15011
rect 8769 14977 8803 15011
rect 11161 14977 11195 15011
rect 11897 14977 11931 15011
rect 12357 14977 12391 15011
rect 13185 14977 13219 15011
rect 13829 14977 13863 15011
rect 14473 14977 14507 15011
rect 2513 14909 2547 14943
rect 2605 14909 2639 14943
rect 6837 14909 6871 14943
rect 8309 14909 8343 14943
rect 9045 14909 9079 14943
rect 10517 14909 10551 14943
rect 13737 14841 13771 14875
rect 3617 14773 3651 14807
rect 5917 14773 5951 14807
rect 11069 14773 11103 14807
rect 11805 14773 11839 14807
rect 12449 14773 12483 14807
rect 13001 14773 13035 14807
rect 15025 14773 15059 14807
rect 1593 14569 1627 14603
rect 3985 14569 4019 14603
rect 8125 14569 8159 14603
rect 9597 14569 9631 14603
rect 10504 14569 10538 14603
rect 4629 14433 4663 14467
rect 14381 14433 14415 14467
rect 2717 14365 2751 14399
rect 2973 14365 3007 14399
rect 8309 14365 8343 14399
rect 9781 14365 9815 14399
rect 10241 14365 10275 14399
rect 12633 14365 12667 14399
rect 13093 14365 13127 14399
rect 14473 14365 14507 14399
rect 4353 14297 4387 14331
rect 5273 14297 5307 14331
rect 4445 14229 4479 14263
rect 6561 14229 6595 14263
rect 11989 14229 12023 14263
rect 12541 14229 12575 14263
rect 13185 14229 13219 14263
rect 15025 14229 15059 14263
rect 1685 14025 1719 14059
rect 2421 14025 2455 14059
rect 4261 14025 4295 14059
rect 6561 14025 6595 14059
rect 8309 14025 8343 14059
rect 11805 14025 11839 14059
rect 3556 13957 3590 13991
rect 1869 13889 1903 13923
rect 3801 13889 3835 13923
rect 7389 13889 7423 13923
rect 9597 13889 9631 13923
rect 10241 13889 10275 13923
rect 10885 13889 10919 13923
rect 11805 13889 11839 13923
rect 12725 13889 12759 13923
rect 13645 13889 13679 13923
rect 14197 13889 14231 13923
rect 5733 13821 5767 13855
rect 6009 13821 6043 13855
rect 10149 13821 10183 13855
rect 10793 13821 10827 13855
rect 7205 13685 7239 13719
rect 12909 13685 12943 13719
rect 13553 13685 13587 13719
rect 14289 13685 14323 13719
rect 14933 13481 14967 13515
rect 4629 13413 4663 13447
rect 2605 13345 2639 13379
rect 6377 13345 6411 13379
rect 1869 13277 1903 13311
rect 2697 13277 2731 13311
rect 2789 13277 2823 13311
rect 3985 13277 4019 13311
rect 6837 13277 6871 13311
rect 9137 13277 9171 13311
rect 10701 13277 10735 13311
rect 11161 13277 11195 13311
rect 13645 13277 13679 13311
rect 14473 13277 14507 13311
rect 15117 13277 15151 13311
rect 4077 13209 4111 13243
rect 6101 13209 6135 13243
rect 7113 13209 7147 13243
rect 11437 13209 11471 13243
rect 1685 13141 1719 13175
rect 3157 13141 3191 13175
rect 8585 13141 8619 13175
rect 9321 13141 9355 13175
rect 10517 13141 10551 13175
rect 12909 13141 12943 13175
rect 13461 13141 13495 13175
rect 14381 13141 14415 13175
rect 2145 12937 2179 12971
rect 15117 12937 15151 12971
rect 2881 12869 2915 12903
rect 6561 12869 6595 12903
rect 8217 12869 8251 12903
rect 11989 12869 12023 12903
rect 13185 12869 13219 12903
rect 2053 12801 2087 12835
rect 4077 12801 4111 12835
rect 4537 12801 4571 12835
rect 4804 12801 4838 12835
rect 6653 12801 6687 12835
rect 6929 12801 6963 12835
rect 7665 12801 7699 12835
rect 8493 12801 8527 12835
rect 9045 12801 9079 12835
rect 12265 12801 12299 12835
rect 12909 12801 12943 12835
rect 15301 12801 15335 12835
rect 2329 12733 2363 12767
rect 9321 12733 9355 12767
rect 10793 12733 10827 12767
rect 14657 12733 14691 12767
rect 3157 12665 3191 12699
rect 3341 12665 3375 12699
rect 5917 12665 5951 12699
rect 1685 12597 1719 12631
rect 3985 12597 4019 12631
rect 7481 12597 7515 12631
rect 1685 12393 1719 12427
rect 15025 12393 15059 12427
rect 11529 12325 11563 12359
rect 3065 12257 3099 12291
rect 5825 12189 5859 12223
rect 6285 12189 6319 12223
rect 11345 12189 11379 12223
rect 12173 12189 12207 12223
rect 13185 12189 13219 12223
rect 14473 12189 14507 12223
rect 15117 12189 15151 12223
rect 15577 12189 15611 12223
rect 2820 12121 2854 12155
rect 4261 12121 4295 12155
rect 6561 12121 6595 12155
rect 10885 12121 10919 12155
rect 8033 12053 8067 12087
rect 9597 12053 9631 12087
rect 12173 12053 12207 12087
rect 13001 12053 13035 12087
rect 14381 12053 14415 12087
rect 5917 11849 5951 11883
rect 6745 11849 6779 11883
rect 7297 11849 7331 11883
rect 8217 11849 8251 11883
rect 16129 11849 16163 11883
rect 1593 11781 1627 11815
rect 12173 11781 12207 11815
rect 1777 11713 1811 11747
rect 2973 11713 3007 11747
rect 5825 11713 5859 11747
rect 6561 11713 6595 11747
rect 7297 11713 7331 11747
rect 7481 11713 7515 11747
rect 8033 11713 8067 11747
rect 9229 11713 9263 11747
rect 3433 11645 3467 11679
rect 3709 11645 3743 11679
rect 14381 11645 14415 11679
rect 14657 11645 14691 11679
rect 2973 11577 3007 11611
rect 1961 11509 1995 11543
rect 5181 11509 5215 11543
rect 10517 11509 10551 11543
rect 13645 11509 13679 11543
rect 2697 11305 2731 11339
rect 5628 11305 5662 11339
rect 9229 11305 9263 11339
rect 10241 11305 10275 11339
rect 1685 11237 1719 11271
rect 4537 11237 4571 11271
rect 7113 11237 7147 11271
rect 8401 11237 8435 11271
rect 13277 11237 13311 11271
rect 3433 11169 3467 11203
rect 10701 11169 10735 11203
rect 1869 11101 1903 11135
rect 2697 11101 2731 11135
rect 3249 11101 3283 11135
rect 4261 11101 4295 11135
rect 4445 11101 4479 11135
rect 5354 11101 5388 11135
rect 8033 11101 8067 11135
rect 8125 11101 8159 11135
rect 9413 11101 9447 11135
rect 9597 11101 9631 11135
rect 10057 11101 10091 11135
rect 12725 11101 12759 11135
rect 13369 11101 13403 11135
rect 14473 11101 14507 11135
rect 14933 11101 14967 11135
rect 15761 11101 15795 11135
rect 7849 11033 7883 11067
rect 8217 11033 8251 11067
rect 12449 11033 12483 11067
rect 15025 11033 15059 11067
rect 15669 11033 15703 11067
rect 14289 10965 14323 10999
rect 2513 10761 2547 10795
rect 7849 10761 7883 10795
rect 3801 10693 3835 10727
rect 4261 10693 4295 10727
rect 6561 10693 6595 10727
rect 11713 10693 11747 10727
rect 10077 10625 10111 10659
rect 10333 10625 10367 10659
rect 10977 10625 11011 10659
rect 13921 10625 13955 10659
rect 16129 10625 16163 10659
rect 6009 10557 6043 10591
rect 14197 10557 14231 10591
rect 8953 10421 8987 10455
rect 10885 10421 10919 10455
rect 13001 10421 13035 10455
rect 15669 10421 15703 10455
rect 16221 10421 16255 10455
rect 2973 10217 3007 10251
rect 5733 10217 5767 10251
rect 10885 10217 10919 10251
rect 13553 10217 13587 10251
rect 7573 10081 7607 10115
rect 7757 10081 7791 10115
rect 16037 10081 16071 10115
rect 1593 10013 1627 10047
rect 4537 10013 4571 10047
rect 7849 10013 7883 10047
rect 9321 10013 9355 10047
rect 9413 10013 9447 10047
rect 12909 10013 12943 10047
rect 13553 10013 13587 10047
rect 14289 10013 14323 10047
rect 1860 9945 1894 9979
rect 4169 9945 4203 9979
rect 4261 9945 4295 9979
rect 7021 9945 7055 9979
rect 12173 9945 12207 9979
rect 3985 9877 4019 9911
rect 4353 9877 4387 9911
rect 8217 9877 8251 9911
rect 9413 9877 9447 9911
rect 12725 9877 12759 9911
rect 3433 9605 3467 9639
rect 6561 9605 6595 9639
rect 2237 9537 2271 9571
rect 5641 9537 5675 9571
rect 5825 9537 5859 9571
rect 6653 9537 6687 9571
rect 6929 9537 6963 9571
rect 7389 9537 7423 9571
rect 8125 9537 8159 9571
rect 10701 9537 10735 9571
rect 10885 9537 10919 9571
rect 14197 9537 14231 9571
rect 3157 9469 3191 9503
rect 8401 9469 8435 9503
rect 11713 9469 11747 9503
rect 13461 9469 13495 9503
rect 13737 9469 13771 9503
rect 14473 9469 14507 9503
rect 2329 9401 2363 9435
rect 5917 9401 5951 9435
rect 10977 9401 11011 9435
rect 4905 9333 4939 9367
rect 7389 9333 7423 9367
rect 9873 9333 9907 9367
rect 15945 9333 15979 9367
rect 11805 9129 11839 9163
rect 13185 9129 13219 9163
rect 15117 9129 15151 9163
rect 12449 9061 12483 9095
rect 4445 8993 4479 9027
rect 6377 8993 6411 9027
rect 6653 8993 6687 9027
rect 10333 8993 10367 9027
rect 2973 8925 3007 8959
rect 4077 8925 4111 8959
rect 4353 8925 4387 8959
rect 8585 8925 8619 8959
rect 9505 8925 9539 8959
rect 9597 8925 9631 8959
rect 10057 8925 10091 8959
rect 12265 8925 12299 8959
rect 13001 8925 13035 8959
rect 14565 8925 14599 8959
rect 15301 8925 15335 8959
rect 15945 8925 15979 8959
rect 2728 8857 2762 8891
rect 8340 8857 8374 8891
rect 1593 8789 1627 8823
rect 4905 8789 4939 8823
rect 7205 8789 7239 8823
rect 14381 8789 14415 8823
rect 15853 8789 15887 8823
rect 1777 8585 1811 8619
rect 5089 8585 5123 8619
rect 15485 8585 15519 8619
rect 6929 8517 6963 8551
rect 1593 8449 1627 8483
rect 2789 8449 2823 8483
rect 5181 8449 5215 8483
rect 5641 8449 5675 8483
rect 5917 8449 5951 8483
rect 9781 8449 9815 8483
rect 11069 8449 11103 8483
rect 11713 8449 11747 8483
rect 11897 8449 11931 8483
rect 14657 8449 14691 8483
rect 15577 8449 15611 8483
rect 3065 8381 3099 8415
rect 7297 8381 7331 8415
rect 14381 8381 14415 8415
rect 4537 8313 4571 8347
rect 5917 8313 5951 8347
rect 11989 8313 12023 8347
rect 6745 8245 6779 8279
rect 6929 8245 6963 8279
rect 8309 8245 8343 8279
rect 11069 8245 11103 8279
rect 12909 8245 12943 8279
rect 1777 8041 1811 8075
rect 9321 8041 9355 8075
rect 13277 8041 13311 8075
rect 2697 7973 2731 8007
rect 4077 7973 4111 8007
rect 12081 7905 12115 7939
rect 1593 7837 1627 7871
rect 2697 7837 2731 7871
rect 3433 7837 3467 7871
rect 4169 7837 4203 7871
rect 4261 7837 4295 7871
rect 7021 7837 7055 7871
rect 8217 7837 8251 7871
rect 8401 7837 8435 7871
rect 8585 7837 8619 7871
rect 9137 7837 9171 7871
rect 13093 7837 13127 7871
rect 8309 7769 8343 7803
rect 11805 7769 11839 7803
rect 3249 7701 3283 7735
rect 5549 7701 5583 7735
rect 8033 7701 8067 7735
rect 10333 7701 10367 7735
rect 1593 7497 1627 7531
rect 3919 7497 3953 7531
rect 8309 7497 8343 7531
rect 10425 7497 10459 7531
rect 11897 7497 11931 7531
rect 2513 7429 2547 7463
rect 3709 7429 3743 7463
rect 9597 7429 9631 7463
rect 10057 7429 10091 7463
rect 1777 7361 1811 7395
rect 2697 7361 2731 7395
rect 2789 7361 2823 7395
rect 4537 7361 4571 7395
rect 5181 7361 5215 7395
rect 5457 7361 5491 7395
rect 5825 7361 5859 7395
rect 6561 7361 6595 7395
rect 10241 7361 10275 7395
rect 10333 7361 10367 7395
rect 11713 7361 11747 7395
rect 12633 7361 12667 7395
rect 13093 7361 13127 7395
rect 13277 7361 13311 7395
rect 2053 7293 2087 7327
rect 6837 7293 6871 7327
rect 10609 7293 10643 7327
rect 2513 7225 2547 7259
rect 5917 7225 5951 7259
rect 6745 7225 6779 7259
rect 13093 7225 13127 7259
rect 1961 7157 1995 7191
rect 3893 7157 3927 7191
rect 4077 7157 4111 7191
rect 6653 7157 6687 7191
rect 12449 7157 12483 7191
rect 1593 6953 1627 6987
rect 1961 6953 1995 6987
rect 4261 6953 4295 6987
rect 11633 6953 11667 6987
rect 4813 6817 4847 6851
rect 5089 6817 5123 6851
rect 6561 6817 6595 6851
rect 9229 6817 9263 6851
rect 1777 6749 1811 6783
rect 2053 6749 2087 6783
rect 2881 6749 2915 6783
rect 2973 6749 3007 6783
rect 3065 6749 3099 6783
rect 3249 6749 3283 6783
rect 4169 6749 4203 6783
rect 4353 6749 4387 6783
rect 7481 6749 7515 6783
rect 7573 6749 7607 6783
rect 9321 6749 9355 6783
rect 11897 6749 11931 6783
rect 12817 6749 12851 6783
rect 12909 6749 12943 6783
rect 7205 6681 7239 6715
rect 7941 6681 7975 6715
rect 8309 6681 8343 6715
rect 2605 6613 2639 6647
rect 8493 6613 8527 6647
rect 10149 6613 10183 6647
rect 1685 6409 1719 6443
rect 2329 6409 2363 6443
rect 3433 6409 3467 6443
rect 6837 6409 6871 6443
rect 8585 6409 8619 6443
rect 11805 6409 11839 6443
rect 5457 6341 5491 6375
rect 7665 6341 7699 6375
rect 7941 6341 7975 6375
rect 1869 6273 1903 6307
rect 2513 6273 2547 6307
rect 2697 6273 2731 6307
rect 2789 6273 2823 6307
rect 3525 6273 3559 6307
rect 5733 6273 5767 6307
rect 7205 6273 7239 6307
rect 7573 6273 7607 6307
rect 9137 6273 9171 6307
rect 9873 6273 9907 6307
rect 10425 6273 10459 6307
rect 10609 6273 10643 6307
rect 11713 6273 11747 6307
rect 11897 6273 11931 6307
rect 3985 6205 4019 6239
rect 8861 6205 8895 6239
rect 10701 6137 10735 6171
rect 6653 6069 6687 6103
rect 8769 6069 8803 6103
rect 9689 6069 9723 6103
rect 7021 5865 7055 5899
rect 11253 5865 11287 5899
rect 2053 5797 2087 5831
rect 1961 5729 1995 5763
rect 4445 5729 4479 5763
rect 9505 5729 9539 5763
rect 9781 5729 9815 5763
rect 1869 5661 1903 5695
rect 2145 5661 2179 5695
rect 2881 5661 2915 5695
rect 3157 5661 3191 5695
rect 4629 5661 4663 5695
rect 4813 5661 4847 5695
rect 5273 5661 5307 5695
rect 7757 5661 7791 5695
rect 8309 5661 8343 5695
rect 8493 5661 8527 5695
rect 3065 5593 3099 5627
rect 5549 5593 5583 5627
rect 1685 5525 1719 5559
rect 2697 5525 2731 5559
rect 7573 5525 7607 5559
rect 8493 5525 8527 5559
rect 3341 5321 3375 5355
rect 4905 5321 4939 5355
rect 5641 5321 5675 5355
rect 6653 5321 6687 5355
rect 10149 5321 10183 5355
rect 4169 5253 4203 5287
rect 4353 5253 4387 5287
rect 7849 5253 7883 5287
rect 9597 5253 9631 5287
rect 1777 5185 1811 5219
rect 2053 5185 2087 5219
rect 2513 5185 2547 5219
rect 2697 5185 2731 5219
rect 2881 5185 2915 5219
rect 3525 5185 3559 5219
rect 4997 5185 5031 5219
rect 5641 5185 5675 5219
rect 6561 5185 6595 5219
rect 6745 5185 6779 5219
rect 10057 5185 10091 5219
rect 1593 4981 1627 5015
rect 1961 4981 1995 5015
rect 3985 4981 4019 5015
rect 3249 4777 3283 4811
rect 3985 4777 4019 4811
rect 5549 4777 5583 4811
rect 9873 4777 9907 4811
rect 1685 4709 1719 4743
rect 2605 4709 2639 4743
rect 4721 4709 4755 4743
rect 2421 4641 2455 4675
rect 1869 4573 1903 4607
rect 2697 4573 2731 4607
rect 3341 4573 3375 4607
rect 4169 4573 4203 4607
rect 4813 4573 4847 4607
rect 5365 4573 5399 4607
rect 7665 4573 7699 4607
rect 9965 4573 9999 4607
rect 7757 4505 7791 4539
rect 2421 4437 2455 4471
rect 4077 4233 4111 4267
rect 7849 4165 7883 4199
rect 1869 4097 1903 4131
rect 2796 4097 2830 4131
rect 3525 4097 3559 4131
rect 3617 4097 3651 4131
rect 4629 4097 4663 4131
rect 4813 4097 4847 4131
rect 7573 4097 7607 4131
rect 2881 4029 2915 4063
rect 9321 4029 9355 4063
rect 1685 3893 1719 3927
rect 2421 3893 2455 3927
rect 4629 3893 4663 3927
rect 1869 3689 1903 3723
rect 2789 3689 2823 3723
rect 3985 3689 4019 3723
rect 4629 3689 4663 3723
rect 3341 3621 3375 3655
rect 2053 3485 2087 3519
rect 2605 3485 2639 3519
rect 2789 3485 2823 3519
rect 3433 3485 3467 3519
rect 3985 3485 4019 3519
rect 4169 3485 4203 3519
rect 3433 3145 3467 3179
rect 4077 3077 4111 3111
rect 1869 3009 1903 3043
rect 3525 3009 3559 3043
rect 3985 3009 4019 3043
rect 4169 3009 4203 3043
rect 1685 2805 1719 2839
rect 1593 2397 1627 2431
rect 1777 2261 1811 2295
<< metal1 >>
rect 4430 15852 4436 15904
rect 4488 15892 4494 15904
rect 13906 15892 13912 15904
rect 4488 15864 13912 15892
rect 4488 15852 4494 15864
rect 13906 15852 13912 15864
rect 13964 15852 13970 15904
rect 1104 15802 16836 15824
rect 1104 15750 2916 15802
rect 2968 15750 2980 15802
rect 3032 15750 3044 15802
rect 3096 15750 3108 15802
rect 3160 15750 3172 15802
rect 3224 15750 6849 15802
rect 6901 15750 6913 15802
rect 6965 15750 6977 15802
rect 7029 15750 7041 15802
rect 7093 15750 7105 15802
rect 7157 15750 10782 15802
rect 10834 15750 10846 15802
rect 10898 15750 10910 15802
rect 10962 15750 10974 15802
rect 11026 15750 11038 15802
rect 11090 15750 14715 15802
rect 14767 15750 14779 15802
rect 14831 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 16836 15802
rect 1104 15728 16836 15750
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 2832 15660 2877 15688
rect 2832 15648 2838 15660
rect 4154 15648 4160 15700
rect 4212 15688 4218 15700
rect 5077 15691 5135 15697
rect 5077 15688 5089 15691
rect 4212 15660 5089 15688
rect 4212 15648 4218 15660
rect 5077 15657 5089 15660
rect 5123 15657 5135 15691
rect 5077 15651 5135 15657
rect 2038 15620 2044 15632
rect 1999 15592 2044 15620
rect 2038 15580 2044 15592
rect 2096 15580 2102 15632
rect 4246 15620 4252 15632
rect 4207 15592 4252 15620
rect 4246 15580 4252 15592
rect 4304 15580 4310 15632
rect 4430 15620 4436 15632
rect 4391 15592 4436 15620
rect 4430 15580 4436 15592
rect 4488 15580 4494 15632
rect 5902 15580 5908 15632
rect 5960 15620 5966 15632
rect 5960 15592 13032 15620
rect 5960 15580 5966 15592
rect 2225 15555 2283 15561
rect 2225 15521 2237 15555
rect 2271 15552 2283 15555
rect 2271 15524 11928 15552
rect 2271 15521 2283 15524
rect 2225 15515 2283 15521
rect 2958 15484 2964 15496
rect 2919 15456 2964 15484
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 4893 15487 4951 15493
rect 4893 15484 4905 15487
rect 3804 15456 4905 15484
rect 1765 15419 1823 15425
rect 1765 15385 1777 15419
rect 1811 15385 1823 15419
rect 1765 15379 1823 15385
rect 1780 15348 1808 15379
rect 2406 15376 2412 15428
rect 2464 15416 2470 15428
rect 3804 15416 3832 15456
rect 4893 15453 4905 15456
rect 4939 15453 4951 15487
rect 4893 15447 4951 15453
rect 5534 15444 5540 15496
rect 5592 15484 5598 15496
rect 5902 15484 5908 15496
rect 5592 15456 5908 15484
rect 5592 15444 5598 15456
rect 5902 15444 5908 15456
rect 5960 15444 5966 15496
rect 8294 15444 8300 15496
rect 8352 15484 8358 15496
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 8352 15456 9137 15484
rect 8352 15444 8358 15456
rect 9125 15453 9137 15456
rect 9171 15453 9183 15487
rect 10318 15484 10324 15496
rect 10279 15456 10324 15484
rect 9125 15447 9183 15453
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 11057 15487 11115 15493
rect 11057 15453 11069 15487
rect 11103 15484 11115 15487
rect 11330 15484 11336 15496
rect 11103 15456 11336 15484
rect 11103 15453 11115 15456
rect 11057 15447 11115 15453
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 11900 15493 11928 15524
rect 11885 15487 11943 15493
rect 11885 15453 11897 15487
rect 11931 15453 11943 15487
rect 12526 15484 12532 15496
rect 12487 15456 12532 15484
rect 11885 15447 11943 15453
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 13004 15493 13032 15592
rect 13814 15512 13820 15564
rect 13872 15552 13878 15564
rect 14277 15555 14335 15561
rect 14277 15552 14289 15555
rect 13872 15524 14289 15552
rect 13872 15512 13878 15524
rect 14277 15521 14289 15524
rect 14323 15552 14335 15555
rect 15565 15555 15623 15561
rect 15565 15552 15577 15555
rect 14323 15524 15577 15552
rect 14323 15521 14335 15524
rect 14277 15515 14335 15521
rect 15565 15521 15577 15524
rect 15611 15521 15623 15555
rect 15565 15515 15623 15521
rect 12989 15487 13047 15493
rect 12989 15453 13001 15487
rect 13035 15453 13047 15487
rect 12989 15447 13047 15453
rect 13998 15444 14004 15496
rect 14056 15484 14062 15496
rect 14553 15487 14611 15493
rect 14553 15484 14565 15487
rect 14056 15456 14565 15484
rect 14056 15444 14062 15456
rect 14553 15453 14565 15456
rect 14599 15453 14611 15487
rect 14553 15447 14611 15453
rect 2464 15388 3832 15416
rect 3973 15419 4031 15425
rect 2464 15376 2470 15388
rect 3973 15385 3985 15419
rect 4019 15385 4031 15419
rect 3973 15379 4031 15385
rect 5997 15419 6055 15425
rect 5997 15385 6009 15419
rect 6043 15416 6055 15419
rect 6362 15416 6368 15428
rect 6043 15388 6368 15416
rect 6043 15385 6055 15388
rect 5997 15379 6055 15385
rect 3234 15348 3240 15360
rect 1780 15320 3240 15348
rect 3234 15308 3240 15320
rect 3292 15348 3298 15360
rect 3988 15348 4016 15379
rect 6362 15376 6368 15388
rect 6420 15376 6426 15428
rect 6546 15416 6552 15428
rect 6507 15388 6552 15416
rect 6546 15376 6552 15388
rect 6604 15376 6610 15428
rect 8662 15376 8668 15428
rect 8720 15416 8726 15428
rect 12437 15419 12495 15425
rect 12437 15416 12449 15419
rect 8720 15388 12449 15416
rect 8720 15376 8726 15388
rect 12437 15385 12449 15388
rect 12483 15385 12495 15419
rect 12437 15379 12495 15385
rect 7834 15348 7840 15360
rect 3292 15320 4016 15348
rect 7795 15320 7840 15348
rect 3292 15308 3298 15320
rect 7834 15308 7840 15320
rect 7892 15308 7898 15360
rect 9306 15348 9312 15360
rect 9267 15320 9312 15348
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 10226 15348 10232 15360
rect 10187 15320 10232 15348
rect 10226 15308 10232 15320
rect 10284 15308 10290 15360
rect 10962 15348 10968 15360
rect 10923 15320 10968 15348
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 11054 15308 11060 15360
rect 11112 15348 11118 15360
rect 11701 15351 11759 15357
rect 11701 15348 11713 15351
rect 11112 15320 11713 15348
rect 11112 15308 11118 15320
rect 11701 15317 11713 15320
rect 11747 15317 11759 15351
rect 11701 15311 11759 15317
rect 13081 15351 13139 15357
rect 13081 15317 13093 15351
rect 13127 15348 13139 15351
rect 13262 15348 13268 15360
rect 13127 15320 13268 15348
rect 13127 15317 13139 15320
rect 13081 15311 13139 15317
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 13725 15351 13783 15357
rect 13725 15317 13737 15351
rect 13771 15348 13783 15351
rect 13814 15348 13820 15360
rect 13771 15320 13820 15348
rect 13771 15317 13783 15320
rect 13725 15311 13783 15317
rect 13814 15308 13820 15320
rect 13872 15308 13878 15360
rect 1104 15258 16995 15280
rect 1104 15206 4882 15258
rect 4934 15206 4946 15258
rect 4998 15206 5010 15258
rect 5062 15206 5074 15258
rect 5126 15206 5138 15258
rect 5190 15206 8815 15258
rect 8867 15206 8879 15258
rect 8931 15206 8943 15258
rect 8995 15206 9007 15258
rect 9059 15206 9071 15258
rect 9123 15206 12748 15258
rect 12800 15206 12812 15258
rect 12864 15206 12876 15258
rect 12928 15206 12940 15258
rect 12992 15206 13004 15258
rect 13056 15206 16681 15258
rect 16733 15206 16745 15258
rect 16797 15206 16809 15258
rect 16861 15206 16873 15258
rect 16925 15206 16937 15258
rect 16989 15206 16995 15258
rect 1104 15184 16995 15206
rect 2038 15144 2044 15156
rect 1999 15116 2044 15144
rect 2038 15104 2044 15116
rect 2096 15104 2102 15156
rect 2406 15144 2412 15156
rect 2367 15116 2412 15144
rect 2406 15104 2412 15116
rect 2464 15104 2470 15156
rect 14369 15147 14427 15153
rect 14369 15144 14381 15147
rect 5000 15116 14381 15144
rect 5000 15017 5028 15116
rect 14369 15113 14381 15116
rect 14415 15113 14427 15147
rect 14369 15107 14427 15113
rect 6730 15076 6736 15088
rect 6012 15048 6736 15076
rect 6012 15017 6040 15048
rect 6730 15036 6736 15048
rect 6788 15036 6794 15088
rect 8662 15076 8668 15088
rect 8050 15048 8668 15076
rect 8662 15036 8668 15048
rect 8720 15036 8726 15088
rect 9306 15076 9312 15088
rect 8772 15048 9312 15076
rect 4729 15011 4787 15017
rect 4729 14977 4741 15011
rect 4775 15008 4787 15011
rect 4985 15011 5043 15017
rect 4775 14980 4936 15008
rect 4775 14977 4787 14980
rect 4729 14971 4787 14977
rect 2501 14943 2559 14949
rect 2501 14909 2513 14943
rect 2547 14909 2559 14943
rect 2501 14903 2559 14909
rect 2516 14872 2544 14903
rect 2590 14900 2596 14952
rect 2648 14940 2654 14952
rect 4908 14940 4936 14980
rect 4985 14977 4997 15011
rect 5031 14977 5043 15011
rect 4985 14971 5043 14977
rect 5997 15011 6055 15017
rect 5997 14977 6009 15011
rect 6043 14977 6055 15011
rect 5997 14971 6055 14977
rect 6362 14968 6368 15020
rect 6420 15008 6426 15020
rect 8772 15017 8800 15048
rect 9306 15036 9312 15048
rect 9364 15036 9370 15088
rect 10962 15076 10968 15088
rect 10258 15048 10968 15076
rect 10962 15036 10968 15048
rect 11020 15036 11026 15088
rect 11072 15048 12388 15076
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 6420 14980 6561 15008
rect 6420 14968 6426 14980
rect 6549 14977 6561 14980
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 8757 15011 8815 15017
rect 8757 14977 8769 15011
rect 8803 14977 8815 15011
rect 8757 14971 8815 14977
rect 10410 14968 10416 15020
rect 10468 15008 10474 15020
rect 11072 15008 11100 15048
rect 10468 14980 11100 15008
rect 11149 15011 11207 15017
rect 10468 14968 10474 14980
rect 11149 14977 11161 15011
rect 11195 15008 11207 15011
rect 11238 15008 11244 15020
rect 11195 14980 11244 15008
rect 11195 14977 11207 14980
rect 11149 14971 11207 14977
rect 11238 14968 11244 14980
rect 11296 14968 11302 15020
rect 11330 14968 11336 15020
rect 11388 15008 11394 15020
rect 12360 15017 12388 15048
rect 11885 15011 11943 15017
rect 11885 15008 11897 15011
rect 11388 14980 11897 15008
rect 11388 14968 11394 14980
rect 11885 14977 11897 14980
rect 11931 14977 11943 15011
rect 11885 14971 11943 14977
rect 12345 15011 12403 15017
rect 12345 14977 12357 15011
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 6454 14940 6460 14952
rect 2648 14912 2693 14940
rect 4908 14912 6460 14940
rect 2648 14900 2654 14912
rect 6454 14900 6460 14912
rect 6512 14900 6518 14952
rect 6825 14943 6883 14949
rect 6825 14909 6837 14943
rect 6871 14940 6883 14943
rect 8110 14940 8116 14952
rect 6871 14912 8116 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 8110 14900 8116 14912
rect 8168 14900 8174 14952
rect 8294 14940 8300 14952
rect 8255 14912 8300 14940
rect 8294 14900 8300 14912
rect 8352 14900 8358 14952
rect 9033 14943 9091 14949
rect 9033 14909 9045 14943
rect 9079 14940 9091 14943
rect 9582 14940 9588 14952
rect 9079 14912 9588 14940
rect 9079 14909 9091 14912
rect 9033 14903 9091 14909
rect 9582 14900 9588 14912
rect 9640 14900 9646 14952
rect 9766 14900 9772 14952
rect 9824 14940 9830 14952
rect 10318 14940 10324 14952
rect 9824 14912 10324 14940
rect 9824 14900 9830 14912
rect 10318 14900 10324 14912
rect 10376 14940 10382 14952
rect 10505 14943 10563 14949
rect 10505 14940 10517 14943
rect 10376 14912 10517 14940
rect 10376 14900 10382 14912
rect 10505 14909 10517 14912
rect 10551 14909 10563 14943
rect 11900 14940 11928 14971
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 13173 15011 13231 15017
rect 13173 15008 13185 15011
rect 12492 14980 13185 15008
rect 12492 14968 12498 14980
rect 13173 14977 13185 14980
rect 13219 14977 13231 15011
rect 13814 15008 13820 15020
rect 13727 14980 13820 15008
rect 13173 14971 13231 14977
rect 13814 14968 13820 14980
rect 13872 15008 13878 15020
rect 14461 15011 14519 15017
rect 14461 15008 14473 15011
rect 13872 14980 14473 15008
rect 13872 14968 13878 14980
rect 14461 14977 14473 14980
rect 14507 15008 14519 15011
rect 14507 14980 15056 15008
rect 14507 14977 14519 14980
rect 14461 14971 14519 14977
rect 12526 14940 12532 14952
rect 11900 14912 12532 14940
rect 10505 14903 10563 14909
rect 12526 14900 12532 14912
rect 12584 14940 12590 14952
rect 13078 14940 13084 14952
rect 12584 14912 13084 14940
rect 12584 14900 12590 14912
rect 13078 14900 13084 14912
rect 13136 14900 13142 14952
rect 13725 14875 13783 14881
rect 13725 14872 13737 14875
rect 2516 14844 2774 14872
rect 2746 14804 2774 14844
rect 5552 14844 6684 14872
rect 2958 14804 2964 14816
rect 2746 14776 2964 14804
rect 2958 14764 2964 14776
rect 3016 14804 3022 14816
rect 3602 14804 3608 14816
rect 3016 14776 3608 14804
rect 3016 14764 3022 14776
rect 3602 14764 3608 14776
rect 3660 14764 3666 14816
rect 3786 14764 3792 14816
rect 3844 14804 3850 14816
rect 5552 14804 5580 14844
rect 3844 14776 5580 14804
rect 3844 14764 3850 14776
rect 5626 14764 5632 14816
rect 5684 14804 5690 14816
rect 5905 14807 5963 14813
rect 5905 14804 5917 14807
rect 5684 14776 5917 14804
rect 5684 14764 5690 14776
rect 5905 14773 5917 14776
rect 5951 14773 5963 14807
rect 6656 14804 6684 14844
rect 8128 14844 8892 14872
rect 8128 14804 8156 14844
rect 6656 14776 8156 14804
rect 8864 14804 8892 14844
rect 10060 14844 13737 14872
rect 10060 14804 10088 14844
rect 13725 14841 13737 14844
rect 13771 14841 13783 14875
rect 13725 14835 13783 14841
rect 8864 14776 10088 14804
rect 5905 14767 5963 14773
rect 10134 14764 10140 14816
rect 10192 14804 10198 14816
rect 10962 14804 10968 14816
rect 10192 14776 10968 14804
rect 10192 14764 10198 14776
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 11057 14807 11115 14813
rect 11057 14773 11069 14807
rect 11103 14804 11115 14807
rect 11146 14804 11152 14816
rect 11103 14776 11152 14804
rect 11103 14773 11115 14776
rect 11057 14767 11115 14773
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 11790 14804 11796 14816
rect 11751 14776 11796 14804
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 12342 14764 12348 14816
rect 12400 14804 12406 14816
rect 12437 14807 12495 14813
rect 12437 14804 12449 14807
rect 12400 14776 12449 14804
rect 12400 14764 12406 14776
rect 12437 14773 12449 14776
rect 12483 14773 12495 14807
rect 12437 14767 12495 14773
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 15028 14813 15056 14980
rect 12989 14807 13047 14813
rect 12989 14804 13001 14807
rect 12676 14776 13001 14804
rect 12676 14764 12682 14776
rect 12989 14773 13001 14776
rect 13035 14773 13047 14807
rect 12989 14767 13047 14773
rect 15013 14807 15071 14813
rect 15013 14773 15025 14807
rect 15059 14804 15071 14807
rect 15102 14804 15108 14816
rect 15059 14776 15108 14804
rect 15059 14773 15071 14776
rect 15013 14767 15071 14773
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 1104 14714 16836 14736
rect 1104 14662 2916 14714
rect 2968 14662 2980 14714
rect 3032 14662 3044 14714
rect 3096 14662 3108 14714
rect 3160 14662 3172 14714
rect 3224 14662 6849 14714
rect 6901 14662 6913 14714
rect 6965 14662 6977 14714
rect 7029 14662 7041 14714
rect 7093 14662 7105 14714
rect 7157 14662 10782 14714
rect 10834 14662 10846 14714
rect 10898 14662 10910 14714
rect 10962 14662 10974 14714
rect 11026 14662 11038 14714
rect 11090 14662 14715 14714
rect 14767 14662 14779 14714
rect 14831 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 16836 14714
rect 1104 14640 16836 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 2314 14600 2320 14612
rect 1627 14572 2320 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 2314 14560 2320 14572
rect 2372 14560 2378 14612
rect 3973 14603 4031 14609
rect 3973 14569 3985 14603
rect 4019 14600 4031 14603
rect 4246 14600 4252 14612
rect 4019 14572 4252 14600
rect 4019 14569 4031 14572
rect 3973 14563 4031 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 8110 14600 8116 14612
rect 8071 14572 8116 14600
rect 8110 14560 8116 14572
rect 8168 14560 8174 14612
rect 9582 14600 9588 14612
rect 9543 14572 9588 14600
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 10492 14603 10550 14609
rect 10492 14569 10504 14603
rect 10538 14600 10550 14603
rect 11606 14600 11612 14612
rect 10538 14572 11612 14600
rect 10538 14569 10550 14572
rect 10492 14563 10550 14569
rect 11606 14560 11612 14572
rect 11664 14560 11670 14612
rect 10134 14532 10140 14544
rect 2976 14504 10140 14532
rect 2976 14464 3004 14504
rect 10134 14492 10140 14504
rect 10192 14492 10198 14544
rect 2884 14436 3004 14464
rect 4617 14467 4675 14473
rect 2705 14399 2763 14405
rect 2705 14365 2717 14399
rect 2751 14396 2763 14399
rect 2884 14396 2912 14436
rect 4617 14433 4629 14467
rect 4663 14464 4675 14467
rect 5810 14464 5816 14476
rect 4663 14436 5816 14464
rect 4663 14433 4675 14436
rect 4617 14427 4675 14433
rect 5810 14424 5816 14436
rect 5868 14424 5874 14476
rect 14369 14467 14427 14473
rect 14369 14464 14381 14467
rect 7852 14436 14381 14464
rect 2751 14368 2912 14396
rect 2961 14399 3019 14405
rect 2751 14365 2763 14368
rect 2705 14359 2763 14365
rect 2961 14365 2973 14399
rect 3007 14396 3019 14399
rect 7852 14396 7880 14436
rect 14369 14433 14381 14436
rect 14415 14433 14427 14467
rect 14369 14427 14427 14433
rect 8294 14396 8300 14408
rect 3007 14368 7880 14396
rect 8255 14368 8300 14396
rect 3007 14365 3019 14368
rect 2961 14359 3019 14365
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 9766 14396 9772 14408
rect 9727 14368 9772 14396
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 10226 14396 10232 14408
rect 10187 14368 10232 14396
rect 10226 14356 10232 14368
rect 10284 14356 10290 14408
rect 12621 14399 12679 14405
rect 12621 14396 12633 14399
rect 11900 14368 12633 14396
rect 3602 14288 3608 14340
rect 3660 14328 3666 14340
rect 4341 14331 4399 14337
rect 4341 14328 4353 14331
rect 3660 14300 4353 14328
rect 3660 14288 3666 14300
rect 4341 14297 4353 14300
rect 4387 14297 4399 14331
rect 4341 14291 4399 14297
rect 4706 14288 4712 14340
rect 4764 14328 4770 14340
rect 5261 14331 5319 14337
rect 5261 14328 5273 14331
rect 4764 14300 5273 14328
rect 4764 14288 4770 14300
rect 5261 14297 5273 14300
rect 5307 14328 5319 14331
rect 5442 14328 5448 14340
rect 5307 14300 5448 14328
rect 5307 14297 5319 14300
rect 5261 14291 5319 14297
rect 5442 14288 5448 14300
rect 5500 14288 5506 14340
rect 6454 14288 6460 14340
rect 6512 14328 6518 14340
rect 11790 14328 11796 14340
rect 6512 14300 10916 14328
rect 11730 14300 11796 14328
rect 6512 14288 6518 14300
rect 10888 14272 10916 14300
rect 11790 14288 11796 14300
rect 11848 14288 11854 14340
rect 3326 14220 3332 14272
rect 3384 14260 3390 14272
rect 4433 14263 4491 14269
rect 4433 14260 4445 14263
rect 3384 14232 4445 14260
rect 3384 14220 3390 14232
rect 4433 14229 4445 14232
rect 4479 14229 4491 14263
rect 6546 14260 6552 14272
rect 6507 14232 6552 14260
rect 4433 14223 4491 14229
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 7374 14220 7380 14272
rect 7432 14260 7438 14272
rect 10410 14260 10416 14272
rect 7432 14232 10416 14260
rect 7432 14220 7438 14232
rect 10410 14220 10416 14232
rect 10468 14220 10474 14272
rect 10870 14220 10876 14272
rect 10928 14220 10934 14272
rect 11238 14220 11244 14272
rect 11296 14260 11302 14272
rect 11900 14260 11928 14368
rect 12621 14365 12633 14368
rect 12667 14365 12679 14399
rect 13078 14396 13084 14408
rect 13039 14368 13084 14396
rect 12621 14359 12679 14365
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14396 14519 14399
rect 14507 14368 15056 14396
rect 14507 14365 14519 14368
rect 14461 14359 14519 14365
rect 11296 14232 11928 14260
rect 11296 14220 11302 14232
rect 11974 14220 11980 14272
rect 12032 14260 12038 14272
rect 12526 14260 12532 14272
rect 12032 14232 12077 14260
rect 12487 14232 12532 14260
rect 12032 14220 12038 14232
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 13170 14260 13176 14272
rect 13131 14232 13176 14260
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 15028 14269 15056 14368
rect 15013 14263 15071 14269
rect 15013 14229 15025 14263
rect 15059 14260 15071 14263
rect 15102 14260 15108 14272
rect 15059 14232 15108 14260
rect 15059 14229 15071 14232
rect 15013 14223 15071 14229
rect 15102 14220 15108 14232
rect 15160 14220 15166 14272
rect 1104 14170 16995 14192
rect 1104 14118 4882 14170
rect 4934 14118 4946 14170
rect 4998 14118 5010 14170
rect 5062 14118 5074 14170
rect 5126 14118 5138 14170
rect 5190 14118 8815 14170
rect 8867 14118 8879 14170
rect 8931 14118 8943 14170
rect 8995 14118 9007 14170
rect 9059 14118 9071 14170
rect 9123 14118 12748 14170
rect 12800 14118 12812 14170
rect 12864 14118 12876 14170
rect 12928 14118 12940 14170
rect 12992 14118 13004 14170
rect 13056 14118 16681 14170
rect 16733 14118 16745 14170
rect 16797 14118 16809 14170
rect 16861 14118 16873 14170
rect 16925 14118 16937 14170
rect 16989 14118 16995 14170
rect 1104 14096 16995 14118
rect 1670 14056 1676 14068
rect 1631 14028 1676 14056
rect 1670 14016 1676 14028
rect 1728 14016 1734 14068
rect 2409 14059 2467 14065
rect 2409 14025 2421 14059
rect 2455 14056 2467 14059
rect 2774 14056 2780 14068
rect 2455 14028 2780 14056
rect 2455 14025 2467 14028
rect 2409 14019 2467 14025
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13920 1915 13923
rect 2424 13920 2452 14019
rect 2774 14016 2780 14028
rect 2832 14056 2838 14068
rect 3326 14056 3332 14068
rect 2832 14028 3332 14056
rect 2832 14016 2838 14028
rect 3326 14016 3332 14028
rect 3384 14016 3390 14068
rect 4249 14059 4307 14065
rect 4249 14025 4261 14059
rect 4295 14056 4307 14059
rect 5350 14056 5356 14068
rect 4295 14028 5356 14056
rect 4295 14025 4307 14028
rect 4249 14019 4307 14025
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 5442 14016 5448 14068
rect 5500 14056 5506 14068
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 5500 14028 6561 14056
rect 5500 14016 5506 14028
rect 6549 14025 6561 14028
rect 6595 14025 6607 14059
rect 6549 14019 6607 14025
rect 6730 14016 6736 14068
rect 6788 14056 6794 14068
rect 8297 14059 8355 14065
rect 8297 14056 8309 14059
rect 6788 14028 8309 14056
rect 6788 14016 6794 14028
rect 8297 14025 8309 14028
rect 8343 14056 8355 14059
rect 11330 14056 11336 14068
rect 8343 14028 11336 14056
rect 8343 14025 8355 14028
rect 8297 14019 8355 14025
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 11606 14016 11612 14068
rect 11664 14056 11670 14068
rect 11793 14059 11851 14065
rect 11793 14056 11805 14059
rect 11664 14028 11805 14056
rect 11664 14016 11670 14028
rect 11793 14025 11805 14028
rect 11839 14025 11851 14059
rect 11793 14019 11851 14025
rect 11882 14016 11888 14068
rect 11940 14056 11946 14068
rect 14550 14056 14556 14068
rect 11940 14028 14556 14056
rect 11940 14016 11946 14028
rect 14550 14016 14556 14028
rect 14608 14016 14614 14068
rect 3544 13991 3602 13997
rect 3544 13957 3556 13991
rect 3590 13988 3602 13991
rect 4062 13988 4068 14000
rect 3590 13960 4068 13988
rect 3590 13957 3602 13960
rect 3544 13951 3602 13957
rect 4062 13948 4068 13960
rect 4120 13948 4126 14000
rect 13170 13988 13176 14000
rect 5290 13960 13176 13988
rect 13170 13948 13176 13960
rect 13228 13948 13234 14000
rect 3786 13920 3792 13932
rect 1903 13892 2452 13920
rect 3747 13892 3792 13920
rect 1903 13889 1915 13892
rect 1857 13883 1915 13889
rect 3786 13880 3792 13892
rect 3844 13880 3850 13932
rect 6086 13880 6092 13932
rect 6144 13920 6150 13932
rect 7374 13920 7380 13932
rect 6144 13892 7380 13920
rect 6144 13880 6150 13892
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 9585 13923 9643 13929
rect 9585 13889 9597 13923
rect 9631 13920 9643 13923
rect 9674 13920 9680 13932
rect 9631 13892 9680 13920
rect 9631 13889 9643 13892
rect 9585 13883 9643 13889
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 9766 13880 9772 13932
rect 9824 13920 9830 13932
rect 10229 13923 10287 13929
rect 10229 13920 10241 13923
rect 9824 13892 10241 13920
rect 9824 13880 9830 13892
rect 10229 13889 10241 13892
rect 10275 13920 10287 13923
rect 10873 13923 10931 13929
rect 10275 13892 10640 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 5721 13855 5779 13861
rect 5721 13821 5733 13855
rect 5767 13852 5779 13855
rect 5997 13855 6055 13861
rect 5767 13824 5948 13852
rect 5767 13821 5779 13824
rect 5721 13815 5779 13821
rect 5920 13784 5948 13824
rect 5997 13821 6009 13855
rect 6043 13852 6055 13855
rect 7834 13852 7840 13864
rect 6043 13824 7840 13852
rect 6043 13821 6055 13824
rect 5997 13815 6055 13821
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 10137 13855 10195 13861
rect 10137 13821 10149 13855
rect 10183 13852 10195 13855
rect 10318 13852 10324 13864
rect 10183 13824 10324 13852
rect 10183 13821 10195 13824
rect 10137 13815 10195 13821
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 10612 13784 10640 13892
rect 10873 13889 10885 13923
rect 10919 13920 10931 13923
rect 11238 13920 11244 13932
rect 10919 13892 11244 13920
rect 10919 13889 10931 13892
rect 10873 13883 10931 13889
rect 11238 13880 11244 13892
rect 11296 13880 11302 13932
rect 11790 13920 11796 13932
rect 11751 13892 11796 13920
rect 11790 13880 11796 13892
rect 11848 13880 11854 13932
rect 12710 13920 12716 13932
rect 12671 13892 12716 13920
rect 12710 13880 12716 13892
rect 12768 13880 12774 13932
rect 13630 13920 13636 13932
rect 13591 13892 13636 13920
rect 13630 13880 13636 13892
rect 13688 13880 13694 13932
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 10686 13812 10692 13864
rect 10744 13852 10750 13864
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 10744 13824 10793 13852
rect 10744 13812 10750 13824
rect 10781 13821 10793 13824
rect 10827 13821 10839 13855
rect 14200 13852 14228 13883
rect 10781 13815 10839 13821
rect 10888 13824 14228 13852
rect 10888 13784 10916 13824
rect 13262 13784 13268 13796
rect 5920 13756 10548 13784
rect 10612 13756 10916 13784
rect 10980 13756 13268 13784
rect 4614 13676 4620 13728
rect 4672 13716 4678 13728
rect 6086 13716 6092 13728
rect 4672 13688 6092 13716
rect 4672 13676 4678 13688
rect 6086 13676 6092 13688
rect 6144 13676 6150 13728
rect 6730 13676 6736 13728
rect 6788 13716 6794 13728
rect 7193 13719 7251 13725
rect 7193 13716 7205 13719
rect 6788 13688 7205 13716
rect 6788 13676 6794 13688
rect 7193 13685 7205 13688
rect 7239 13685 7251 13719
rect 7193 13679 7251 13685
rect 7742 13676 7748 13728
rect 7800 13716 7806 13728
rect 10410 13716 10416 13728
rect 7800 13688 10416 13716
rect 7800 13676 7806 13688
rect 10410 13676 10416 13688
rect 10468 13676 10474 13728
rect 10520 13716 10548 13756
rect 10980 13716 11008 13756
rect 13262 13744 13268 13756
rect 13320 13744 13326 13796
rect 10520 13688 11008 13716
rect 11054 13676 11060 13728
rect 11112 13716 11118 13728
rect 12342 13716 12348 13728
rect 11112 13688 12348 13716
rect 11112 13676 11118 13688
rect 12342 13676 12348 13688
rect 12400 13676 12406 13728
rect 12897 13719 12955 13725
rect 12897 13685 12909 13719
rect 12943 13716 12955 13719
rect 13078 13716 13084 13728
rect 12943 13688 13084 13716
rect 12943 13685 12955 13688
rect 12897 13679 12955 13685
rect 13078 13676 13084 13688
rect 13136 13676 13142 13728
rect 13170 13676 13176 13728
rect 13228 13716 13234 13728
rect 13541 13719 13599 13725
rect 13541 13716 13553 13719
rect 13228 13688 13553 13716
rect 13228 13676 13234 13688
rect 13541 13685 13553 13688
rect 13587 13685 13599 13719
rect 13541 13679 13599 13685
rect 13814 13676 13820 13728
rect 13872 13716 13878 13728
rect 14277 13719 14335 13725
rect 14277 13716 14289 13719
rect 13872 13688 14289 13716
rect 13872 13676 13878 13688
rect 14277 13685 14289 13688
rect 14323 13685 14335 13719
rect 14277 13679 14335 13685
rect 1104 13626 16836 13648
rect 1104 13574 2916 13626
rect 2968 13574 2980 13626
rect 3032 13574 3044 13626
rect 3096 13574 3108 13626
rect 3160 13574 3172 13626
rect 3224 13574 6849 13626
rect 6901 13574 6913 13626
rect 6965 13574 6977 13626
rect 7029 13574 7041 13626
rect 7093 13574 7105 13626
rect 7157 13574 10782 13626
rect 10834 13574 10846 13626
rect 10898 13574 10910 13626
rect 10962 13574 10974 13626
rect 11026 13574 11038 13626
rect 11090 13574 14715 13626
rect 14767 13574 14779 13626
rect 14831 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 16836 13626
rect 1104 13552 16836 13574
rect 4798 13472 4804 13524
rect 4856 13512 4862 13524
rect 10594 13512 10600 13524
rect 4856 13484 10600 13512
rect 4856 13472 4862 13484
rect 10594 13472 10600 13484
rect 10652 13472 10658 13524
rect 11054 13472 11060 13524
rect 11112 13512 11118 13524
rect 11790 13512 11796 13524
rect 11112 13484 11796 13512
rect 11112 13472 11118 13484
rect 11790 13472 11796 13484
rect 11848 13472 11854 13524
rect 14550 13472 14556 13524
rect 14608 13512 14614 13524
rect 14921 13515 14979 13521
rect 14921 13512 14933 13515
rect 14608 13484 14933 13512
rect 14608 13472 14614 13484
rect 14921 13481 14933 13484
rect 14967 13481 14979 13515
rect 14921 13475 14979 13481
rect 4614 13444 4620 13456
rect 4575 13416 4620 13444
rect 4614 13404 4620 13416
rect 4672 13404 4678 13456
rect 11146 13444 11152 13456
rect 8220 13416 11152 13444
rect 2314 13336 2320 13388
rect 2372 13376 2378 13388
rect 2590 13376 2596 13388
rect 2372 13348 2596 13376
rect 2372 13336 2378 13348
rect 2590 13336 2596 13348
rect 2648 13376 2654 13388
rect 5718 13376 5724 13388
rect 2648 13348 5724 13376
rect 2648 13336 2654 13348
rect 5718 13336 5724 13348
rect 5776 13336 5782 13388
rect 6365 13379 6423 13385
rect 6365 13345 6377 13379
rect 6411 13376 6423 13379
rect 7834 13376 7840 13388
rect 6411 13348 7840 13376
rect 6411 13345 6423 13348
rect 6365 13339 6423 13345
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 1857 13311 1915 13317
rect 1857 13277 1869 13311
rect 1903 13308 1915 13311
rect 2038 13308 2044 13320
rect 1903 13280 2044 13308
rect 1903 13277 1915 13280
rect 1857 13271 1915 13277
rect 2038 13268 2044 13280
rect 2096 13308 2102 13320
rect 2685 13311 2743 13317
rect 2685 13308 2697 13311
rect 2096 13280 2697 13308
rect 2096 13268 2102 13280
rect 2685 13277 2697 13280
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 2774 13268 2780 13320
rect 2832 13308 2838 13320
rect 2832 13280 2877 13308
rect 2832 13268 2838 13280
rect 3326 13268 3332 13320
rect 3384 13308 3390 13320
rect 3973 13311 4031 13317
rect 3973 13308 3985 13311
rect 3384 13280 3985 13308
rect 3384 13268 3390 13280
rect 3973 13277 3985 13280
rect 4019 13308 4031 13311
rect 4798 13308 4804 13320
rect 4019 13280 4804 13308
rect 4019 13277 4031 13280
rect 3973 13271 4031 13277
rect 4798 13268 4804 13280
rect 4856 13268 4862 13320
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 6825 13311 6883 13317
rect 6825 13308 6837 13311
rect 6788 13280 6837 13308
rect 6788 13268 6794 13280
rect 6825 13277 6837 13280
rect 6871 13277 6883 13311
rect 8220 13294 8248 13416
rect 11146 13404 11152 13416
rect 11204 13404 11210 13456
rect 12434 13376 12440 13388
rect 8404 13348 12440 13376
rect 6825 13271 6883 13277
rect 4065 13243 4123 13249
rect 4065 13209 4077 13243
rect 4111 13240 4123 13243
rect 4111 13212 4844 13240
rect 4111 13209 4123 13212
rect 4065 13203 4123 13209
rect 1670 13172 1676 13184
rect 1631 13144 1676 13172
rect 1670 13132 1676 13144
rect 1728 13132 1734 13184
rect 3142 13172 3148 13184
rect 3103 13144 3148 13172
rect 3142 13132 3148 13144
rect 3200 13132 3206 13184
rect 4816 13172 4844 13212
rect 5626 13200 5632 13252
rect 5684 13200 5690 13252
rect 6089 13243 6147 13249
rect 6089 13209 6101 13243
rect 6135 13240 6147 13243
rect 7098 13240 7104 13252
rect 6135 13212 6960 13240
rect 7059 13212 7104 13240
rect 6135 13209 6147 13212
rect 6089 13203 6147 13209
rect 6730 13172 6736 13184
rect 4816 13144 6736 13172
rect 6730 13132 6736 13144
rect 6788 13132 6794 13184
rect 6932 13172 6960 13212
rect 7098 13200 7104 13212
rect 7156 13200 7162 13252
rect 7742 13172 7748 13184
rect 6932 13144 7748 13172
rect 7742 13132 7748 13144
rect 7800 13132 7806 13184
rect 7834 13132 7840 13184
rect 7892 13172 7898 13184
rect 8404 13172 8432 13348
rect 12434 13336 12440 13348
rect 12492 13336 12498 13388
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 13964 13348 15148 13376
rect 13964 13336 13970 13348
rect 9125 13311 9183 13317
rect 9125 13308 9137 13311
rect 8680 13280 9137 13308
rect 7892 13144 8432 13172
rect 7892 13132 7898 13144
rect 8478 13132 8484 13184
rect 8536 13172 8542 13184
rect 8573 13175 8631 13181
rect 8573 13172 8585 13175
rect 8536 13144 8585 13172
rect 8536 13132 8542 13144
rect 8573 13141 8585 13144
rect 8619 13172 8631 13175
rect 8680 13172 8708 13280
rect 9125 13277 9137 13280
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 10689 13311 10747 13317
rect 10689 13277 10701 13311
rect 10735 13308 10747 13311
rect 10962 13308 10968 13320
rect 10735 13280 10968 13308
rect 10735 13277 10747 13280
rect 10689 13271 10747 13277
rect 10962 13268 10968 13280
rect 11020 13268 11026 13320
rect 11149 13311 11207 13317
rect 11149 13308 11161 13311
rect 11072 13280 11161 13308
rect 9306 13172 9312 13184
rect 8619 13144 8708 13172
rect 9267 13144 9312 13172
rect 8619 13141 8631 13144
rect 8573 13135 8631 13141
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 10505 13175 10563 13181
rect 10505 13141 10517 13175
rect 10551 13172 10563 13175
rect 11072 13172 11100 13280
rect 11149 13277 11161 13280
rect 11195 13277 11207 13311
rect 11149 13271 11207 13277
rect 12526 13268 12532 13320
rect 12584 13268 12590 13320
rect 13630 13308 13636 13320
rect 13591 13280 13636 13308
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 14458 13308 14464 13320
rect 14419 13280 14464 13308
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 15120 13317 15148 13348
rect 15105 13311 15163 13317
rect 15105 13277 15117 13311
rect 15151 13277 15163 13311
rect 15105 13271 15163 13277
rect 11422 13240 11428 13252
rect 11383 13212 11428 13240
rect 11422 13200 11428 13212
rect 11480 13200 11486 13252
rect 10551 13144 11100 13172
rect 10551 13141 10563 13144
rect 10505 13135 10563 13141
rect 12434 13132 12440 13184
rect 12492 13172 12498 13184
rect 12710 13172 12716 13184
rect 12492 13144 12716 13172
rect 12492 13132 12498 13144
rect 12710 13132 12716 13144
rect 12768 13172 12774 13184
rect 12897 13175 12955 13181
rect 12897 13172 12909 13175
rect 12768 13144 12909 13172
rect 12768 13132 12774 13144
rect 12897 13141 12909 13144
rect 12943 13141 12955 13175
rect 12897 13135 12955 13141
rect 13449 13175 13507 13181
rect 13449 13141 13461 13175
rect 13495 13172 13507 13175
rect 14182 13172 14188 13184
rect 13495 13144 14188 13172
rect 13495 13141 13507 13144
rect 13449 13135 13507 13141
rect 14182 13132 14188 13144
rect 14240 13132 14246 13184
rect 14274 13132 14280 13184
rect 14332 13172 14338 13184
rect 14369 13175 14427 13181
rect 14369 13172 14381 13175
rect 14332 13144 14381 13172
rect 14332 13132 14338 13144
rect 14369 13141 14381 13144
rect 14415 13141 14427 13175
rect 14369 13135 14427 13141
rect 1104 13082 16995 13104
rect 1104 13030 4882 13082
rect 4934 13030 4946 13082
rect 4998 13030 5010 13082
rect 5062 13030 5074 13082
rect 5126 13030 5138 13082
rect 5190 13030 8815 13082
rect 8867 13030 8879 13082
rect 8931 13030 8943 13082
rect 8995 13030 9007 13082
rect 9059 13030 9071 13082
rect 9123 13030 12748 13082
rect 12800 13030 12812 13082
rect 12864 13030 12876 13082
rect 12928 13030 12940 13082
rect 12992 13030 13004 13082
rect 13056 13030 16681 13082
rect 16733 13030 16745 13082
rect 16797 13030 16809 13082
rect 16861 13030 16873 13082
rect 16925 13030 16937 13082
rect 16989 13030 16995 13082
rect 1104 13008 16995 13030
rect 2133 12971 2191 12977
rect 2133 12937 2145 12971
rect 2179 12968 2191 12971
rect 2406 12968 2412 12980
rect 2179 12940 2412 12968
rect 2179 12937 2191 12940
rect 2133 12931 2191 12937
rect 2406 12928 2412 12940
rect 2464 12928 2470 12980
rect 13814 12968 13820 12980
rect 4448 12940 13820 12968
rect 2869 12903 2927 12909
rect 2869 12869 2881 12903
rect 2915 12900 2927 12903
rect 3234 12900 3240 12912
rect 2915 12872 3240 12900
rect 2915 12869 2927 12872
rect 2869 12863 2927 12869
rect 3234 12860 3240 12872
rect 3292 12860 3298 12912
rect 2038 12832 2044 12844
rect 1999 12804 2044 12832
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 4062 12832 4068 12844
rect 4023 12804 4068 12832
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 4448 12830 4476 12940
rect 13814 12928 13820 12940
rect 13872 12928 13878 12980
rect 14090 12928 14096 12980
rect 14148 12968 14154 12980
rect 15105 12971 15163 12977
rect 15105 12968 15117 12971
rect 14148 12940 15117 12968
rect 14148 12928 14154 12940
rect 15105 12937 15117 12940
rect 15151 12937 15163 12971
rect 15105 12931 15163 12937
rect 5810 12860 5816 12912
rect 5868 12900 5874 12912
rect 6549 12903 6607 12909
rect 6549 12900 6561 12903
rect 5868 12872 6561 12900
rect 5868 12860 5874 12872
rect 6549 12869 6561 12872
rect 6595 12869 6607 12903
rect 6549 12863 6607 12869
rect 7098 12860 7104 12912
rect 7156 12900 7162 12912
rect 8205 12903 8263 12909
rect 8205 12900 8217 12903
rect 7156 12872 8217 12900
rect 7156 12860 7162 12872
rect 8205 12869 8217 12872
rect 8251 12869 8263 12903
rect 9306 12900 9312 12912
rect 8205 12863 8263 12869
rect 9048 12872 9312 12900
rect 4798 12841 4804 12844
rect 4525 12835 4583 12841
rect 4525 12830 4537 12835
rect 4448 12802 4537 12830
rect 4525 12801 4537 12802
rect 4571 12801 4583 12835
rect 4792 12832 4804 12841
rect 4759 12804 4804 12832
rect 4525 12795 4583 12801
rect 4792 12795 4804 12804
rect 4798 12792 4804 12795
rect 4856 12792 4862 12844
rect 5074 12792 5080 12844
rect 5132 12832 5138 12844
rect 6641 12835 6699 12841
rect 6641 12832 6653 12835
rect 5132 12804 5856 12832
rect 5132 12792 5138 12804
rect 2314 12764 2320 12776
rect 2275 12736 2320 12764
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 3142 12696 3148 12708
rect 3103 12668 3148 12696
rect 3142 12656 3148 12668
rect 3200 12656 3206 12708
rect 3329 12699 3387 12705
rect 3329 12665 3341 12699
rect 3375 12696 3387 12699
rect 4522 12696 4528 12708
rect 3375 12668 4528 12696
rect 3375 12665 3387 12668
rect 3329 12659 3387 12665
rect 4522 12656 4528 12668
rect 4580 12656 4586 12708
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 3973 12631 4031 12637
rect 3973 12597 3985 12631
rect 4019 12628 4031 12631
rect 5626 12628 5632 12640
rect 4019 12600 5632 12628
rect 4019 12597 4031 12600
rect 3973 12591 4031 12597
rect 5626 12588 5632 12600
rect 5684 12588 5690 12640
rect 5828 12628 5856 12804
rect 5920 12804 6653 12832
rect 5920 12705 5948 12804
rect 6641 12801 6653 12804
rect 6687 12801 6699 12835
rect 6641 12795 6699 12801
rect 6730 12792 6736 12844
rect 6788 12832 6794 12844
rect 6917 12835 6975 12841
rect 6917 12832 6929 12835
rect 6788 12804 6929 12832
rect 6788 12792 6794 12804
rect 6917 12801 6929 12804
rect 6963 12801 6975 12835
rect 6917 12795 6975 12801
rect 7653 12835 7711 12841
rect 7653 12801 7665 12835
rect 7699 12832 7711 12835
rect 8018 12832 8024 12844
rect 7699 12804 8024 12832
rect 7699 12801 7711 12804
rect 7653 12795 7711 12801
rect 6932 12764 6960 12795
rect 8018 12792 8024 12804
rect 8076 12792 8082 12844
rect 8478 12832 8484 12844
rect 8439 12804 8484 12832
rect 8478 12792 8484 12804
rect 8536 12792 8542 12844
rect 9048 12841 9076 12872
rect 9306 12860 9312 12872
rect 9364 12860 9370 12912
rect 10686 12900 10692 12912
rect 10534 12872 10692 12900
rect 10686 12860 10692 12872
rect 10744 12860 10750 12912
rect 11422 12860 11428 12912
rect 11480 12900 11486 12912
rect 11977 12903 12035 12909
rect 11977 12900 11989 12903
rect 11480 12872 11989 12900
rect 11480 12860 11486 12872
rect 11977 12869 11989 12872
rect 12023 12869 12035 12903
rect 13078 12900 13084 12912
rect 11977 12863 12035 12869
rect 12912 12872 13084 12900
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12801 9091 12835
rect 9033 12795 9091 12801
rect 12253 12835 12311 12841
rect 12253 12801 12265 12835
rect 12299 12832 12311 12835
rect 12434 12832 12440 12844
rect 12299 12804 12440 12832
rect 12299 12801 12311 12804
rect 12253 12795 12311 12801
rect 12434 12792 12440 12804
rect 12492 12792 12498 12844
rect 12912 12841 12940 12872
rect 13078 12860 13084 12872
rect 13136 12860 13142 12912
rect 13170 12860 13176 12912
rect 13228 12900 13234 12912
rect 13228 12872 13273 12900
rect 13228 12860 13234 12872
rect 12897 12835 12955 12841
rect 12897 12801 12909 12835
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 14274 12792 14280 12844
rect 14332 12792 14338 12844
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12801 15347 12835
rect 15289 12795 15347 12801
rect 9309 12767 9367 12773
rect 9309 12764 9321 12767
rect 6932 12736 9321 12764
rect 9309 12733 9321 12736
rect 9355 12733 9367 12767
rect 9309 12727 9367 12733
rect 10594 12724 10600 12776
rect 10652 12764 10658 12776
rect 10781 12767 10839 12773
rect 10781 12764 10793 12767
rect 10652 12736 10793 12764
rect 10652 12724 10658 12736
rect 10781 12733 10793 12736
rect 10827 12733 10839 12767
rect 10781 12727 10839 12733
rect 13630 12724 13636 12776
rect 13688 12764 13694 12776
rect 14645 12767 14703 12773
rect 14645 12764 14657 12767
rect 13688 12736 14657 12764
rect 13688 12724 13694 12736
rect 14645 12733 14657 12736
rect 14691 12733 14703 12767
rect 14645 12727 14703 12733
rect 5905 12699 5963 12705
rect 5905 12665 5917 12699
rect 5951 12665 5963 12699
rect 15304 12696 15332 12795
rect 5905 12659 5963 12665
rect 7116 12668 7880 12696
rect 7116 12628 7144 12668
rect 5828 12600 7144 12628
rect 7190 12588 7196 12640
rect 7248 12628 7254 12640
rect 7469 12631 7527 12637
rect 7469 12628 7481 12631
rect 7248 12600 7481 12628
rect 7248 12588 7254 12600
rect 7469 12597 7481 12600
rect 7515 12597 7527 12631
rect 7852 12628 7880 12668
rect 14200 12668 15332 12696
rect 14200 12628 14228 12668
rect 7852 12600 14228 12628
rect 7469 12591 7527 12597
rect 1104 12538 16836 12560
rect 1104 12486 2916 12538
rect 2968 12486 2980 12538
rect 3032 12486 3044 12538
rect 3096 12486 3108 12538
rect 3160 12486 3172 12538
rect 3224 12486 6849 12538
rect 6901 12486 6913 12538
rect 6965 12486 6977 12538
rect 7029 12486 7041 12538
rect 7093 12486 7105 12538
rect 7157 12486 10782 12538
rect 10834 12486 10846 12538
rect 10898 12486 10910 12538
rect 10962 12486 10974 12538
rect 11026 12486 11038 12538
rect 11090 12486 14715 12538
rect 14767 12486 14779 12538
rect 14831 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 16836 12538
rect 1104 12464 16836 12486
rect 1673 12427 1731 12433
rect 1673 12393 1685 12427
rect 1719 12424 1731 12427
rect 2038 12424 2044 12436
rect 1719 12396 2044 12424
rect 1719 12393 1731 12396
rect 1673 12387 1731 12393
rect 2038 12384 2044 12396
rect 2096 12384 2102 12436
rect 15013 12427 15071 12433
rect 15013 12424 15025 12427
rect 3068 12396 15025 12424
rect 3068 12297 3096 12396
rect 15013 12393 15025 12396
rect 15059 12393 15071 12427
rect 15013 12387 15071 12393
rect 11517 12359 11575 12365
rect 11517 12325 11529 12359
rect 11563 12356 11575 12359
rect 12526 12356 12532 12368
rect 11563 12328 12532 12356
rect 11563 12325 11575 12328
rect 11517 12319 11575 12325
rect 12526 12316 12532 12328
rect 12584 12316 12590 12368
rect 3053 12291 3111 12297
rect 3053 12257 3065 12291
rect 3099 12257 3111 12291
rect 3053 12251 3111 12257
rect 5828 12260 12434 12288
rect 5828 12229 5856 12260
rect 5813 12223 5871 12229
rect 5813 12189 5825 12223
rect 5859 12189 5871 12223
rect 5813 12183 5871 12189
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 6273 12223 6331 12229
rect 6273 12220 6285 12223
rect 5960 12192 6285 12220
rect 5960 12180 5966 12192
rect 6273 12189 6285 12192
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 10594 12180 10600 12232
rect 10652 12220 10658 12232
rect 11333 12223 11391 12229
rect 11333 12220 11345 12223
rect 10652 12192 11345 12220
rect 10652 12180 10658 12192
rect 11333 12189 11345 12192
rect 11379 12189 11391 12223
rect 11333 12183 11391 12189
rect 12161 12223 12219 12229
rect 12161 12189 12173 12223
rect 12207 12189 12219 12223
rect 12161 12183 12219 12189
rect 2808 12155 2866 12161
rect 2808 12121 2820 12155
rect 2854 12152 2866 12155
rect 3234 12152 3240 12164
rect 2854 12124 3240 12152
rect 2854 12121 2866 12124
rect 2808 12115 2866 12121
rect 3234 12112 3240 12124
rect 3292 12112 3298 12164
rect 4246 12152 4252 12164
rect 4207 12124 4252 12152
rect 4246 12112 4252 12124
rect 4304 12112 4310 12164
rect 6549 12155 6607 12161
rect 6549 12121 6561 12155
rect 6595 12121 6607 12155
rect 6549 12115 6607 12121
rect 6564 12084 6592 12115
rect 7282 12112 7288 12164
rect 7340 12112 7346 12164
rect 10226 12112 10232 12164
rect 10284 12152 10290 12164
rect 10873 12155 10931 12161
rect 10873 12152 10885 12155
rect 10284 12124 10885 12152
rect 10284 12112 10290 12124
rect 10873 12121 10885 12124
rect 10919 12121 10931 12155
rect 10873 12115 10931 12121
rect 11238 12112 11244 12164
rect 11296 12152 11302 12164
rect 12176 12152 12204 12183
rect 11296 12124 12204 12152
rect 12406 12152 12434 12260
rect 13173 12223 13231 12229
rect 13173 12189 13185 12223
rect 13219 12220 13231 12223
rect 13354 12220 13360 12232
rect 13219 12192 13360 12220
rect 13219 12189 13231 12192
rect 13173 12183 13231 12189
rect 13354 12180 13360 12192
rect 13412 12180 13418 12232
rect 14458 12220 14464 12232
rect 14419 12192 14464 12220
rect 14458 12180 14464 12192
rect 14516 12180 14522 12232
rect 15102 12220 15108 12232
rect 15063 12192 15108 12220
rect 15102 12180 15108 12192
rect 15160 12220 15166 12232
rect 15565 12223 15623 12229
rect 15565 12220 15577 12223
rect 15160 12192 15577 12220
rect 15160 12180 15166 12192
rect 15565 12189 15577 12192
rect 15611 12189 15623 12223
rect 15565 12183 15623 12189
rect 12618 12152 12624 12164
rect 12406 12124 12624 12152
rect 11296 12112 11302 12124
rect 12618 12112 12624 12124
rect 12676 12112 12682 12164
rect 7190 12084 7196 12096
rect 6564 12056 7196 12084
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 8018 12084 8024 12096
rect 7979 12056 8024 12084
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 9585 12087 9643 12093
rect 9585 12053 9597 12087
rect 9631 12084 9643 12087
rect 9674 12084 9680 12096
rect 9631 12056 9680 12084
rect 9631 12053 9643 12056
rect 9585 12047 9643 12053
rect 9674 12044 9680 12056
rect 9732 12044 9738 12096
rect 12161 12087 12219 12093
rect 12161 12053 12173 12087
rect 12207 12084 12219 12087
rect 12434 12084 12440 12096
rect 12207 12056 12440 12084
rect 12207 12053 12219 12056
rect 12161 12047 12219 12053
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 12989 12087 13047 12093
rect 12989 12053 13001 12087
rect 13035 12084 13047 12087
rect 13906 12084 13912 12096
rect 13035 12056 13912 12084
rect 13035 12053 13047 12056
rect 12989 12047 13047 12053
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 14366 12084 14372 12096
rect 14327 12056 14372 12084
rect 14366 12044 14372 12056
rect 14424 12044 14430 12096
rect 1104 11994 16995 12016
rect 1104 11942 4882 11994
rect 4934 11942 4946 11994
rect 4998 11942 5010 11994
rect 5062 11942 5074 11994
rect 5126 11942 5138 11994
rect 5190 11942 8815 11994
rect 8867 11942 8879 11994
rect 8931 11942 8943 11994
rect 8995 11942 9007 11994
rect 9059 11942 9071 11994
rect 9123 11942 12748 11994
rect 12800 11942 12812 11994
rect 12864 11942 12876 11994
rect 12928 11942 12940 11994
rect 12992 11942 13004 11994
rect 13056 11942 16681 11994
rect 16733 11942 16745 11994
rect 16797 11942 16809 11994
rect 16861 11942 16873 11994
rect 16925 11942 16937 11994
rect 16989 11942 16995 11994
rect 1104 11920 16995 11942
rect 5258 11880 5264 11892
rect 2976 11852 5264 11880
rect 1581 11815 1639 11821
rect 1581 11781 1593 11815
rect 1627 11812 1639 11815
rect 1670 11812 1676 11824
rect 1627 11784 1676 11812
rect 1627 11781 1639 11784
rect 1581 11775 1639 11781
rect 1670 11772 1676 11784
rect 1728 11772 1734 11824
rect 2976 11753 3004 11852
rect 5258 11840 5264 11852
rect 5316 11840 5322 11892
rect 5902 11880 5908 11892
rect 5863 11852 5908 11880
rect 5902 11840 5908 11852
rect 5960 11840 5966 11892
rect 6733 11883 6791 11889
rect 6733 11849 6745 11883
rect 6779 11849 6791 11883
rect 7282 11880 7288 11892
rect 7243 11852 7288 11880
rect 6733 11843 6791 11849
rect 4430 11772 4436 11824
rect 4488 11772 4494 11824
rect 6748 11812 6776 11843
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 8110 11840 8116 11892
rect 8168 11880 8174 11892
rect 8205 11883 8263 11889
rect 8205 11880 8217 11883
rect 8168 11852 8217 11880
rect 8168 11840 8174 11852
rect 8205 11849 8217 11852
rect 8251 11849 8263 11883
rect 8205 11843 8263 11849
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 16117 11883 16175 11889
rect 16117 11880 16129 11883
rect 13412 11852 16129 11880
rect 13412 11840 13418 11852
rect 16117 11849 16129 11852
rect 16163 11849 16175 11883
rect 16117 11843 16175 11849
rect 12161 11815 12219 11821
rect 12161 11812 12173 11815
rect 6748 11784 12173 11812
rect 12161 11781 12173 11784
rect 12207 11781 12219 11815
rect 13998 11812 14004 11824
rect 12161 11775 12219 11781
rect 12406 11784 14004 11812
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11744 1823 11747
rect 2961 11747 3019 11753
rect 1811 11716 2636 11744
rect 1811 11713 1823 11716
rect 1765 11707 1823 11713
rect 1949 11543 2007 11549
rect 1949 11509 1961 11543
rect 1995 11540 2007 11543
rect 2130 11540 2136 11552
rect 1995 11512 2136 11540
rect 1995 11509 2007 11512
rect 1949 11503 2007 11509
rect 2130 11500 2136 11512
rect 2188 11500 2194 11552
rect 2608 11540 2636 11716
rect 2961 11713 2973 11747
rect 3007 11713 3019 11747
rect 5813 11747 5871 11753
rect 5813 11744 5825 11747
rect 2961 11707 3019 11713
rect 5644 11716 5825 11744
rect 2682 11636 2688 11688
rect 2740 11676 2746 11688
rect 3421 11679 3479 11685
rect 3421 11676 3433 11679
rect 2740 11648 3433 11676
rect 2740 11636 2746 11648
rect 3421 11645 3433 11648
rect 3467 11645 3479 11679
rect 3697 11679 3755 11685
rect 3697 11676 3709 11679
rect 3421 11639 3479 11645
rect 3528 11648 3709 11676
rect 2961 11611 3019 11617
rect 2961 11577 2973 11611
rect 3007 11608 3019 11611
rect 3528 11608 3556 11648
rect 3697 11645 3709 11648
rect 3743 11645 3755 11679
rect 3697 11639 3755 11645
rect 4062 11636 4068 11688
rect 4120 11676 4126 11688
rect 5644 11676 5672 11716
rect 5813 11713 5825 11716
rect 5859 11713 5871 11747
rect 5813 11707 5871 11713
rect 5902 11704 5908 11756
rect 5960 11744 5966 11756
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 5960 11716 6561 11744
rect 5960 11704 5966 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 7285 11747 7343 11753
rect 7285 11713 7297 11747
rect 7331 11744 7343 11747
rect 7469 11747 7527 11753
rect 7331 11716 7420 11744
rect 7331 11713 7343 11716
rect 7285 11707 7343 11713
rect 4120 11648 5672 11676
rect 4120 11636 4126 11648
rect 5644 11608 5672 11648
rect 6730 11608 6736 11620
rect 3007 11580 3556 11608
rect 5092 11580 5396 11608
rect 5644 11580 6736 11608
rect 3007 11577 3019 11580
rect 2961 11571 3019 11577
rect 3142 11540 3148 11552
rect 2608 11512 3148 11540
rect 3142 11500 3148 11512
rect 3200 11540 3206 11552
rect 5092 11540 5120 11580
rect 3200 11512 5120 11540
rect 5169 11543 5227 11549
rect 3200 11500 3206 11512
rect 5169 11509 5181 11543
rect 5215 11540 5227 11543
rect 5258 11540 5264 11552
rect 5215 11512 5264 11540
rect 5215 11509 5227 11512
rect 5169 11503 5227 11509
rect 5258 11500 5264 11512
rect 5316 11500 5322 11552
rect 5368 11540 5396 11580
rect 6730 11568 6736 11580
rect 6788 11568 6794 11620
rect 7392 11608 7420 11716
rect 7469 11713 7481 11747
rect 7515 11713 7527 11747
rect 7469 11707 7527 11713
rect 7484 11676 7512 11707
rect 7650 11704 7656 11756
rect 7708 11744 7714 11756
rect 8018 11744 8024 11756
rect 7708 11716 8024 11744
rect 7708 11704 7714 11716
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 9214 11744 9220 11756
rect 9175 11716 9220 11744
rect 9214 11704 9220 11716
rect 9272 11704 9278 11756
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 12406 11744 12434 11784
rect 13998 11772 14004 11784
rect 14056 11772 14062 11824
rect 14366 11772 14372 11824
rect 14424 11812 14430 11824
rect 14424 11784 15134 11812
rect 14424 11772 14430 11784
rect 9640 11716 12434 11744
rect 9640 11704 9646 11716
rect 9490 11676 9496 11688
rect 7484 11648 9496 11676
rect 9490 11636 9496 11648
rect 9548 11636 9554 11688
rect 14182 11636 14188 11688
rect 14240 11676 14246 11688
rect 14369 11679 14427 11685
rect 14369 11676 14381 11679
rect 14240 11648 14381 11676
rect 14240 11636 14246 11648
rect 14369 11645 14381 11648
rect 14415 11645 14427 11679
rect 14645 11679 14703 11685
rect 14645 11676 14657 11679
rect 14369 11639 14427 11645
rect 14476 11648 14657 11676
rect 8294 11608 8300 11620
rect 7392 11580 8300 11608
rect 8294 11568 8300 11580
rect 8352 11568 8358 11620
rect 13262 11568 13268 11620
rect 13320 11608 13326 11620
rect 14476 11608 14504 11648
rect 14645 11645 14657 11648
rect 14691 11645 14703 11679
rect 14645 11639 14703 11645
rect 13320 11580 14504 11608
rect 13320 11568 13326 11580
rect 9582 11540 9588 11552
rect 5368 11512 9588 11540
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 10410 11500 10416 11552
rect 10468 11540 10474 11552
rect 10505 11543 10563 11549
rect 10505 11540 10517 11543
rect 10468 11512 10517 11540
rect 10468 11500 10474 11512
rect 10505 11509 10517 11512
rect 10551 11509 10563 11543
rect 13630 11540 13636 11552
rect 13591 11512 13636 11540
rect 10505 11503 10563 11509
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 1104 11450 16836 11472
rect 1104 11398 2916 11450
rect 2968 11398 2980 11450
rect 3032 11398 3044 11450
rect 3096 11398 3108 11450
rect 3160 11398 3172 11450
rect 3224 11398 6849 11450
rect 6901 11398 6913 11450
rect 6965 11398 6977 11450
rect 7029 11398 7041 11450
rect 7093 11398 7105 11450
rect 7157 11398 10782 11450
rect 10834 11398 10846 11450
rect 10898 11398 10910 11450
rect 10962 11398 10974 11450
rect 11026 11398 11038 11450
rect 11090 11398 14715 11450
rect 14767 11398 14779 11450
rect 14831 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 16836 11450
rect 1104 11376 16836 11398
rect 2682 11336 2688 11348
rect 2643 11308 2688 11336
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 5626 11345 5632 11348
rect 5616 11339 5632 11345
rect 5616 11336 5628 11339
rect 5539 11308 5628 11336
rect 5616 11305 5628 11308
rect 5684 11336 5690 11348
rect 9214 11336 9220 11348
rect 5684 11308 8156 11336
rect 9175 11308 9220 11336
rect 5616 11299 5632 11305
rect 5626 11296 5632 11299
rect 5684 11296 5690 11308
rect 1670 11268 1676 11280
rect 1631 11240 1676 11268
rect 1670 11228 1676 11240
rect 1728 11228 1734 11280
rect 4430 11228 4436 11280
rect 4488 11268 4494 11280
rect 4525 11271 4583 11277
rect 4525 11268 4537 11271
rect 4488 11240 4537 11268
rect 4488 11228 4494 11240
rect 4525 11237 4537 11240
rect 4571 11237 4583 11271
rect 4525 11231 4583 11237
rect 6730 11228 6736 11280
rect 6788 11268 6794 11280
rect 7101 11271 7159 11277
rect 7101 11268 7113 11271
rect 6788 11240 7113 11268
rect 6788 11228 6794 11240
rect 7101 11237 7113 11240
rect 7147 11268 7159 11271
rect 7282 11268 7288 11280
rect 7147 11240 7288 11268
rect 7147 11237 7159 11240
rect 7101 11231 7159 11237
rect 7282 11228 7288 11240
rect 7340 11228 7346 11280
rect 3326 11200 3332 11212
rect 1872 11172 3332 11200
rect 1872 11141 1900 11172
rect 3326 11160 3332 11172
rect 3384 11160 3390 11212
rect 3421 11203 3479 11209
rect 3421 11169 3433 11203
rect 3467 11200 3479 11203
rect 6270 11200 6276 11212
rect 3467 11172 6276 11200
rect 3467 11169 3479 11172
rect 3421 11163 3479 11169
rect 6270 11160 6276 11172
rect 6328 11160 6334 11212
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11101 1915 11135
rect 1857 11095 1915 11101
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 4249 11135 4307 11141
rect 3283 11104 4200 11132
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 2700 11064 2728 11095
rect 4062 11064 4068 11076
rect 2700 11036 4068 11064
rect 4062 11024 4068 11036
rect 4120 11024 4126 11076
rect 4172 10996 4200 11104
rect 4249 11101 4261 11135
rect 4295 11101 4307 11135
rect 4249 11095 4307 11101
rect 4264 11064 4292 11095
rect 4338 11092 4344 11144
rect 4396 11132 4402 11144
rect 4433 11135 4491 11141
rect 4433 11132 4445 11135
rect 4396 11104 4445 11132
rect 4396 11092 4402 11104
rect 4433 11101 4445 11104
rect 4479 11101 4491 11135
rect 5342 11135 5400 11141
rect 5342 11132 5354 11135
rect 4433 11095 4491 11101
rect 4632 11104 5354 11132
rect 4632 11076 4660 11104
rect 5342 11101 5354 11104
rect 5388 11101 5400 11135
rect 5342 11095 5400 11101
rect 7650 11092 7656 11144
rect 7708 11132 7714 11144
rect 8128 11141 8156 11308
rect 9214 11296 9220 11308
rect 9272 11296 9278 11348
rect 10226 11336 10232 11348
rect 10187 11308 10232 11336
rect 10226 11296 10232 11308
rect 10284 11296 10290 11348
rect 13446 11336 13452 11348
rect 11440 11308 13452 11336
rect 8389 11271 8447 11277
rect 8389 11237 8401 11271
rect 8435 11268 8447 11271
rect 11440 11268 11468 11308
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 13262 11268 13268 11280
rect 8435 11240 11468 11268
rect 13223 11240 13268 11268
rect 8435 11237 8447 11240
rect 8389 11231 8447 11237
rect 13262 11228 13268 11240
rect 13320 11228 13326 11280
rect 13372 11240 13676 11268
rect 9766 11200 9772 11212
rect 9416 11172 9772 11200
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 7708 11104 8033 11132
rect 7708 11092 7714 11104
rect 8021 11101 8033 11104
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11101 8171 11135
rect 8113 11095 8171 11101
rect 9306 11092 9312 11144
rect 9364 11132 9370 11144
rect 9416 11141 9444 11172
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 10689 11203 10747 11209
rect 10689 11169 10701 11203
rect 10735 11200 10747 11203
rect 11238 11200 11244 11212
rect 10735 11172 11244 11200
rect 10735 11169 10747 11172
rect 10689 11163 10747 11169
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 11422 11160 11428 11212
rect 11480 11200 11486 11212
rect 13372 11200 13400 11240
rect 11480 11172 13400 11200
rect 13648 11200 13676 11240
rect 14458 11228 14464 11280
rect 14516 11268 14522 11280
rect 14516 11240 15424 11268
rect 14516 11228 14522 11240
rect 13648 11172 14964 11200
rect 11480 11160 11486 11172
rect 9401 11135 9459 11141
rect 9401 11132 9413 11135
rect 9364 11104 9413 11132
rect 9364 11092 9370 11104
rect 9401 11101 9413 11104
rect 9447 11101 9459 11135
rect 9582 11132 9588 11144
rect 9543 11104 9588 11132
rect 9401 11095 9459 11101
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11132 10103 11135
rect 11146 11132 11152 11144
rect 10091 11104 11152 11132
rect 10091 11101 10103 11104
rect 10045 11095 10103 11101
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 12710 11092 12716 11144
rect 12768 11132 12774 11144
rect 13354 11132 13360 11144
rect 12768 11104 12813 11132
rect 13315 11104 13360 11132
rect 12768 11092 12774 11104
rect 13354 11092 13360 11104
rect 13412 11092 13418 11144
rect 13446 11092 13452 11144
rect 13504 11132 13510 11144
rect 14936 11141 14964 11172
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 13504 11104 14473 11132
rect 13504 11092 13510 11104
rect 14461 11101 14473 11104
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11101 14979 11135
rect 15396 11132 15424 11240
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15396 11104 15761 11132
rect 14921 11095 14979 11101
rect 15749 11101 15761 11104
rect 15795 11132 15807 11135
rect 16114 11132 16120 11144
rect 15795 11104 16120 11132
rect 15795 11101 15807 11104
rect 15749 11095 15807 11101
rect 16114 11092 16120 11104
rect 16172 11092 16178 11144
rect 4614 11064 4620 11076
rect 4264 11036 4620 11064
rect 4614 11024 4620 11036
rect 4672 11024 4678 11076
rect 6362 11024 6368 11076
rect 6420 11024 6426 11076
rect 7837 11067 7895 11073
rect 7837 11033 7849 11067
rect 7883 11033 7895 11067
rect 7837 11027 7895 11033
rect 4522 10996 4528 11008
rect 4172 10968 4528 10996
rect 4522 10956 4528 10968
rect 4580 10956 4586 11008
rect 7742 10956 7748 11008
rect 7800 10996 7806 11008
rect 7852 10996 7880 11027
rect 7926 11024 7932 11076
rect 7984 11064 7990 11076
rect 8205 11067 8263 11073
rect 8205 11064 8217 11067
rect 7984 11036 8217 11064
rect 7984 11024 7990 11036
rect 8205 11033 8217 11036
rect 8251 11033 8263 11067
rect 12006 11036 12388 11064
rect 8205 11027 8263 11033
rect 11054 10996 11060 11008
rect 7800 10968 11060 10996
rect 7800 10956 7806 10968
rect 11054 10956 11060 10968
rect 11112 10956 11118 11008
rect 12360 10996 12388 11036
rect 12434 11024 12440 11076
rect 12492 11064 12498 11076
rect 15013 11067 15071 11073
rect 15013 11064 15025 11067
rect 12492 11036 12537 11064
rect 12636 11036 15025 11064
rect 12492 11024 12498 11036
rect 12636 10996 12664 11036
rect 15013 11033 15025 11036
rect 15059 11033 15071 11067
rect 15654 11064 15660 11076
rect 15615 11036 15660 11064
rect 15013 11027 15071 11033
rect 15654 11024 15660 11036
rect 15712 11024 15718 11076
rect 12360 10968 12664 10996
rect 13814 10956 13820 11008
rect 13872 10996 13878 11008
rect 14277 10999 14335 11005
rect 14277 10996 14289 10999
rect 13872 10968 14289 10996
rect 13872 10956 13878 10968
rect 14277 10965 14289 10968
rect 14323 10965 14335 10999
rect 14277 10959 14335 10965
rect 1104 10906 16995 10928
rect 1104 10854 4882 10906
rect 4934 10854 4946 10906
rect 4998 10854 5010 10906
rect 5062 10854 5074 10906
rect 5126 10854 5138 10906
rect 5190 10854 8815 10906
rect 8867 10854 8879 10906
rect 8931 10854 8943 10906
rect 8995 10854 9007 10906
rect 9059 10854 9071 10906
rect 9123 10854 12748 10906
rect 12800 10854 12812 10906
rect 12864 10854 12876 10906
rect 12928 10854 12940 10906
rect 12992 10854 13004 10906
rect 13056 10854 16681 10906
rect 16733 10854 16745 10906
rect 16797 10854 16809 10906
rect 16861 10854 16873 10906
rect 16925 10854 16937 10906
rect 16989 10854 16995 10906
rect 1104 10832 16995 10854
rect 2501 10795 2559 10801
rect 2501 10761 2513 10795
rect 2547 10792 2559 10795
rect 4062 10792 4068 10804
rect 2547 10764 4068 10792
rect 2547 10761 2559 10764
rect 2501 10755 2559 10761
rect 4062 10752 4068 10764
rect 4120 10752 4126 10804
rect 7834 10792 7840 10804
rect 7795 10764 7840 10792
rect 7834 10752 7840 10764
rect 7892 10752 7898 10804
rect 10318 10752 10324 10804
rect 10376 10752 10382 10804
rect 3789 10727 3847 10733
rect 3789 10693 3801 10727
rect 3835 10724 3847 10727
rect 4246 10724 4252 10736
rect 3835 10696 4252 10724
rect 3835 10693 3847 10696
rect 3789 10687 3847 10693
rect 4246 10684 4252 10696
rect 4304 10684 4310 10736
rect 6546 10724 6552 10736
rect 6507 10696 6552 10724
rect 6546 10684 6552 10696
rect 6604 10684 6610 10736
rect 10336 10665 10364 10752
rect 10410 10684 10416 10736
rect 10468 10724 10474 10736
rect 11701 10727 11759 10733
rect 11701 10724 11713 10727
rect 10468 10696 11713 10724
rect 10468 10684 10474 10696
rect 11701 10693 11713 10696
rect 11747 10693 11759 10727
rect 15654 10724 15660 10736
rect 15410 10696 15660 10724
rect 11701 10687 11759 10693
rect 15654 10684 15660 10696
rect 15712 10684 15718 10736
rect 10065 10659 10123 10665
rect 10065 10625 10077 10659
rect 10111 10656 10123 10659
rect 10321 10659 10379 10665
rect 10111 10628 10272 10656
rect 10111 10625 10123 10628
rect 10065 10619 10123 10625
rect 5997 10591 6055 10597
rect 5997 10557 6009 10591
rect 6043 10588 6055 10591
rect 9306 10588 9312 10600
rect 6043 10560 9312 10588
rect 6043 10557 6055 10560
rect 5997 10551 6055 10557
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 10244 10588 10272 10628
rect 10321 10625 10333 10659
rect 10367 10625 10379 10659
rect 10321 10619 10379 10625
rect 10965 10659 11023 10665
rect 10965 10625 10977 10659
rect 11011 10656 11023 10659
rect 11054 10656 11060 10668
rect 11011 10628 11060 10656
rect 11011 10625 11023 10628
rect 10965 10619 11023 10625
rect 11054 10616 11060 10628
rect 11112 10656 11118 10668
rect 11790 10656 11796 10668
rect 11112 10628 11796 10656
rect 11112 10616 11118 10628
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 13906 10656 13912 10668
rect 13867 10628 13912 10656
rect 13906 10616 13912 10628
rect 13964 10616 13970 10668
rect 16114 10656 16120 10668
rect 16075 10628 16120 10656
rect 16114 10616 16120 10628
rect 16172 10616 16178 10668
rect 14182 10588 14188 10600
rect 10244 10560 12434 10588
rect 14143 10560 14188 10588
rect 12406 10520 12434 10560
rect 14182 10548 14188 10560
rect 14240 10548 14246 10600
rect 13814 10520 13820 10532
rect 12406 10492 13820 10520
rect 13814 10480 13820 10492
rect 13872 10480 13878 10532
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 8941 10455 8999 10461
rect 8941 10452 8953 10455
rect 8352 10424 8953 10452
rect 8352 10412 8358 10424
rect 8941 10421 8953 10424
rect 8987 10452 8999 10455
rect 9398 10452 9404 10464
rect 8987 10424 9404 10452
rect 8987 10421 8999 10424
rect 8941 10415 8999 10421
rect 9398 10412 9404 10424
rect 9456 10412 9462 10464
rect 10318 10412 10324 10464
rect 10376 10452 10382 10464
rect 10873 10455 10931 10461
rect 10873 10452 10885 10455
rect 10376 10424 10885 10452
rect 10376 10412 10382 10424
rect 10873 10421 10885 10424
rect 10919 10421 10931 10455
rect 10873 10415 10931 10421
rect 11146 10412 11152 10464
rect 11204 10452 11210 10464
rect 12989 10455 13047 10461
rect 12989 10452 13001 10455
rect 11204 10424 13001 10452
rect 11204 10412 11210 10424
rect 12989 10421 13001 10424
rect 13035 10421 13047 10455
rect 12989 10415 13047 10421
rect 13538 10412 13544 10464
rect 13596 10452 13602 10464
rect 15657 10455 15715 10461
rect 15657 10452 15669 10455
rect 13596 10424 15669 10452
rect 13596 10412 13602 10424
rect 15657 10421 15669 10424
rect 15703 10421 15715 10455
rect 16206 10452 16212 10464
rect 16167 10424 16212 10452
rect 15657 10415 15715 10421
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 1104 10362 16836 10384
rect 1104 10310 2916 10362
rect 2968 10310 2980 10362
rect 3032 10310 3044 10362
rect 3096 10310 3108 10362
rect 3160 10310 3172 10362
rect 3224 10310 6849 10362
rect 6901 10310 6913 10362
rect 6965 10310 6977 10362
rect 7029 10310 7041 10362
rect 7093 10310 7105 10362
rect 7157 10310 10782 10362
rect 10834 10310 10846 10362
rect 10898 10310 10910 10362
rect 10962 10310 10974 10362
rect 11026 10310 11038 10362
rect 11090 10310 14715 10362
rect 14767 10310 14779 10362
rect 14831 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 16836 10362
rect 1104 10288 16836 10310
rect 2961 10251 3019 10257
rect 2961 10217 2973 10251
rect 3007 10248 3019 10251
rect 4614 10248 4620 10260
rect 3007 10220 4620 10248
rect 3007 10217 3019 10220
rect 2961 10211 3019 10217
rect 4614 10208 4620 10220
rect 4672 10248 4678 10260
rect 5350 10248 5356 10260
rect 4672 10220 5356 10248
rect 4672 10208 4678 10220
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 5718 10248 5724 10260
rect 5631 10220 5724 10248
rect 5718 10208 5724 10220
rect 5776 10248 5782 10260
rect 5902 10248 5908 10260
rect 5776 10220 5908 10248
rect 5776 10208 5782 10220
rect 5902 10208 5908 10220
rect 5960 10208 5966 10260
rect 10873 10251 10931 10257
rect 10873 10217 10885 10251
rect 10919 10248 10931 10251
rect 11422 10248 11428 10260
rect 10919 10220 11428 10248
rect 10919 10217 10931 10220
rect 10873 10211 10931 10217
rect 11422 10208 11428 10220
rect 11480 10208 11486 10260
rect 13541 10251 13599 10257
rect 13541 10217 13553 10251
rect 13587 10248 13599 10251
rect 14182 10248 14188 10260
rect 13587 10220 14188 10248
rect 13587 10217 13599 10220
rect 13541 10211 13599 10217
rect 14182 10208 14188 10220
rect 14240 10208 14246 10260
rect 4062 10140 4068 10192
rect 4120 10180 4126 10192
rect 15102 10180 15108 10192
rect 4120 10152 15108 10180
rect 4120 10140 4126 10152
rect 15102 10140 15108 10152
rect 15160 10140 15166 10192
rect 7558 10112 7564 10124
rect 7519 10084 7564 10112
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 7742 10112 7748 10124
rect 7703 10084 7748 10112
rect 7742 10072 7748 10084
rect 7800 10072 7806 10124
rect 9490 10112 9496 10124
rect 9324 10084 9496 10112
rect 1578 10044 1584 10056
rect 1539 10016 1584 10044
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10044 4583 10047
rect 5258 10044 5264 10056
rect 4571 10016 5264 10044
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 5258 10004 5264 10016
rect 5316 10044 5322 10056
rect 9324 10053 9352 10084
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 16025 10115 16083 10121
rect 16025 10081 16037 10115
rect 16071 10112 16083 10115
rect 16114 10112 16120 10124
rect 16071 10084 16120 10112
rect 16071 10081 16083 10084
rect 16025 10075 16083 10081
rect 16114 10072 16120 10084
rect 16172 10072 16178 10124
rect 7837 10047 7895 10053
rect 7837 10044 7849 10047
rect 5316 10016 7849 10044
rect 5316 10004 5322 10016
rect 7837 10013 7849 10016
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 9398 10004 9404 10056
rect 9456 10044 9462 10056
rect 12897 10047 12955 10053
rect 9456 10016 9501 10044
rect 9456 10004 9462 10016
rect 12897 10013 12909 10047
rect 12943 10044 12955 10047
rect 13538 10044 13544 10056
rect 12943 10016 13544 10044
rect 12943 10013 12955 10016
rect 12897 10007 12955 10013
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 13630 10004 13636 10056
rect 13688 10044 13694 10056
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 13688 10016 14289 10044
rect 13688 10004 13694 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 1848 9979 1906 9985
rect 1848 9945 1860 9979
rect 1894 9976 1906 9979
rect 1946 9976 1952 9988
rect 1894 9948 1952 9976
rect 1894 9945 1906 9948
rect 1848 9939 1906 9945
rect 1946 9936 1952 9948
rect 2004 9936 2010 9988
rect 3326 9936 3332 9988
rect 3384 9976 3390 9988
rect 4157 9979 4215 9985
rect 4157 9976 4169 9979
rect 3384 9948 4169 9976
rect 3384 9936 3390 9948
rect 4157 9945 4169 9948
rect 4203 9945 4215 9979
rect 4157 9939 4215 9945
rect 4249 9979 4307 9985
rect 4249 9945 4261 9979
rect 4295 9976 4307 9979
rect 4614 9976 4620 9988
rect 4295 9948 4620 9976
rect 4295 9945 4307 9948
rect 4249 9939 4307 9945
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 7009 9979 7067 9985
rect 7009 9945 7021 9979
rect 7055 9976 7067 9979
rect 10410 9976 10416 9988
rect 7055 9948 10416 9976
rect 7055 9945 7067 9948
rect 7009 9939 7067 9945
rect 10410 9936 10416 9948
rect 10468 9936 10474 9988
rect 12161 9979 12219 9985
rect 12161 9945 12173 9979
rect 12207 9976 12219 9979
rect 13648 9976 13676 10004
rect 12207 9948 13676 9976
rect 12207 9945 12219 9948
rect 12161 9939 12219 9945
rect 3970 9908 3976 9920
rect 3931 9880 3976 9908
rect 3970 9868 3976 9880
rect 4028 9868 4034 9920
rect 4341 9911 4399 9917
rect 4341 9877 4353 9911
rect 4387 9908 4399 9911
rect 4522 9908 4528 9920
rect 4387 9880 4528 9908
rect 4387 9877 4399 9880
rect 4341 9871 4399 9877
rect 4522 9868 4528 9880
rect 4580 9868 4586 9920
rect 8205 9911 8263 9917
rect 8205 9877 8217 9911
rect 8251 9908 8263 9911
rect 8386 9908 8392 9920
rect 8251 9880 8392 9908
rect 8251 9877 8263 9880
rect 8205 9871 8263 9877
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 9398 9908 9404 9920
rect 9359 9880 9404 9908
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 12713 9911 12771 9917
rect 12713 9877 12725 9911
rect 12759 9908 12771 9911
rect 14182 9908 14188 9920
rect 12759 9880 14188 9908
rect 12759 9877 12771 9880
rect 12713 9871 12771 9877
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 1104 9818 16995 9840
rect 1104 9766 4882 9818
rect 4934 9766 4946 9818
rect 4998 9766 5010 9818
rect 5062 9766 5074 9818
rect 5126 9766 5138 9818
rect 5190 9766 8815 9818
rect 8867 9766 8879 9818
rect 8931 9766 8943 9818
rect 8995 9766 9007 9818
rect 9059 9766 9071 9818
rect 9123 9766 12748 9818
rect 12800 9766 12812 9818
rect 12864 9766 12876 9818
rect 12928 9766 12940 9818
rect 12992 9766 13004 9818
rect 13056 9766 16681 9818
rect 16733 9766 16745 9818
rect 16797 9766 16809 9818
rect 16861 9766 16873 9818
rect 16925 9766 16937 9818
rect 16989 9766 16995 9818
rect 1104 9744 16995 9766
rect 16206 9704 16212 9716
rect 8312 9676 9720 9704
rect 8312 9648 8340 9676
rect 3326 9596 3332 9648
rect 3384 9636 3390 9648
rect 3421 9639 3479 9645
rect 3421 9636 3433 9639
rect 3384 9608 3433 9636
rect 3384 9596 3390 9608
rect 3421 9605 3433 9608
rect 3467 9605 3479 9639
rect 3421 9599 3479 9605
rect 4430 9596 4436 9648
rect 4488 9596 4494 9648
rect 6362 9596 6368 9648
rect 6420 9636 6426 9648
rect 6549 9639 6607 9645
rect 6549 9636 6561 9639
rect 6420 9608 6561 9636
rect 6420 9596 6426 9608
rect 6549 9605 6561 9608
rect 6595 9605 6607 9639
rect 8294 9636 8300 9648
rect 6549 9599 6607 9605
rect 6932 9608 8300 9636
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9537 2283 9571
rect 2225 9531 2283 9537
rect 2240 9364 2268 9531
rect 5350 9528 5356 9580
rect 5408 9568 5414 9580
rect 5629 9571 5687 9577
rect 5629 9568 5641 9571
rect 5408 9540 5641 9568
rect 5408 9528 5414 9540
rect 5629 9537 5641 9540
rect 5675 9537 5687 9571
rect 5810 9568 5816 9580
rect 5771 9540 5816 9568
rect 5629 9531 5687 9537
rect 5810 9528 5816 9540
rect 5868 9528 5874 9580
rect 6932 9577 6960 9608
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 9398 9596 9404 9648
rect 9456 9596 9462 9648
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9537 6699 9571
rect 6641 9531 6699 9537
rect 6917 9571 6975 9577
rect 6917 9537 6929 9571
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 8110 9568 8116 9580
rect 8071 9540 8116 9568
rect 7377 9531 7435 9537
rect 3145 9503 3203 9509
rect 3145 9500 3157 9503
rect 2332 9472 3157 9500
rect 2332 9441 2360 9472
rect 3145 9469 3157 9472
rect 3191 9469 3203 9503
rect 3145 9463 3203 9469
rect 4154 9460 4160 9512
rect 4212 9500 4218 9512
rect 4212 9472 4844 9500
rect 4212 9460 4218 9472
rect 2317 9435 2375 9441
rect 2317 9401 2329 9435
rect 2363 9401 2375 9435
rect 2317 9395 2375 9401
rect 4816 9376 4844 9472
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 6656 9500 6684 9531
rect 5132 9472 6684 9500
rect 5132 9460 5138 9472
rect 5902 9432 5908 9444
rect 5863 9404 5908 9432
rect 5902 9392 5908 9404
rect 5960 9392 5966 9444
rect 7392 9432 7420 9531
rect 8110 9528 8116 9540
rect 8168 9528 8174 9580
rect 9692 9568 9720 9676
rect 14844 9676 16212 9704
rect 14844 9636 14872 9676
rect 16206 9664 16212 9676
rect 16264 9664 16270 9716
rect 13018 9608 14872 9636
rect 15470 9596 15476 9648
rect 15528 9596 15534 9648
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 9692 9540 10701 9568
rect 10689 9537 10701 9540
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 10873 9571 10931 9577
rect 10873 9537 10885 9571
rect 10919 9537 10931 9571
rect 14182 9568 14188 9580
rect 14143 9540 14188 9568
rect 10873 9531 10931 9537
rect 7926 9460 7932 9512
rect 7984 9500 7990 9512
rect 8389 9503 8447 9509
rect 8389 9500 8401 9503
rect 7984 9472 8401 9500
rect 7984 9460 7990 9472
rect 8389 9469 8401 9472
rect 8435 9469 8447 9503
rect 8389 9463 8447 9469
rect 9582 9460 9588 9512
rect 9640 9500 9646 9512
rect 10888 9500 10916 9531
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 9640 9472 10916 9500
rect 11701 9503 11759 9509
rect 9640 9460 9646 9472
rect 11701 9469 11713 9503
rect 11747 9469 11759 9503
rect 13446 9500 13452 9512
rect 13407 9472 13452 9500
rect 11701 9463 11759 9469
rect 6012 9404 7420 9432
rect 10965 9435 11023 9441
rect 4522 9364 4528 9376
rect 2240 9336 4528 9364
rect 4522 9324 4528 9336
rect 4580 9324 4586 9376
rect 4798 9324 4804 9376
rect 4856 9364 4862 9376
rect 4893 9367 4951 9373
rect 4893 9364 4905 9367
rect 4856 9336 4905 9364
rect 4856 9324 4862 9336
rect 4893 9333 4905 9336
rect 4939 9333 4951 9367
rect 4893 9327 4951 9333
rect 5258 9324 5264 9376
rect 5316 9364 5322 9376
rect 6012 9364 6040 9404
rect 10965 9401 10977 9435
rect 11011 9432 11023 9435
rect 11422 9432 11428 9444
rect 11011 9404 11428 9432
rect 11011 9401 11023 9404
rect 10965 9395 11023 9401
rect 11422 9392 11428 9404
rect 11480 9392 11486 9444
rect 11716 9432 11744 9463
rect 13446 9460 13452 9472
rect 13504 9460 13510 9512
rect 13722 9500 13728 9512
rect 13683 9472 13728 9500
rect 13722 9460 13728 9472
rect 13780 9460 13786 9512
rect 14461 9503 14519 9509
rect 14461 9469 14473 9503
rect 14507 9500 14519 9503
rect 15102 9500 15108 9512
rect 14507 9472 15108 9500
rect 14507 9469 14519 9472
rect 14461 9463 14519 9469
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 12342 9432 12348 9444
rect 11716 9404 12348 9432
rect 12342 9392 12348 9404
rect 12400 9392 12406 9444
rect 5316 9336 6040 9364
rect 5316 9324 5322 9336
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 7377 9367 7435 9373
rect 7377 9364 7389 9367
rect 6696 9336 7389 9364
rect 6696 9324 6702 9336
rect 7377 9333 7389 9336
rect 7423 9333 7435 9367
rect 9858 9364 9864 9376
rect 9819 9336 9864 9364
rect 7377 9327 7435 9333
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 15562 9324 15568 9376
rect 15620 9364 15626 9376
rect 15933 9367 15991 9373
rect 15933 9364 15945 9367
rect 15620 9336 15945 9364
rect 15620 9324 15626 9336
rect 15933 9333 15945 9336
rect 15979 9333 15991 9367
rect 15933 9327 15991 9333
rect 1104 9274 16836 9296
rect 1104 9222 2916 9274
rect 2968 9222 2980 9274
rect 3032 9222 3044 9274
rect 3096 9222 3108 9274
rect 3160 9222 3172 9274
rect 3224 9222 6849 9274
rect 6901 9222 6913 9274
rect 6965 9222 6977 9274
rect 7029 9222 7041 9274
rect 7093 9222 7105 9274
rect 7157 9222 10782 9274
rect 10834 9222 10846 9274
rect 10898 9222 10910 9274
rect 10962 9222 10974 9274
rect 11026 9222 11038 9274
rect 11090 9222 14715 9274
rect 14767 9222 14779 9274
rect 14831 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 16836 9274
rect 1104 9200 16836 9222
rect 7558 9120 7564 9172
rect 7616 9160 7622 9172
rect 11790 9160 11796 9172
rect 7616 9132 11376 9160
rect 11751 9132 11796 9160
rect 7616 9120 7622 9132
rect 4246 9092 4252 9104
rect 4159 9064 4252 9092
rect 2961 8959 3019 8965
rect 2961 8925 2973 8959
rect 3007 8956 3019 8959
rect 3510 8956 3516 8968
rect 3007 8928 3516 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 3510 8916 3516 8928
rect 3568 8916 3574 8968
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8956 4123 8959
rect 4172 8956 4200 9064
rect 4246 9052 4252 9064
rect 4304 9092 4310 9104
rect 5350 9092 5356 9104
rect 4304 9064 5356 9092
rect 4304 9052 4310 9064
rect 5350 9052 5356 9064
rect 5408 9052 5414 9104
rect 11348 9036 11376 9132
rect 11790 9120 11796 9132
rect 11848 9120 11854 9172
rect 13173 9163 13231 9169
rect 13173 9129 13185 9163
rect 13219 9160 13231 9163
rect 13446 9160 13452 9172
rect 13219 9132 13452 9160
rect 13219 9129 13231 9132
rect 13173 9123 13231 9129
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 15102 9160 15108 9172
rect 15063 9132 15108 9160
rect 15102 9120 15108 9132
rect 15160 9120 15166 9172
rect 12437 9095 12495 9101
rect 12437 9061 12449 9095
rect 12483 9092 12495 9095
rect 13722 9092 13728 9104
rect 12483 9064 13728 9092
rect 12483 9061 12495 9064
rect 12437 9055 12495 9061
rect 13722 9052 13728 9064
rect 13780 9052 13786 9104
rect 4430 9024 4436 9036
rect 4391 8996 4436 9024
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 6270 8984 6276 9036
rect 6328 9024 6334 9036
rect 6365 9027 6423 9033
rect 6365 9024 6377 9027
rect 6328 8996 6377 9024
rect 6328 8984 6334 8996
rect 6365 8993 6377 8996
rect 6411 8993 6423 9027
rect 6638 9024 6644 9036
rect 6599 8996 6644 9024
rect 6365 8987 6423 8993
rect 6638 8984 6644 8996
rect 6696 8984 6702 9036
rect 9858 9024 9864 9036
rect 8496 8996 9864 9024
rect 4338 8956 4344 8968
rect 4111 8928 4200 8956
rect 4299 8928 4344 8956
rect 4111 8925 4123 8928
rect 4065 8919 4123 8925
rect 4338 8916 4344 8928
rect 4396 8956 4402 8968
rect 5074 8956 5080 8968
rect 4396 8928 5080 8956
rect 4396 8916 4402 8928
rect 5074 8916 5080 8928
rect 5132 8916 5138 8968
rect 7466 8916 7472 8968
rect 7524 8956 7530 8968
rect 8496 8956 8524 8996
rect 7524 8928 8524 8956
rect 8573 8959 8631 8965
rect 7524 8916 7530 8928
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 9214 8956 9220 8968
rect 8619 8928 9220 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 9508 8965 9536 8996
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 10318 9024 10324 9036
rect 10279 8996 10324 9024
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 11330 8984 11336 9036
rect 11388 9024 11394 9036
rect 11388 8996 12296 9024
rect 11388 8984 11394 8996
rect 9493 8959 9551 8965
rect 9493 8925 9505 8959
rect 9539 8925 9551 8959
rect 9493 8919 9551 8925
rect 9585 8959 9643 8965
rect 9585 8925 9597 8959
rect 9631 8956 9643 8959
rect 10045 8959 10103 8965
rect 10045 8956 10057 8959
rect 9631 8928 10057 8956
rect 9631 8925 9643 8928
rect 9585 8919 9643 8925
rect 10045 8925 10057 8928
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 11422 8916 11428 8968
rect 11480 8916 11486 8968
rect 12268 8965 12296 8996
rect 12253 8959 12311 8965
rect 12253 8925 12265 8959
rect 12299 8925 12311 8959
rect 12253 8919 12311 8925
rect 2716 8891 2774 8897
rect 2716 8857 2728 8891
rect 2762 8888 2774 8891
rect 3694 8888 3700 8900
rect 2762 8860 3700 8888
rect 2762 8857 2774 8860
rect 2716 8851 2774 8857
rect 3694 8848 3700 8860
rect 3752 8848 3758 8900
rect 5902 8848 5908 8900
rect 5960 8848 5966 8900
rect 8328 8891 8386 8897
rect 8328 8857 8340 8891
rect 8374 8888 8386 8891
rect 10226 8888 10232 8900
rect 8374 8860 10232 8888
rect 8374 8857 8386 8860
rect 8328 8851 8386 8857
rect 10226 8848 10232 8860
rect 10284 8848 10290 8900
rect 12268 8888 12296 8919
rect 12342 8916 12348 8968
rect 12400 8956 12406 8968
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 12400 8928 13001 8956
rect 12400 8916 12406 8928
rect 12989 8925 13001 8928
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8956 14611 8959
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 14599 8928 15301 8956
rect 14599 8925 14611 8928
rect 14553 8919 14611 8925
rect 15289 8925 15301 8928
rect 15335 8956 15347 8959
rect 15562 8956 15568 8968
rect 15335 8928 15568 8956
rect 15335 8925 15347 8928
rect 15289 8919 15347 8925
rect 15562 8916 15568 8928
rect 15620 8916 15626 8968
rect 15933 8959 15991 8965
rect 15933 8925 15945 8959
rect 15979 8956 15991 8959
rect 16114 8956 16120 8968
rect 15979 8928 16120 8956
rect 15979 8925 15991 8928
rect 15933 8919 15991 8925
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 13262 8888 13268 8900
rect 12268 8860 13268 8888
rect 13262 8848 13268 8860
rect 13320 8848 13326 8900
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 2590 8820 2596 8832
rect 1627 8792 2596 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 2590 8780 2596 8792
rect 2648 8780 2654 8832
rect 4522 8780 4528 8832
rect 4580 8820 4586 8832
rect 4893 8823 4951 8829
rect 4893 8820 4905 8823
rect 4580 8792 4905 8820
rect 4580 8780 4586 8792
rect 4893 8789 4905 8792
rect 4939 8820 4951 8823
rect 5442 8820 5448 8832
rect 4939 8792 5448 8820
rect 4939 8789 4951 8792
rect 4893 8783 4951 8789
rect 5442 8780 5448 8792
rect 5500 8780 5506 8832
rect 6086 8780 6092 8832
rect 6144 8820 6150 8832
rect 7193 8823 7251 8829
rect 7193 8820 7205 8823
rect 6144 8792 7205 8820
rect 6144 8780 6150 8792
rect 7193 8789 7205 8792
rect 7239 8789 7251 8823
rect 7193 8783 7251 8789
rect 14369 8823 14427 8829
rect 14369 8789 14381 8823
rect 14415 8820 14427 8823
rect 14642 8820 14648 8832
rect 14415 8792 14648 8820
rect 14415 8789 14427 8792
rect 14369 8783 14427 8789
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 15838 8820 15844 8832
rect 15799 8792 15844 8820
rect 15838 8780 15844 8792
rect 15896 8780 15902 8832
rect 1104 8730 16995 8752
rect 1104 8678 4882 8730
rect 4934 8678 4946 8730
rect 4998 8678 5010 8730
rect 5062 8678 5074 8730
rect 5126 8678 5138 8730
rect 5190 8678 8815 8730
rect 8867 8678 8879 8730
rect 8931 8678 8943 8730
rect 8995 8678 9007 8730
rect 9059 8678 9071 8730
rect 9123 8678 12748 8730
rect 12800 8678 12812 8730
rect 12864 8678 12876 8730
rect 12928 8678 12940 8730
rect 12992 8678 13004 8730
rect 13056 8678 16681 8730
rect 16733 8678 16745 8730
rect 16797 8678 16809 8730
rect 16861 8678 16873 8730
rect 16925 8678 16937 8730
rect 16989 8678 16995 8730
rect 1104 8656 16995 8678
rect 1762 8616 1768 8628
rect 1723 8588 1768 8616
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 5077 8619 5135 8625
rect 2792 8588 4384 8616
rect 1486 8440 1492 8492
rect 1544 8480 1550 8492
rect 1581 8483 1639 8489
rect 1581 8480 1593 8483
rect 1544 8452 1593 8480
rect 1544 8440 1550 8452
rect 1581 8449 1593 8452
rect 1627 8449 1639 8483
rect 1581 8443 1639 8449
rect 2590 8440 2596 8492
rect 2648 8480 2654 8492
rect 2792 8489 2820 8588
rect 4356 8548 4384 8588
rect 5077 8585 5089 8619
rect 5123 8616 5135 8619
rect 7926 8616 7932 8628
rect 5123 8588 7932 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 15470 8616 15476 8628
rect 15431 8588 15476 8616
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 6917 8551 6975 8557
rect 4356 8520 5396 8548
rect 5368 8492 5396 8520
rect 6917 8517 6929 8551
rect 6963 8548 6975 8551
rect 7558 8548 7564 8560
rect 6963 8520 7564 8548
rect 6963 8517 6975 8520
rect 6917 8511 6975 8517
rect 7558 8508 7564 8520
rect 7616 8508 7622 8560
rect 9490 8508 9496 8560
rect 9548 8548 9554 8560
rect 15838 8548 15844 8560
rect 9548 8520 11928 8548
rect 13938 8520 15844 8548
rect 9548 8508 9554 8520
rect 2777 8483 2835 8489
rect 2777 8480 2789 8483
rect 2648 8452 2789 8480
rect 2648 8440 2654 8452
rect 2777 8449 2789 8452
rect 2823 8449 2835 8483
rect 2777 8443 2835 8449
rect 4154 8440 4160 8492
rect 4212 8440 4218 8492
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8449 5227 8483
rect 5169 8443 5227 8449
rect 3053 8415 3111 8421
rect 3053 8381 3065 8415
rect 3099 8412 3111 8415
rect 4614 8412 4620 8424
rect 3099 8384 4620 8412
rect 3099 8381 3111 8384
rect 3053 8375 3111 8381
rect 4614 8372 4620 8384
rect 4672 8372 4678 8424
rect 5184 8412 5212 8443
rect 5350 8440 5356 8492
rect 5408 8480 5414 8492
rect 5629 8483 5687 8489
rect 5629 8480 5641 8483
rect 5408 8452 5641 8480
rect 5408 8440 5414 8452
rect 5629 8449 5641 8452
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 5810 8440 5816 8492
rect 5868 8480 5874 8492
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5868 8452 5917 8480
rect 5868 8440 5874 8452
rect 5905 8449 5917 8452
rect 5951 8480 5963 8483
rect 9508 8480 9536 8508
rect 9766 8480 9772 8492
rect 5951 8452 9536 8480
rect 9727 8452 9772 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 11057 8483 11115 8489
rect 11057 8449 11069 8483
rect 11103 8480 11115 8483
rect 11238 8480 11244 8492
rect 11103 8452 11244 8480
rect 11103 8449 11115 8452
rect 11057 8443 11115 8449
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11698 8480 11704 8492
rect 11659 8452 11704 8480
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 11900 8489 11928 8520
rect 15838 8508 15844 8520
rect 15896 8508 15902 8560
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8449 11943 8483
rect 11885 8443 11943 8449
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 15565 8483 15623 8489
rect 14700 8452 14745 8480
rect 14700 8440 14706 8452
rect 15565 8449 15577 8483
rect 15611 8480 15623 8483
rect 16114 8480 16120 8492
rect 15611 8452 16120 8480
rect 15611 8449 15623 8452
rect 15565 8443 15623 8449
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 7282 8412 7288 8424
rect 5184 8384 6132 8412
rect 7243 8384 7288 8412
rect 4430 8304 4436 8356
rect 4488 8344 4494 8356
rect 4525 8347 4583 8353
rect 4525 8344 4537 8347
rect 4488 8316 4537 8344
rect 4488 8304 4494 8316
rect 4525 8313 4537 8316
rect 4571 8344 4583 8347
rect 5258 8344 5264 8356
rect 4571 8316 5264 8344
rect 4571 8313 4583 8316
rect 4525 8307 4583 8313
rect 5258 8304 5264 8316
rect 5316 8304 5322 8356
rect 5810 8304 5816 8356
rect 5868 8344 5874 8356
rect 5905 8347 5963 8353
rect 5905 8344 5917 8347
rect 5868 8316 5917 8344
rect 5868 8304 5874 8316
rect 5905 8313 5917 8316
rect 5951 8313 5963 8347
rect 6104 8344 6132 8384
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 14366 8412 14372 8424
rect 14327 8384 14372 8412
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 7466 8344 7472 8356
rect 6104 8316 7472 8344
rect 5905 8307 5963 8313
rect 7466 8304 7472 8316
rect 7524 8304 7530 8356
rect 8128 8316 8432 8344
rect 5994 8236 6000 8288
rect 6052 8276 6058 8288
rect 6733 8279 6791 8285
rect 6733 8276 6745 8279
rect 6052 8248 6745 8276
rect 6052 8236 6058 8248
rect 6733 8245 6745 8248
rect 6779 8245 6791 8279
rect 6733 8239 6791 8245
rect 6917 8279 6975 8285
rect 6917 8245 6929 8279
rect 6963 8276 6975 8279
rect 8128 8276 8156 8316
rect 8294 8276 8300 8288
rect 6963 8248 8156 8276
rect 8255 8248 8300 8276
rect 6963 8245 6975 8248
rect 6917 8239 6975 8245
rect 8294 8236 8300 8248
rect 8352 8236 8358 8288
rect 8404 8276 8432 8316
rect 11330 8304 11336 8356
rect 11388 8344 11394 8356
rect 11977 8347 12035 8353
rect 11977 8344 11989 8347
rect 11388 8316 11989 8344
rect 11388 8304 11394 8316
rect 11977 8313 11989 8316
rect 12023 8313 12035 8347
rect 11977 8307 12035 8313
rect 8478 8276 8484 8288
rect 8404 8248 8484 8276
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 11057 8279 11115 8285
rect 11057 8245 11069 8279
rect 11103 8276 11115 8279
rect 12066 8276 12072 8288
rect 11103 8248 12072 8276
rect 11103 8245 11115 8248
rect 11057 8239 11115 8245
rect 12066 8236 12072 8248
rect 12124 8236 12130 8288
rect 12894 8276 12900 8288
rect 12855 8248 12900 8276
rect 12894 8236 12900 8248
rect 12952 8236 12958 8288
rect 1104 8186 16836 8208
rect 1104 8134 2916 8186
rect 2968 8134 2980 8186
rect 3032 8134 3044 8186
rect 3096 8134 3108 8186
rect 3160 8134 3172 8186
rect 3224 8134 6849 8186
rect 6901 8134 6913 8186
rect 6965 8134 6977 8186
rect 7029 8134 7041 8186
rect 7093 8134 7105 8186
rect 7157 8134 10782 8186
rect 10834 8134 10846 8186
rect 10898 8134 10910 8186
rect 10962 8134 10974 8186
rect 11026 8134 11038 8186
rect 11090 8134 14715 8186
rect 14767 8134 14779 8186
rect 14831 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 16836 8186
rect 1104 8112 16836 8134
rect 1762 8072 1768 8084
rect 1723 8044 1768 8072
rect 1762 8032 1768 8044
rect 1820 8032 1826 8084
rect 9309 8075 9367 8081
rect 9309 8041 9321 8075
rect 9355 8072 9367 8075
rect 9766 8072 9772 8084
rect 9355 8044 9772 8072
rect 9355 8041 9367 8044
rect 9309 8035 9367 8041
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 12342 8072 12348 8084
rect 9876 8044 12348 8072
rect 2685 8007 2743 8013
rect 2685 7973 2697 8007
rect 2731 8004 2743 8007
rect 3786 8004 3792 8016
rect 2731 7976 3792 8004
rect 2731 7973 2743 7976
rect 2685 7967 2743 7973
rect 3786 7964 3792 7976
rect 3844 7964 3850 8016
rect 4065 8007 4123 8013
rect 4065 7973 4077 8007
rect 4111 8004 4123 8007
rect 4154 8004 4160 8016
rect 4111 7976 4160 8004
rect 4111 7973 4123 7976
rect 4065 7967 4123 7973
rect 4154 7964 4160 7976
rect 4212 7964 4218 8016
rect 5718 7964 5724 8016
rect 5776 8004 5782 8016
rect 9122 8004 9128 8016
rect 5776 7976 9128 8004
rect 5776 7964 5782 7976
rect 9122 7964 9128 7976
rect 9180 7964 9186 8016
rect 8294 7936 8300 7948
rect 7024 7908 8300 7936
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 1670 7868 1676 7880
rect 1627 7840 1676 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 1670 7828 1676 7840
rect 1728 7828 1734 7880
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7868 2743 7871
rect 3142 7868 3148 7880
rect 2731 7840 3148 7868
rect 2731 7837 2743 7840
rect 2685 7831 2743 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7868 3479 7871
rect 3878 7868 3884 7880
rect 3467 7840 3884 7868
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 3878 7828 3884 7840
rect 3936 7828 3942 7880
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 4172 7800 4200 7831
rect 4246 7828 4252 7880
rect 4304 7868 4310 7880
rect 4304 7840 4349 7868
rect 4304 7828 4310 7840
rect 5442 7828 5448 7880
rect 5500 7868 5506 7880
rect 7024 7877 7052 7908
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 9876 7936 9904 8044
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 13265 8075 13323 8081
rect 13265 8041 13277 8075
rect 13311 8072 13323 8075
rect 14366 8072 14372 8084
rect 13311 8044 14372 8072
rect 13311 8041 13323 8044
rect 13265 8035 13323 8041
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 12066 7936 12072 7948
rect 8588 7908 9904 7936
rect 12027 7908 12072 7936
rect 7009 7871 7067 7877
rect 5500 7840 5764 7868
rect 5500 7828 5506 7840
rect 4338 7800 4344 7812
rect 4172 7772 4344 7800
rect 4338 7760 4344 7772
rect 4396 7800 4402 7812
rect 5736 7800 5764 7840
rect 7009 7837 7021 7871
rect 7055 7837 7067 7871
rect 8202 7868 8208 7880
rect 8163 7840 8208 7868
rect 7009 7831 7067 7837
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 8386 7868 8392 7880
rect 8347 7840 8392 7868
rect 8386 7828 8392 7840
rect 8444 7828 8450 7880
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 8588 7877 8616 7908
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 8573 7871 8631 7877
rect 8573 7868 8585 7871
rect 8536 7840 8585 7868
rect 8536 7828 8542 7840
rect 8573 7837 8585 7840
rect 8619 7837 8631 7871
rect 8573 7831 8631 7837
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 9180 7840 9225 7868
rect 9180 7828 9186 7840
rect 12894 7828 12900 7880
rect 12952 7868 12958 7880
rect 13078 7868 13084 7880
rect 12952 7840 13084 7868
rect 12952 7828 12958 7840
rect 13078 7828 13084 7840
rect 13136 7828 13142 7880
rect 7742 7800 7748 7812
rect 4396 7772 5580 7800
rect 5736 7772 7748 7800
rect 4396 7760 4402 7772
rect 5552 7744 5580 7772
rect 7742 7760 7748 7772
rect 7800 7760 7806 7812
rect 8297 7803 8355 7809
rect 8297 7769 8309 7803
rect 8343 7800 8355 7803
rect 10042 7800 10048 7812
rect 8343 7772 10048 7800
rect 8343 7769 8355 7772
rect 8297 7763 8355 7769
rect 10042 7760 10048 7772
rect 10100 7800 10106 7812
rect 10100 7772 10364 7800
rect 10100 7760 10106 7772
rect 3237 7735 3295 7741
rect 3237 7701 3249 7735
rect 3283 7732 3295 7735
rect 3970 7732 3976 7744
rect 3283 7704 3976 7732
rect 3283 7701 3295 7704
rect 3237 7695 3295 7701
rect 3970 7692 3976 7704
rect 4028 7692 4034 7744
rect 5534 7732 5540 7744
rect 5495 7704 5540 7732
rect 5534 7692 5540 7704
rect 5592 7692 5598 7744
rect 8018 7732 8024 7744
rect 7979 7704 8024 7732
rect 8018 7692 8024 7704
rect 8076 7692 8082 7744
rect 10336 7741 10364 7772
rect 11330 7760 11336 7812
rect 11388 7760 11394 7812
rect 11793 7803 11851 7809
rect 11793 7769 11805 7803
rect 11839 7800 11851 7803
rect 11882 7800 11888 7812
rect 11839 7772 11888 7800
rect 11839 7769 11851 7772
rect 11793 7763 11851 7769
rect 11882 7760 11888 7772
rect 11940 7760 11946 7812
rect 10321 7735 10379 7741
rect 10321 7701 10333 7735
rect 10367 7701 10379 7735
rect 10321 7695 10379 7701
rect 1104 7642 16995 7664
rect 1104 7590 4882 7642
rect 4934 7590 4946 7642
rect 4998 7590 5010 7642
rect 5062 7590 5074 7642
rect 5126 7590 5138 7642
rect 5190 7590 8815 7642
rect 8867 7590 8879 7642
rect 8931 7590 8943 7642
rect 8995 7590 9007 7642
rect 9059 7590 9071 7642
rect 9123 7590 12748 7642
rect 12800 7590 12812 7642
rect 12864 7590 12876 7642
rect 12928 7590 12940 7642
rect 12992 7590 13004 7642
rect 13056 7590 16681 7642
rect 16733 7590 16745 7642
rect 16797 7590 16809 7642
rect 16861 7590 16873 7642
rect 16925 7590 16937 7642
rect 16989 7590 16995 7642
rect 1104 7568 16995 7590
rect 1486 7488 1492 7540
rect 1544 7528 1550 7540
rect 1581 7531 1639 7537
rect 1581 7528 1593 7531
rect 1544 7500 1593 7528
rect 1544 7488 1550 7500
rect 1581 7497 1593 7500
rect 1627 7497 1639 7531
rect 2774 7528 2780 7540
rect 1581 7491 1639 7497
rect 2516 7500 2780 7528
rect 2516 7469 2544 7500
rect 2774 7488 2780 7500
rect 2832 7488 2838 7540
rect 3907 7531 3965 7537
rect 3907 7497 3919 7531
rect 3953 7528 3965 7531
rect 5442 7528 5448 7540
rect 3953 7500 5448 7528
rect 3953 7497 3965 7500
rect 3907 7491 3965 7497
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 8297 7531 8355 7537
rect 5644 7500 8248 7528
rect 2501 7463 2559 7469
rect 2501 7429 2513 7463
rect 2547 7429 2559 7463
rect 2501 7423 2559 7429
rect 3142 7420 3148 7472
rect 3200 7460 3206 7472
rect 3697 7463 3755 7469
rect 3697 7460 3709 7463
rect 3200 7432 3709 7460
rect 3200 7420 3206 7432
rect 3697 7429 3709 7432
rect 3743 7460 3755 7463
rect 4706 7460 4712 7472
rect 3743 7432 4712 7460
rect 3743 7429 3755 7432
rect 3697 7423 3755 7429
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 5644 7460 5672 7500
rect 5460 7432 5672 7460
rect 8220 7460 8248 7500
rect 8297 7497 8309 7531
rect 8343 7528 8355 7531
rect 9490 7528 9496 7540
rect 8343 7500 9496 7528
rect 8343 7497 8355 7500
rect 8297 7491 8355 7497
rect 9490 7488 9496 7500
rect 9548 7488 9554 7540
rect 9766 7488 9772 7540
rect 9824 7528 9830 7540
rect 10413 7531 10471 7537
rect 10413 7528 10425 7531
rect 9824 7500 10425 7528
rect 9824 7488 9830 7500
rect 10413 7497 10425 7500
rect 10459 7497 10471 7531
rect 11882 7528 11888 7540
rect 11843 7500 11888 7528
rect 10413 7491 10471 7497
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 8570 7460 8576 7472
rect 8220 7432 8576 7460
rect 1762 7392 1768 7404
rect 1723 7364 1768 7392
rect 1762 7352 1768 7364
rect 1820 7352 1826 7404
rect 2590 7352 2596 7404
rect 2648 7392 2654 7404
rect 2685 7395 2743 7401
rect 2685 7392 2697 7395
rect 2648 7364 2697 7392
rect 2648 7352 2654 7364
rect 2685 7361 2697 7364
rect 2731 7361 2743 7395
rect 2685 7355 2743 7361
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7361 2835 7395
rect 4522 7392 4528 7404
rect 4483 7364 4528 7392
rect 2777 7355 2835 7361
rect 2038 7324 2044 7336
rect 1951 7296 2044 7324
rect 2038 7284 2044 7296
rect 2096 7324 2102 7336
rect 2792 7324 2820 7355
rect 4522 7352 4528 7364
rect 4580 7352 4586 7404
rect 5166 7392 5172 7404
rect 5127 7364 5172 7392
rect 5166 7352 5172 7364
rect 5224 7352 5230 7404
rect 5460 7401 5488 7432
rect 8570 7420 8576 7432
rect 8628 7420 8634 7472
rect 9585 7463 9643 7469
rect 9585 7429 9597 7463
rect 9631 7460 9643 7463
rect 9674 7460 9680 7472
rect 9631 7432 9680 7460
rect 9631 7429 9643 7432
rect 9585 7423 9643 7429
rect 9674 7420 9680 7432
rect 9732 7420 9738 7472
rect 10042 7460 10048 7472
rect 10003 7432 10048 7460
rect 10042 7420 10048 7432
rect 10100 7460 10106 7472
rect 10100 7432 11744 7460
rect 10100 7420 10106 7432
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 5994 7392 6000 7404
rect 5859 7364 6000 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 6546 7392 6552 7404
rect 6459 7364 6552 7392
rect 6546 7352 6552 7364
rect 6604 7392 6610 7404
rect 8478 7392 8484 7404
rect 6604 7364 8484 7392
rect 6604 7352 6610 7364
rect 8478 7352 8484 7364
rect 8536 7352 8542 7404
rect 9858 7352 9864 7404
rect 9916 7392 9922 7404
rect 10229 7395 10287 7401
rect 10229 7392 10241 7395
rect 9916 7364 10241 7392
rect 9916 7352 9922 7364
rect 10229 7361 10241 7364
rect 10275 7361 10287 7395
rect 10229 7355 10287 7361
rect 10318 7352 10324 7404
rect 10376 7392 10382 7404
rect 11716 7401 11744 7432
rect 12342 7420 12348 7472
rect 12400 7460 12406 7472
rect 12400 7432 13124 7460
rect 12400 7420 12406 7432
rect 13096 7401 13124 7432
rect 11701 7395 11759 7401
rect 10376 7364 10421 7392
rect 10376 7352 10382 7364
rect 11701 7361 11713 7395
rect 11747 7361 11759 7395
rect 12621 7395 12679 7401
rect 12621 7392 12633 7395
rect 11701 7355 11759 7361
rect 12406 7364 12633 7392
rect 3602 7324 3608 7336
rect 2096 7296 2544 7324
rect 2792 7296 3608 7324
rect 2096 7284 2102 7296
rect 2516 7265 2544 7296
rect 3602 7284 3608 7296
rect 3660 7324 3666 7336
rect 6825 7327 6883 7333
rect 3660 7296 5948 7324
rect 3660 7284 3666 7296
rect 2501 7259 2559 7265
rect 2501 7225 2513 7259
rect 2547 7225 2559 7259
rect 5626 7256 5632 7268
rect 2501 7219 2559 7225
rect 3896 7228 5632 7256
rect 3896 7200 3924 7228
rect 5626 7216 5632 7228
rect 5684 7216 5690 7268
rect 5920 7265 5948 7296
rect 6825 7293 6837 7327
rect 6871 7324 6883 7327
rect 7558 7324 7564 7336
rect 6871 7296 7564 7324
rect 6871 7293 6883 7296
rect 6825 7287 6883 7293
rect 7558 7284 7564 7296
rect 7616 7284 7622 7336
rect 10597 7327 10655 7333
rect 10597 7293 10609 7327
rect 10643 7324 10655 7327
rect 12406 7324 12434 7364
rect 12621 7361 12633 7364
rect 12667 7361 12679 7395
rect 12621 7355 12679 7361
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7361 13139 7395
rect 13262 7392 13268 7404
rect 13223 7364 13268 7392
rect 13081 7355 13139 7361
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 10643 7296 12434 7324
rect 10643 7293 10655 7296
rect 10597 7287 10655 7293
rect 5905 7259 5963 7265
rect 5905 7225 5917 7259
rect 5951 7225 5963 7259
rect 6730 7256 6736 7268
rect 6691 7228 6736 7256
rect 5905 7219 5963 7225
rect 6730 7216 6736 7228
rect 6788 7216 6794 7268
rect 8202 7216 8208 7268
rect 8260 7256 8266 7268
rect 13081 7259 13139 7265
rect 13081 7256 13093 7259
rect 8260 7228 13093 7256
rect 8260 7216 8266 7228
rect 13081 7225 13093 7228
rect 13127 7225 13139 7259
rect 13081 7219 13139 7225
rect 1949 7191 2007 7197
rect 1949 7157 1961 7191
rect 1995 7188 2007 7191
rect 2314 7188 2320 7200
rect 1995 7160 2320 7188
rect 1995 7157 2007 7160
rect 1949 7151 2007 7157
rect 2314 7148 2320 7160
rect 2372 7148 2378 7200
rect 3878 7188 3884 7200
rect 3839 7160 3884 7188
rect 3878 7148 3884 7160
rect 3936 7148 3942 7200
rect 4065 7191 4123 7197
rect 4065 7157 4077 7191
rect 4111 7188 4123 7191
rect 4154 7188 4160 7200
rect 4111 7160 4160 7188
rect 4111 7157 4123 7160
rect 4065 7151 4123 7157
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 5350 7148 5356 7200
rect 5408 7188 5414 7200
rect 6641 7191 6699 7197
rect 6641 7188 6653 7191
rect 5408 7160 6653 7188
rect 5408 7148 5414 7160
rect 6641 7157 6653 7160
rect 6687 7157 6699 7191
rect 6641 7151 6699 7157
rect 10226 7148 10232 7200
rect 10284 7188 10290 7200
rect 12437 7191 12495 7197
rect 12437 7188 12449 7191
rect 10284 7160 12449 7188
rect 10284 7148 10290 7160
rect 12437 7157 12449 7160
rect 12483 7157 12495 7191
rect 12437 7151 12495 7157
rect 1104 7098 16836 7120
rect 1104 7046 2916 7098
rect 2968 7046 2980 7098
rect 3032 7046 3044 7098
rect 3096 7046 3108 7098
rect 3160 7046 3172 7098
rect 3224 7046 6849 7098
rect 6901 7046 6913 7098
rect 6965 7046 6977 7098
rect 7029 7046 7041 7098
rect 7093 7046 7105 7098
rect 7157 7046 10782 7098
rect 10834 7046 10846 7098
rect 10898 7046 10910 7098
rect 10962 7046 10974 7098
rect 11026 7046 11038 7098
rect 11090 7046 14715 7098
rect 14767 7046 14779 7098
rect 14831 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 16836 7098
rect 1104 7024 16836 7046
rect 1581 6987 1639 6993
rect 1581 6953 1593 6987
rect 1627 6984 1639 6987
rect 1670 6984 1676 6996
rect 1627 6956 1676 6984
rect 1627 6953 1639 6956
rect 1581 6947 1639 6953
rect 1670 6944 1676 6956
rect 1728 6944 1734 6996
rect 1949 6987 2007 6993
rect 1949 6953 1961 6987
rect 1995 6984 2007 6987
rect 2038 6984 2044 6996
rect 1995 6956 2044 6984
rect 1995 6953 2007 6956
rect 1949 6947 2007 6953
rect 2038 6944 2044 6956
rect 2096 6944 2102 6996
rect 4249 6987 4307 6993
rect 4249 6953 4261 6987
rect 4295 6984 4307 6987
rect 4522 6984 4528 6996
rect 4295 6956 4528 6984
rect 4295 6953 4307 6956
rect 4249 6947 4307 6953
rect 4522 6944 4528 6956
rect 4580 6944 4586 6996
rect 5166 6944 5172 6996
rect 5224 6984 5230 6996
rect 6546 6984 6552 6996
rect 5224 6956 6552 6984
rect 5224 6944 5230 6956
rect 6546 6944 6552 6956
rect 6604 6944 6610 6996
rect 10318 6944 10324 6996
rect 10376 6984 10382 6996
rect 11621 6987 11679 6993
rect 11621 6984 11633 6987
rect 10376 6956 11633 6984
rect 10376 6944 10382 6956
rect 11621 6953 11633 6956
rect 11667 6953 11679 6987
rect 11621 6947 11679 6953
rect 3970 6876 3976 6928
rect 4028 6916 4034 6928
rect 4028 6888 4936 6916
rect 4028 6876 4034 6888
rect 1780 6820 3280 6848
rect 1780 6792 1808 6820
rect 1762 6780 1768 6792
rect 1723 6752 1768 6780
rect 1762 6740 1768 6752
rect 1820 6740 1826 6792
rect 2038 6780 2044 6792
rect 1999 6752 2044 6780
rect 2038 6740 2044 6752
rect 2096 6740 2102 6792
rect 2590 6740 2596 6792
rect 2648 6780 2654 6792
rect 3252 6789 3280 6820
rect 3786 6808 3792 6860
rect 3844 6848 3850 6860
rect 4801 6851 4859 6857
rect 4801 6848 4813 6851
rect 3844 6820 4813 6848
rect 3844 6808 3850 6820
rect 4801 6817 4813 6820
rect 4847 6817 4859 6851
rect 4908 6848 4936 6888
rect 5077 6851 5135 6857
rect 5077 6848 5089 6851
rect 4908 6820 5089 6848
rect 4801 6811 4859 6817
rect 5077 6817 5089 6820
rect 5123 6817 5135 6851
rect 5077 6811 5135 6817
rect 5626 6808 5632 6860
rect 5684 6848 5690 6860
rect 6549 6851 6607 6857
rect 6549 6848 6561 6851
rect 5684 6820 6561 6848
rect 5684 6808 5690 6820
rect 6549 6817 6561 6820
rect 6595 6817 6607 6851
rect 8478 6848 8484 6860
rect 8234 6820 8484 6848
rect 6549 6811 6607 6817
rect 2869 6783 2927 6789
rect 2869 6780 2881 6783
rect 2648 6752 2881 6780
rect 2648 6740 2654 6752
rect 2869 6749 2881 6752
rect 2915 6749 2927 6783
rect 2869 6743 2927 6749
rect 2961 6783 3019 6789
rect 2961 6749 2973 6783
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 3053 6783 3111 6789
rect 3053 6749 3065 6783
rect 3099 6749 3111 6783
rect 3053 6743 3111 6749
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6749 3295 6783
rect 3237 6743 3295 6749
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6780 4399 6783
rect 4387 6752 4844 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 2682 6672 2688 6724
rect 2740 6712 2746 6724
rect 2976 6712 3004 6743
rect 2740 6684 3004 6712
rect 3068 6712 3096 6743
rect 3418 6712 3424 6724
rect 3068 6684 3424 6712
rect 2740 6672 2746 6684
rect 3418 6672 3424 6684
rect 3476 6672 3482 6724
rect 4172 6712 4200 6743
rect 4430 6712 4436 6724
rect 4172 6684 4436 6712
rect 4430 6672 4436 6684
rect 4488 6672 4494 6724
rect 4816 6712 4844 6752
rect 5166 6712 5172 6724
rect 4816 6684 5172 6712
rect 5166 6672 5172 6684
rect 5224 6672 5230 6724
rect 5810 6672 5816 6724
rect 5868 6672 5874 6724
rect 6564 6712 6592 6811
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 9214 6848 9220 6860
rect 9175 6820 9220 6848
rect 9214 6808 9220 6820
rect 9272 6808 9278 6860
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 7466 6780 7472 6792
rect 6696 6752 7328 6780
rect 7427 6752 7472 6780
rect 6696 6740 6702 6752
rect 7193 6715 7251 6721
rect 7193 6712 7205 6715
rect 6564 6684 7205 6712
rect 7193 6681 7205 6684
rect 7239 6681 7251 6715
rect 7300 6712 7328 6752
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 7558 6740 7564 6792
rect 7616 6780 7622 6792
rect 9306 6780 9312 6792
rect 7616 6752 7661 6780
rect 9267 6752 9312 6780
rect 7616 6740 7622 6752
rect 9306 6740 9312 6752
rect 9364 6740 9370 6792
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6780 11943 6783
rect 12805 6783 12863 6789
rect 12805 6780 12817 6783
rect 11931 6752 12817 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 12805 6749 12817 6752
rect 12851 6749 12863 6783
rect 12805 6743 12863 6749
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6780 12955 6783
rect 13078 6780 13084 6792
rect 12943 6752 13084 6780
rect 12943 6749 12955 6752
rect 12897 6743 12955 6749
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 7929 6715 7987 6721
rect 7929 6712 7941 6715
rect 7300 6684 7941 6712
rect 7193 6675 7251 6681
rect 7929 6681 7941 6684
rect 7975 6681 7987 6715
rect 7929 6675 7987 6681
rect 8297 6715 8355 6721
rect 8297 6681 8309 6715
rect 8343 6712 8355 6715
rect 8343 6684 10272 6712
rect 8343 6681 8355 6684
rect 8297 6675 8355 6681
rect 1854 6604 1860 6656
rect 1912 6644 1918 6656
rect 2593 6647 2651 6653
rect 2593 6644 2605 6647
rect 1912 6616 2605 6644
rect 1912 6604 1918 6616
rect 2593 6613 2605 6616
rect 2639 6613 2651 6647
rect 2593 6607 2651 6613
rect 4338 6604 4344 6656
rect 4396 6644 4402 6656
rect 8481 6647 8539 6653
rect 8481 6644 8493 6647
rect 4396 6616 8493 6644
rect 4396 6604 4402 6616
rect 8481 6613 8493 6616
rect 8527 6613 8539 6647
rect 10134 6644 10140 6656
rect 10095 6616 10140 6644
rect 8481 6607 8539 6613
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 10244 6644 10272 6684
rect 11146 6672 11152 6724
rect 11204 6672 11210 6724
rect 11238 6644 11244 6656
rect 10244 6616 11244 6644
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 1104 6554 16995 6576
rect 1104 6502 4882 6554
rect 4934 6502 4946 6554
rect 4998 6502 5010 6554
rect 5062 6502 5074 6554
rect 5126 6502 5138 6554
rect 5190 6502 8815 6554
rect 8867 6502 8879 6554
rect 8931 6502 8943 6554
rect 8995 6502 9007 6554
rect 9059 6502 9071 6554
rect 9123 6502 12748 6554
rect 12800 6502 12812 6554
rect 12864 6502 12876 6554
rect 12928 6502 12940 6554
rect 12992 6502 13004 6554
rect 13056 6502 16681 6554
rect 16733 6502 16745 6554
rect 16797 6502 16809 6554
rect 16861 6502 16873 6554
rect 16925 6502 16937 6554
rect 16989 6502 16995 6554
rect 1104 6480 16995 6502
rect 1670 6440 1676 6452
rect 1631 6412 1676 6440
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 2314 6440 2320 6452
rect 2275 6412 2320 6440
rect 2314 6400 2320 6412
rect 2372 6400 2378 6452
rect 3326 6400 3332 6452
rect 3384 6440 3390 6452
rect 3421 6443 3479 6449
rect 3421 6440 3433 6443
rect 3384 6412 3433 6440
rect 3384 6400 3390 6412
rect 3421 6409 3433 6412
rect 3467 6409 3479 6443
rect 4798 6440 4804 6452
rect 3421 6403 3479 6409
rect 3528 6412 4804 6440
rect 1854 6304 1860 6316
rect 1815 6276 1860 6304
rect 1854 6264 1860 6276
rect 1912 6264 1918 6316
rect 2406 6264 2412 6316
rect 2464 6304 2470 6316
rect 2501 6307 2559 6313
rect 2501 6304 2513 6307
rect 2464 6276 2513 6304
rect 2464 6264 2470 6276
rect 2501 6273 2513 6276
rect 2547 6273 2559 6307
rect 2682 6304 2688 6316
rect 2643 6276 2688 6304
rect 2501 6267 2559 6273
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3528 6313 3556 6412
rect 4798 6400 4804 6412
rect 4856 6440 4862 6452
rect 6638 6440 6644 6452
rect 4856 6412 6644 6440
rect 4856 6400 4862 6412
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 6825 6443 6883 6449
rect 6825 6409 6837 6443
rect 6871 6440 6883 6443
rect 8570 6440 8576 6452
rect 6871 6412 8432 6440
rect 8531 6412 8576 6440
rect 6871 6409 6883 6412
rect 6825 6403 6883 6409
rect 4430 6332 4436 6384
rect 4488 6332 4494 6384
rect 5442 6372 5448 6384
rect 5403 6344 5448 6372
rect 5442 6332 5448 6344
rect 5500 6332 5506 6384
rect 7650 6372 7656 6384
rect 7611 6344 7656 6372
rect 7650 6332 7656 6344
rect 7708 6332 7714 6384
rect 7742 6332 7748 6384
rect 7800 6372 7806 6384
rect 7929 6375 7987 6381
rect 7929 6372 7941 6375
rect 7800 6344 7941 6372
rect 7800 6332 7806 6344
rect 7929 6341 7941 6344
rect 7975 6341 7987 6375
rect 8404 6372 8432 6412
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 10134 6440 10140 6452
rect 9140 6412 10140 6440
rect 8404 6344 8984 6372
rect 7929 6335 7987 6341
rect 3513 6307 3571 6313
rect 2832 6276 2877 6304
rect 2832 6264 2838 6276
rect 3513 6273 3525 6307
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 5721 6307 5779 6313
rect 5721 6273 5733 6307
rect 5767 6304 5779 6307
rect 6086 6304 6092 6316
rect 5767 6276 6092 6304
rect 5767 6273 5779 6276
rect 5721 6267 5779 6273
rect 6086 6264 6092 6276
rect 6144 6304 6150 6316
rect 6638 6304 6644 6316
rect 6144 6276 6644 6304
rect 6144 6264 6150 6276
rect 6638 6264 6644 6276
rect 6696 6264 6702 6316
rect 7190 6304 7196 6316
rect 7151 6276 7196 6304
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6304 7619 6307
rect 8036 6304 8248 6310
rect 8478 6304 8484 6316
rect 7607 6302 7880 6304
rect 7944 6302 8484 6304
rect 7607 6282 8484 6302
rect 7607 6276 8064 6282
rect 8220 6276 8484 6282
rect 7607 6273 7619 6276
rect 7852 6274 7972 6276
rect 7561 6267 7619 6273
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 3973 6239 4031 6245
rect 3973 6205 3985 6239
rect 4019 6236 4031 6239
rect 5350 6236 5356 6248
rect 4019 6208 5356 6236
rect 4019 6205 4031 6208
rect 3973 6199 4031 6205
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 7650 6196 7656 6248
rect 7708 6196 7714 6248
rect 8849 6239 8907 6245
rect 8849 6236 8861 6239
rect 8142 6208 8861 6236
rect 8849 6205 8861 6208
rect 8895 6205 8907 6239
rect 8956 6236 8984 6344
rect 9140 6313 9168 6412
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 11146 6400 11152 6452
rect 11204 6440 11210 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11204 6412 11805 6440
rect 11204 6400 11210 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 11793 6403 11851 6409
rect 9582 6332 9588 6384
rect 9640 6372 9646 6384
rect 9640 6344 11928 6372
rect 9640 6332 9646 6344
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 9306 6264 9312 6316
rect 9364 6304 9370 6316
rect 9858 6304 9864 6316
rect 9364 6276 9864 6304
rect 9364 6264 9370 6276
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 10612 6313 10640 6344
rect 10413 6307 10471 6313
rect 10413 6304 10425 6307
rect 9968 6276 10425 6304
rect 9324 6236 9352 6264
rect 8956 6208 9352 6236
rect 8849 6199 8907 6205
rect 8386 6128 8392 6180
rect 8444 6168 8450 6180
rect 9968 6168 9996 6276
rect 10413 6273 10425 6276
rect 10459 6273 10471 6307
rect 10413 6267 10471 6273
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6273 10655 6307
rect 11698 6304 11704 6316
rect 11611 6276 11704 6304
rect 10597 6267 10655 6273
rect 10428 6236 10456 6267
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 11900 6313 11928 6344
rect 11885 6307 11943 6313
rect 11885 6273 11897 6307
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 11716 6236 11744 6264
rect 10428 6208 11744 6236
rect 8444 6140 9996 6168
rect 8444 6128 8450 6140
rect 10502 6128 10508 6180
rect 10560 6168 10566 6180
rect 10689 6171 10747 6177
rect 10689 6168 10701 6171
rect 10560 6140 10701 6168
rect 10560 6128 10566 6140
rect 10689 6137 10701 6140
rect 10735 6137 10747 6171
rect 10689 6131 10747 6137
rect 4246 6060 4252 6112
rect 4304 6100 4310 6112
rect 6641 6103 6699 6109
rect 6641 6100 6653 6103
rect 4304 6072 6653 6100
rect 4304 6060 4310 6072
rect 6641 6069 6653 6072
rect 6687 6069 6699 6103
rect 6641 6063 6699 6069
rect 8478 6060 8484 6112
rect 8536 6100 8542 6112
rect 8757 6103 8815 6109
rect 8757 6100 8769 6103
rect 8536 6072 8769 6100
rect 8536 6060 8542 6072
rect 8757 6069 8769 6072
rect 8803 6069 8815 6103
rect 8757 6063 8815 6069
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 9677 6103 9735 6109
rect 9677 6100 9689 6103
rect 9548 6072 9689 6100
rect 9548 6060 9554 6072
rect 9677 6069 9689 6072
rect 9723 6069 9735 6103
rect 9677 6063 9735 6069
rect 1104 6010 16836 6032
rect 1104 5958 2916 6010
rect 2968 5958 2980 6010
rect 3032 5958 3044 6010
rect 3096 5958 3108 6010
rect 3160 5958 3172 6010
rect 3224 5958 6849 6010
rect 6901 5958 6913 6010
rect 6965 5958 6977 6010
rect 7029 5958 7041 6010
rect 7093 5958 7105 6010
rect 7157 5958 10782 6010
rect 10834 5958 10846 6010
rect 10898 5958 10910 6010
rect 10962 5958 10974 6010
rect 11026 5958 11038 6010
rect 11090 5958 14715 6010
rect 14767 5958 14779 6010
rect 14831 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 16836 6010
rect 1104 5936 16836 5958
rect 4706 5856 4712 5908
rect 4764 5896 4770 5908
rect 7009 5899 7067 5905
rect 7009 5896 7021 5899
rect 4764 5868 7021 5896
rect 4764 5856 4770 5868
rect 7009 5865 7021 5868
rect 7055 5896 7067 5899
rect 7190 5896 7196 5908
rect 7055 5868 7196 5896
rect 7055 5865 7067 5868
rect 7009 5859 7067 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 11238 5896 11244 5908
rect 11199 5868 11244 5896
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 2041 5831 2099 5837
rect 2041 5797 2053 5831
rect 2087 5828 2099 5831
rect 2314 5828 2320 5840
rect 2087 5800 2320 5828
rect 2087 5797 2099 5800
rect 2041 5791 2099 5797
rect 2314 5788 2320 5800
rect 2372 5788 2378 5840
rect 2498 5788 2504 5840
rect 2556 5828 2562 5840
rect 2682 5828 2688 5840
rect 2556 5800 2688 5828
rect 2556 5788 2562 5800
rect 2682 5788 2688 5800
rect 2740 5828 2746 5840
rect 2740 5800 3096 5828
rect 2740 5788 2746 5800
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5760 2007 5763
rect 2590 5760 2596 5772
rect 1995 5732 2596 5760
rect 1995 5729 2007 5732
rect 1949 5723 2007 5729
rect 2590 5720 2596 5732
rect 2648 5720 2654 5772
rect 2958 5760 2964 5772
rect 2700 5732 2964 5760
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 2222 5692 2228 5704
rect 2179 5664 2228 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 1872 5624 1900 5655
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 2700 5624 2728 5732
rect 2958 5720 2964 5732
rect 3016 5720 3022 5772
rect 2774 5652 2780 5704
rect 2832 5692 2838 5704
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 2832 5664 2881 5692
rect 2832 5652 2838 5664
rect 2869 5661 2881 5664
rect 2915 5692 2927 5695
rect 2915 5664 3004 5692
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 1872 5596 2728 5624
rect 1673 5559 1731 5565
rect 1673 5525 1685 5559
rect 1719 5556 1731 5559
rect 1854 5556 1860 5568
rect 1719 5528 1860 5556
rect 1719 5525 1731 5528
rect 1673 5519 1731 5525
rect 1854 5516 1860 5528
rect 1912 5516 1918 5568
rect 2682 5556 2688 5568
rect 2643 5528 2688 5556
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 2976 5556 3004 5664
rect 3068 5633 3096 5800
rect 6638 5788 6644 5840
rect 6696 5828 6702 5840
rect 8386 5828 8392 5840
rect 6696 5800 8392 5828
rect 6696 5788 6702 5800
rect 4430 5760 4436 5772
rect 4391 5732 4436 5760
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 5534 5760 5540 5772
rect 4632 5732 5540 5760
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5692 3203 5695
rect 3602 5692 3608 5704
rect 3191 5664 3608 5692
rect 3191 5661 3203 5664
rect 3145 5655 3203 5661
rect 3602 5652 3608 5664
rect 3660 5652 3666 5704
rect 4632 5701 4660 5732
rect 5534 5720 5540 5732
rect 5592 5760 5598 5772
rect 6730 5760 6736 5772
rect 5592 5732 6736 5760
rect 5592 5720 5598 5732
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5661 4675 5695
rect 4798 5692 4804 5704
rect 4759 5664 4804 5692
rect 4617 5655 4675 5661
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5661 5319 5695
rect 5261 5655 5319 5661
rect 3053 5627 3111 5633
rect 3053 5593 3065 5627
rect 3099 5624 3111 5627
rect 4246 5624 4252 5636
rect 3099 5596 4252 5624
rect 3099 5593 3111 5596
rect 3053 5587 3111 5593
rect 4246 5584 4252 5596
rect 4304 5584 4310 5636
rect 3326 5556 3332 5568
rect 2976 5528 3332 5556
rect 3326 5516 3332 5528
rect 3384 5516 3390 5568
rect 5276 5556 5304 5655
rect 6638 5652 6644 5704
rect 6696 5652 6702 5704
rect 8312 5701 8340 5800
rect 8386 5788 8392 5800
rect 8444 5788 8450 5840
rect 9490 5760 9496 5772
rect 9451 5732 9496 5760
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 9766 5760 9772 5772
rect 9727 5732 9772 5760
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5661 7803 5695
rect 7745 5655 7803 5661
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 9398 5692 9404 5704
rect 8527 5664 9404 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 5534 5624 5540 5636
rect 5495 5596 5540 5624
rect 5534 5584 5540 5596
rect 5592 5584 5598 5636
rect 7760 5624 7788 5655
rect 9398 5652 9404 5664
rect 9456 5652 9462 5704
rect 7760 5596 10180 5624
rect 10152 5568 10180 5596
rect 10502 5584 10508 5636
rect 10560 5584 10566 5636
rect 5626 5556 5632 5568
rect 5276 5528 5632 5556
rect 5626 5516 5632 5528
rect 5684 5516 5690 5568
rect 7558 5556 7564 5568
rect 7519 5528 7564 5556
rect 7558 5516 7564 5528
rect 7616 5516 7622 5568
rect 8478 5556 8484 5568
rect 8439 5528 8484 5556
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 10134 5516 10140 5568
rect 10192 5516 10198 5568
rect 1104 5466 16995 5488
rect 1104 5414 4882 5466
rect 4934 5414 4946 5466
rect 4998 5414 5010 5466
rect 5062 5414 5074 5466
rect 5126 5414 5138 5466
rect 5190 5414 8815 5466
rect 8867 5414 8879 5466
rect 8931 5414 8943 5466
rect 8995 5414 9007 5466
rect 9059 5414 9071 5466
rect 9123 5414 12748 5466
rect 12800 5414 12812 5466
rect 12864 5414 12876 5466
rect 12928 5414 12940 5466
rect 12992 5414 13004 5466
rect 13056 5414 16681 5466
rect 16733 5414 16745 5466
rect 16797 5414 16809 5466
rect 16861 5414 16873 5466
rect 16925 5414 16937 5466
rect 16989 5414 16995 5466
rect 1104 5392 16995 5414
rect 2222 5352 2228 5364
rect 1780 5324 2228 5352
rect 1780 5228 1808 5324
rect 2222 5312 2228 5324
rect 2280 5312 2286 5364
rect 3234 5312 3240 5364
rect 3292 5352 3298 5364
rect 3329 5355 3387 5361
rect 3329 5352 3341 5355
rect 3292 5324 3341 5352
rect 3292 5312 3298 5324
rect 3329 5321 3341 5324
rect 3375 5321 3387 5355
rect 3329 5315 3387 5321
rect 4614 5312 4620 5364
rect 4672 5352 4678 5364
rect 4893 5355 4951 5361
rect 4893 5352 4905 5355
rect 4672 5324 4905 5352
rect 4672 5312 4678 5324
rect 4893 5321 4905 5324
rect 4939 5321 4951 5355
rect 5626 5352 5632 5364
rect 5587 5324 5632 5352
rect 4893 5315 4951 5321
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 6638 5352 6644 5364
rect 6599 5324 6644 5352
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 10137 5355 10195 5361
rect 10137 5321 10149 5355
rect 10183 5352 10195 5355
rect 10318 5352 10324 5364
rect 10183 5324 10324 5352
rect 10183 5321 10195 5324
rect 10137 5315 10195 5321
rect 10318 5312 10324 5324
rect 10376 5312 10382 5364
rect 2130 5244 2136 5296
rect 2188 5284 2194 5296
rect 4157 5287 4215 5293
rect 2188 5256 3556 5284
rect 2188 5244 2194 5256
rect 1762 5216 1768 5228
rect 1723 5188 1768 5216
rect 1762 5176 1768 5188
rect 1820 5176 1826 5228
rect 2038 5216 2044 5228
rect 1999 5188 2044 5216
rect 2038 5176 2044 5188
rect 2096 5216 2102 5228
rect 2498 5216 2504 5228
rect 2096 5188 2504 5216
rect 2096 5176 2102 5188
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 2774 5216 2780 5228
rect 2731 5188 2780 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 2774 5176 2780 5188
rect 2832 5176 2838 5228
rect 3528 5225 3556 5256
rect 4157 5253 4169 5287
rect 4203 5284 4215 5287
rect 4246 5284 4252 5296
rect 4203 5256 4252 5284
rect 4203 5253 4215 5256
rect 4157 5247 4215 5253
rect 4246 5244 4252 5256
rect 4304 5244 4310 5296
rect 4338 5244 4344 5296
rect 4396 5284 4402 5296
rect 4396 5256 4441 5284
rect 4396 5244 4402 5256
rect 4798 5244 4804 5296
rect 4856 5284 4862 5296
rect 5258 5284 5264 5296
rect 4856 5256 5264 5284
rect 4856 5244 4862 5256
rect 5258 5244 5264 5256
rect 5316 5284 5322 5296
rect 7837 5287 7895 5293
rect 5316 5256 6592 5284
rect 5316 5244 5322 5256
rect 2869 5219 2927 5225
rect 2869 5185 2881 5219
rect 2915 5185 2927 5219
rect 2869 5179 2927 5185
rect 3513 5219 3571 5225
rect 3513 5185 3525 5219
rect 3559 5185 3571 5219
rect 3513 5179 3571 5185
rect 2314 5108 2320 5160
rect 2372 5148 2378 5160
rect 2884 5148 2912 5179
rect 4522 5176 4528 5228
rect 4580 5216 4586 5228
rect 4985 5219 5043 5225
rect 4985 5216 4997 5219
rect 4580 5188 4997 5216
rect 4580 5176 4586 5188
rect 4985 5185 4997 5188
rect 5031 5185 5043 5219
rect 4985 5179 5043 5185
rect 5350 5176 5356 5228
rect 5408 5216 5414 5228
rect 6564 5225 6592 5256
rect 7837 5253 7849 5287
rect 7883 5284 7895 5287
rect 8294 5284 8300 5296
rect 7883 5256 8300 5284
rect 7883 5253 7895 5256
rect 7837 5247 7895 5253
rect 8294 5244 8300 5256
rect 8352 5244 8358 5296
rect 9582 5284 9588 5296
rect 9543 5256 9588 5284
rect 9582 5244 9588 5256
rect 9640 5244 9646 5296
rect 5629 5219 5687 5225
rect 5629 5216 5641 5219
rect 5408 5188 5641 5216
rect 5408 5176 5414 5188
rect 5629 5185 5641 5188
rect 5675 5185 5687 5219
rect 5629 5179 5687 5185
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5185 6607 5219
rect 6730 5216 6736 5228
rect 6691 5188 6736 5216
rect 6549 5179 6607 5185
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 10045 5219 10103 5225
rect 10045 5185 10057 5219
rect 10091 5216 10103 5219
rect 10134 5216 10140 5228
rect 10091 5188 10140 5216
rect 10091 5185 10103 5188
rect 10045 5179 10103 5185
rect 10134 5176 10140 5188
rect 10192 5176 10198 5228
rect 4246 5148 4252 5160
rect 2372 5120 4252 5148
rect 2372 5108 2378 5120
rect 4246 5108 4252 5120
rect 4304 5148 4310 5160
rect 8018 5148 8024 5160
rect 4304 5120 8024 5148
rect 4304 5108 4310 5120
rect 8018 5108 8024 5120
rect 8076 5108 8082 5160
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 1670 5012 1676 5024
rect 1627 4984 1676 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 1670 4972 1676 4984
rect 1728 4972 1734 5024
rect 1949 5015 2007 5021
rect 1949 4981 1961 5015
rect 1995 5012 2007 5015
rect 2682 5012 2688 5024
rect 1995 4984 2688 5012
rect 1995 4981 2007 4984
rect 1949 4975 2007 4981
rect 2682 4972 2688 4984
rect 2740 4972 2746 5024
rect 3970 5012 3976 5024
rect 3931 4984 3976 5012
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 1104 4922 16836 4944
rect 1104 4870 2916 4922
rect 2968 4870 2980 4922
rect 3032 4870 3044 4922
rect 3096 4870 3108 4922
rect 3160 4870 3172 4922
rect 3224 4870 6849 4922
rect 6901 4870 6913 4922
rect 6965 4870 6977 4922
rect 7029 4870 7041 4922
rect 7093 4870 7105 4922
rect 7157 4870 10782 4922
rect 10834 4870 10846 4922
rect 10898 4870 10910 4922
rect 10962 4870 10974 4922
rect 11026 4870 11038 4922
rect 11090 4870 14715 4922
rect 14767 4870 14779 4922
rect 14831 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 16836 4922
rect 1104 4848 16836 4870
rect 1578 4768 1584 4820
rect 1636 4808 1642 4820
rect 3237 4811 3295 4817
rect 3237 4808 3249 4811
rect 1636 4780 3249 4808
rect 1636 4768 1642 4780
rect 3237 4777 3249 4780
rect 3283 4777 3295 4811
rect 3237 4771 3295 4777
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 3973 4811 4031 4817
rect 3973 4808 3985 4811
rect 3752 4780 3985 4808
rect 3752 4768 3758 4780
rect 3973 4777 3985 4780
rect 4019 4777 4031 4811
rect 5534 4808 5540 4820
rect 5495 4780 5540 4808
rect 3973 4771 4031 4777
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 9861 4811 9919 4817
rect 9861 4808 9873 4811
rect 9824 4780 9873 4808
rect 9824 4768 9830 4780
rect 9861 4777 9873 4780
rect 9907 4777 9919 4811
rect 9861 4771 9919 4777
rect 1486 4700 1492 4752
rect 1544 4740 1550 4752
rect 1673 4743 1731 4749
rect 1673 4740 1685 4743
rect 1544 4712 1685 4740
rect 1544 4700 1550 4712
rect 1673 4709 1685 4712
rect 1719 4709 1731 4743
rect 2590 4740 2596 4752
rect 2503 4712 2596 4740
rect 1673 4703 1731 4709
rect 2590 4700 2596 4712
rect 2648 4740 2654 4752
rect 3786 4740 3792 4752
rect 2648 4712 3792 4740
rect 2648 4700 2654 4712
rect 3786 4700 3792 4712
rect 3844 4700 3850 4752
rect 4709 4743 4767 4749
rect 4709 4709 4721 4743
rect 4755 4740 4767 4743
rect 5442 4740 5448 4752
rect 4755 4712 5448 4740
rect 4755 4709 4767 4712
rect 4709 4703 4767 4709
rect 5442 4700 5448 4712
rect 5500 4700 5506 4752
rect 2409 4675 2467 4681
rect 2409 4641 2421 4675
rect 2455 4672 2467 4675
rect 3050 4672 3056 4684
rect 2455 4644 3056 4672
rect 2455 4641 2467 4644
rect 2409 4635 2467 4641
rect 3050 4632 3056 4644
rect 3108 4632 3114 4684
rect 1854 4604 1860 4616
rect 1815 4576 1860 4604
rect 1854 4564 1860 4576
rect 1912 4564 1918 4616
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4573 2743 4607
rect 2685 4567 2743 4573
rect 3329 4607 3387 4613
rect 3329 4573 3341 4607
rect 3375 4604 3387 4607
rect 4062 4604 4068 4616
rect 3375 4576 4068 4604
rect 3375 4573 3387 4576
rect 3329 4567 3387 4573
rect 2314 4496 2320 4548
rect 2372 4536 2378 4548
rect 2700 4536 2728 4567
rect 4062 4564 4068 4576
rect 4120 4564 4126 4616
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4801 4607 4859 4613
rect 4212 4576 4257 4604
rect 4212 4564 4218 4576
rect 4801 4573 4813 4607
rect 4847 4604 4859 4607
rect 5258 4604 5264 4616
rect 4847 4576 5264 4604
rect 4847 4573 4859 4576
rect 4801 4567 4859 4573
rect 5258 4564 5264 4576
rect 5316 4564 5322 4616
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4573 5411 4607
rect 5353 4567 5411 4573
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4604 7711 4607
rect 9306 4604 9312 4616
rect 7699 4576 9312 4604
rect 7699 4573 7711 4576
rect 7653 4567 7711 4573
rect 2372 4508 2728 4536
rect 2372 4496 2378 4508
rect 4706 4496 4712 4548
rect 4764 4536 4770 4548
rect 5368 4536 5396 4567
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 9953 4607 10011 4613
rect 9953 4573 9965 4607
rect 9999 4604 10011 4607
rect 11238 4604 11244 4616
rect 9999 4576 11244 4604
rect 9999 4573 10011 4576
rect 9953 4567 10011 4573
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 7742 4536 7748 4548
rect 4764 4508 5396 4536
rect 7703 4508 7748 4536
rect 4764 4496 4770 4508
rect 7742 4496 7748 4508
rect 7800 4496 7806 4548
rect 1854 4428 1860 4480
rect 1912 4468 1918 4480
rect 2409 4471 2467 4477
rect 2409 4468 2421 4471
rect 1912 4440 2421 4468
rect 1912 4428 1918 4440
rect 2409 4437 2421 4440
rect 2455 4437 2467 4471
rect 2409 4431 2467 4437
rect 1104 4378 16995 4400
rect 1104 4326 4882 4378
rect 4934 4326 4946 4378
rect 4998 4326 5010 4378
rect 5062 4326 5074 4378
rect 5126 4326 5138 4378
rect 5190 4326 8815 4378
rect 8867 4326 8879 4378
rect 8931 4326 8943 4378
rect 8995 4326 9007 4378
rect 9059 4326 9071 4378
rect 9123 4326 12748 4378
rect 12800 4326 12812 4378
rect 12864 4326 12876 4378
rect 12928 4326 12940 4378
rect 12992 4326 13004 4378
rect 13056 4326 16681 4378
rect 16733 4326 16745 4378
rect 16797 4326 16809 4378
rect 16861 4326 16873 4378
rect 16925 4326 16937 4378
rect 16989 4326 16995 4378
rect 1104 4304 16995 4326
rect 4062 4264 4068 4276
rect 4023 4236 4068 4264
rect 4062 4224 4068 4236
rect 4120 4224 4126 4276
rect 3970 4196 3976 4208
rect 3252 4168 3976 4196
rect 1854 4128 1860 4140
rect 1815 4100 1860 4128
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 2784 4131 2842 4137
rect 2784 4097 2796 4131
rect 2830 4128 2842 4131
rect 3050 4128 3056 4140
rect 2830 4100 3056 4128
rect 2830 4097 2842 4100
rect 2784 4091 2842 4097
rect 3050 4088 3056 4100
rect 3108 4128 3114 4140
rect 3252 4128 3280 4168
rect 3970 4156 3976 4168
rect 4028 4156 4034 4208
rect 3510 4128 3516 4140
rect 3108 4100 3280 4128
rect 3471 4100 3516 4128
rect 3108 4088 3114 4100
rect 3510 4088 3516 4100
rect 3568 4088 3574 4140
rect 3605 4131 3663 4137
rect 3605 4097 3617 4131
rect 3651 4128 3663 4131
rect 4080 4128 4108 4224
rect 3651 4100 4108 4128
rect 4540 4168 4844 4196
rect 3651 4097 3663 4100
rect 3605 4091 3663 4097
rect 2498 4020 2504 4072
rect 2556 4060 2562 4072
rect 2869 4063 2927 4069
rect 2869 4060 2881 4063
rect 2556 4032 2881 4060
rect 2556 4020 2562 4032
rect 2869 4029 2881 4032
rect 2915 4029 2927 4063
rect 2869 4023 2927 4029
rect 2958 4020 2964 4072
rect 3016 4060 3022 4072
rect 4540 4060 4568 4168
rect 4816 4137 4844 4168
rect 7742 4156 7748 4208
rect 7800 4196 7806 4208
rect 7837 4199 7895 4205
rect 7837 4196 7849 4199
rect 7800 4168 7849 4196
rect 7800 4156 7806 4168
rect 7837 4165 7849 4168
rect 7883 4165 7895 4199
rect 7837 4159 7895 4165
rect 8478 4156 8484 4208
rect 8536 4156 8542 4208
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 4801 4131 4859 4137
rect 4801 4097 4813 4131
rect 4847 4097 4859 4131
rect 7558 4128 7564 4140
rect 7519 4100 7564 4128
rect 4801 4091 4859 4097
rect 3016 4032 4568 4060
rect 3016 4020 3022 4032
rect 2682 3952 2688 4004
rect 2740 3992 2746 4004
rect 4632 3992 4660 4091
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 9306 4060 9312 4072
rect 9267 4032 9312 4060
rect 9306 4020 9312 4032
rect 9364 4020 9370 4072
rect 2740 3964 4660 3992
rect 2740 3952 2746 3964
rect 1394 3884 1400 3936
rect 1452 3924 1458 3936
rect 1673 3927 1731 3933
rect 1673 3924 1685 3927
rect 1452 3896 1685 3924
rect 1452 3884 1458 3896
rect 1673 3893 1685 3896
rect 1719 3893 1731 3927
rect 1673 3887 1731 3893
rect 1854 3884 1860 3936
rect 1912 3924 1918 3936
rect 2409 3927 2467 3933
rect 2409 3924 2421 3927
rect 1912 3896 2421 3924
rect 1912 3884 1918 3896
rect 2409 3893 2421 3896
rect 2455 3893 2467 3927
rect 2409 3887 2467 3893
rect 3234 3884 3240 3936
rect 3292 3924 3298 3936
rect 4617 3927 4675 3933
rect 4617 3924 4629 3927
rect 3292 3896 4629 3924
rect 3292 3884 3298 3896
rect 4617 3893 4629 3896
rect 4663 3893 4675 3927
rect 4617 3887 4675 3893
rect 1104 3834 16836 3856
rect 1104 3782 2916 3834
rect 2968 3782 2980 3834
rect 3032 3782 3044 3834
rect 3096 3782 3108 3834
rect 3160 3782 3172 3834
rect 3224 3782 6849 3834
rect 6901 3782 6913 3834
rect 6965 3782 6977 3834
rect 7029 3782 7041 3834
rect 7093 3782 7105 3834
rect 7157 3782 10782 3834
rect 10834 3782 10846 3834
rect 10898 3782 10910 3834
rect 10962 3782 10974 3834
rect 11026 3782 11038 3834
rect 11090 3782 14715 3834
rect 14767 3782 14779 3834
rect 14831 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 16836 3834
rect 1104 3760 16836 3782
rect 1857 3723 1915 3729
rect 1857 3689 1869 3723
rect 1903 3720 1915 3723
rect 1946 3720 1952 3732
rect 1903 3692 1952 3720
rect 1903 3689 1915 3692
rect 1857 3683 1915 3689
rect 1946 3680 1952 3692
rect 2004 3680 2010 3732
rect 2774 3720 2780 3732
rect 2735 3692 2780 3720
rect 2774 3680 2780 3692
rect 2832 3680 2838 3732
rect 3786 3680 3792 3732
rect 3844 3720 3850 3732
rect 3973 3723 4031 3729
rect 3973 3720 3985 3723
rect 3844 3692 3985 3720
rect 3844 3680 3850 3692
rect 3973 3689 3985 3692
rect 4019 3689 4031 3723
rect 3973 3683 4031 3689
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 4617 3723 4675 3729
rect 4617 3720 4629 3723
rect 4120 3692 4629 3720
rect 4120 3680 4126 3692
rect 4617 3689 4629 3692
rect 4663 3689 4675 3723
rect 4617 3683 4675 3689
rect 3326 3652 3332 3664
rect 3287 3624 3332 3652
rect 3326 3612 3332 3624
rect 3384 3612 3390 3664
rect 3436 3556 4200 3584
rect 2038 3516 2044 3528
rect 1999 3488 2044 3516
rect 2038 3476 2044 3488
rect 2096 3476 2102 3528
rect 2406 3476 2412 3528
rect 2464 3516 2470 3528
rect 3436 3525 3464 3556
rect 4172 3525 4200 3556
rect 2593 3519 2651 3525
rect 2593 3516 2605 3519
rect 2464 3488 2605 3516
rect 2464 3476 2470 3488
rect 2593 3485 2605 3488
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3485 2835 3519
rect 2777 3479 2835 3485
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3516 4215 3519
rect 4338 3516 4344 3528
rect 4203 3488 4344 3516
rect 4203 3485 4215 3488
rect 4157 3479 4215 3485
rect 2792 3448 2820 3479
rect 3602 3448 3608 3460
rect 2792 3420 3608 3448
rect 3602 3408 3608 3420
rect 3660 3448 3666 3460
rect 3988 3448 4016 3479
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 3660 3420 4016 3448
rect 3660 3408 3666 3420
rect 1104 3290 16995 3312
rect 1104 3238 4882 3290
rect 4934 3238 4946 3290
rect 4998 3238 5010 3290
rect 5062 3238 5074 3290
rect 5126 3238 5138 3290
rect 5190 3238 8815 3290
rect 8867 3238 8879 3290
rect 8931 3238 8943 3290
rect 8995 3238 9007 3290
rect 9059 3238 9071 3290
rect 9123 3238 12748 3290
rect 12800 3238 12812 3290
rect 12864 3238 12876 3290
rect 12928 3238 12940 3290
rect 12992 3238 13004 3290
rect 13056 3238 16681 3290
rect 16733 3238 16745 3290
rect 16797 3238 16809 3290
rect 16861 3238 16873 3290
rect 16925 3238 16937 3290
rect 16989 3238 16995 3290
rect 1104 3216 16995 3238
rect 3418 3176 3424 3188
rect 3379 3148 3424 3176
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 1762 3068 1768 3120
rect 1820 3108 1826 3120
rect 4065 3111 4123 3117
rect 4065 3108 4077 3111
rect 1820 3080 4077 3108
rect 1820 3068 1826 3080
rect 4065 3077 4077 3080
rect 4111 3077 4123 3111
rect 4065 3071 4123 3077
rect 1854 3040 1860 3052
rect 1815 3012 1860 3040
rect 1854 3000 1860 3012
rect 1912 3000 1918 3052
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3040 3571 3043
rect 3602 3040 3608 3052
rect 3559 3012 3608 3040
rect 3559 3009 3571 3012
rect 3513 3003 3571 3009
rect 3602 3000 3608 3012
rect 3660 3000 3666 3052
rect 3970 3040 3976 3052
rect 3931 3012 3976 3040
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3040 4215 3043
rect 4246 3040 4252 3052
rect 4203 3012 4252 3040
rect 4203 3009 4215 3012
rect 4157 3003 4215 3009
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 1673 2839 1731 2845
rect 1673 2836 1685 2839
rect 1452 2808 1685 2836
rect 1452 2796 1458 2808
rect 1673 2805 1685 2808
rect 1719 2805 1731 2839
rect 1673 2799 1731 2805
rect 1104 2746 16836 2768
rect 1104 2694 2916 2746
rect 2968 2694 2980 2746
rect 3032 2694 3044 2746
rect 3096 2694 3108 2746
rect 3160 2694 3172 2746
rect 3224 2694 6849 2746
rect 6901 2694 6913 2746
rect 6965 2694 6977 2746
rect 7029 2694 7041 2746
rect 7093 2694 7105 2746
rect 7157 2694 10782 2746
rect 10834 2694 10846 2746
rect 10898 2694 10910 2746
rect 10962 2694 10974 2746
rect 11026 2694 11038 2746
rect 11090 2694 14715 2746
rect 14767 2694 14779 2746
rect 14831 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 16836 2746
rect 1104 2672 16836 2694
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2428 1639 2431
rect 1670 2428 1676 2440
rect 1627 2400 1676 2428
rect 1627 2397 1639 2400
rect 1581 2391 1639 2397
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 1762 2292 1768 2304
rect 1723 2264 1768 2292
rect 1762 2252 1768 2264
rect 1820 2252 1826 2304
rect 1104 2202 16995 2224
rect 1104 2150 4882 2202
rect 4934 2150 4946 2202
rect 4998 2150 5010 2202
rect 5062 2150 5074 2202
rect 5126 2150 5138 2202
rect 5190 2150 8815 2202
rect 8867 2150 8879 2202
rect 8931 2150 8943 2202
rect 8995 2150 9007 2202
rect 9059 2150 9071 2202
rect 9123 2150 12748 2202
rect 12800 2150 12812 2202
rect 12864 2150 12876 2202
rect 12928 2150 12940 2202
rect 12992 2150 13004 2202
rect 13056 2150 16681 2202
rect 16733 2150 16745 2202
rect 16797 2150 16809 2202
rect 16861 2150 16873 2202
rect 16925 2150 16937 2202
rect 16989 2150 16995 2202
rect 1104 2128 16995 2150
<< via1 >>
rect 4436 15852 4488 15904
rect 13912 15852 13964 15904
rect 2916 15750 2968 15802
rect 2980 15750 3032 15802
rect 3044 15750 3096 15802
rect 3108 15750 3160 15802
rect 3172 15750 3224 15802
rect 6849 15750 6901 15802
rect 6913 15750 6965 15802
rect 6977 15750 7029 15802
rect 7041 15750 7093 15802
rect 7105 15750 7157 15802
rect 10782 15750 10834 15802
rect 10846 15750 10898 15802
rect 10910 15750 10962 15802
rect 10974 15750 11026 15802
rect 11038 15750 11090 15802
rect 14715 15750 14767 15802
rect 14779 15750 14831 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 2780 15691 2832 15700
rect 2780 15657 2789 15691
rect 2789 15657 2823 15691
rect 2823 15657 2832 15691
rect 2780 15648 2832 15657
rect 4160 15648 4212 15700
rect 2044 15623 2096 15632
rect 2044 15589 2053 15623
rect 2053 15589 2087 15623
rect 2087 15589 2096 15623
rect 2044 15580 2096 15589
rect 4252 15623 4304 15632
rect 4252 15589 4261 15623
rect 4261 15589 4295 15623
rect 4295 15589 4304 15623
rect 4252 15580 4304 15589
rect 4436 15623 4488 15632
rect 4436 15589 4445 15623
rect 4445 15589 4479 15623
rect 4479 15589 4488 15623
rect 4436 15580 4488 15589
rect 5908 15580 5960 15632
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 2412 15376 2464 15428
rect 5540 15444 5592 15496
rect 5908 15487 5960 15496
rect 5908 15453 5917 15487
rect 5917 15453 5951 15487
rect 5951 15453 5960 15487
rect 5908 15444 5960 15453
rect 8300 15444 8352 15496
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 11336 15444 11388 15496
rect 12532 15487 12584 15496
rect 12532 15453 12541 15487
rect 12541 15453 12575 15487
rect 12575 15453 12584 15487
rect 12532 15444 12584 15453
rect 13820 15512 13872 15564
rect 14004 15444 14056 15496
rect 3240 15308 3292 15360
rect 6368 15376 6420 15428
rect 6552 15419 6604 15428
rect 6552 15385 6561 15419
rect 6561 15385 6595 15419
rect 6595 15385 6604 15419
rect 6552 15376 6604 15385
rect 8668 15376 8720 15428
rect 7840 15351 7892 15360
rect 7840 15317 7849 15351
rect 7849 15317 7883 15351
rect 7883 15317 7892 15351
rect 7840 15308 7892 15317
rect 9312 15351 9364 15360
rect 9312 15317 9321 15351
rect 9321 15317 9355 15351
rect 9355 15317 9364 15351
rect 9312 15308 9364 15317
rect 10232 15351 10284 15360
rect 10232 15317 10241 15351
rect 10241 15317 10275 15351
rect 10275 15317 10284 15351
rect 10232 15308 10284 15317
rect 10968 15351 11020 15360
rect 10968 15317 10977 15351
rect 10977 15317 11011 15351
rect 11011 15317 11020 15351
rect 10968 15308 11020 15317
rect 11060 15308 11112 15360
rect 13268 15308 13320 15360
rect 13820 15308 13872 15360
rect 4882 15206 4934 15258
rect 4946 15206 4998 15258
rect 5010 15206 5062 15258
rect 5074 15206 5126 15258
rect 5138 15206 5190 15258
rect 8815 15206 8867 15258
rect 8879 15206 8931 15258
rect 8943 15206 8995 15258
rect 9007 15206 9059 15258
rect 9071 15206 9123 15258
rect 12748 15206 12800 15258
rect 12812 15206 12864 15258
rect 12876 15206 12928 15258
rect 12940 15206 12992 15258
rect 13004 15206 13056 15258
rect 16681 15206 16733 15258
rect 16745 15206 16797 15258
rect 16809 15206 16861 15258
rect 16873 15206 16925 15258
rect 16937 15206 16989 15258
rect 2044 15147 2096 15156
rect 2044 15113 2053 15147
rect 2053 15113 2087 15147
rect 2087 15113 2096 15147
rect 2044 15104 2096 15113
rect 2412 15147 2464 15156
rect 2412 15113 2421 15147
rect 2421 15113 2455 15147
rect 2455 15113 2464 15147
rect 2412 15104 2464 15113
rect 6736 15036 6788 15088
rect 8668 15036 8720 15088
rect 2596 14943 2648 14952
rect 2596 14909 2605 14943
rect 2605 14909 2639 14943
rect 2639 14909 2648 14943
rect 6368 14968 6420 15020
rect 9312 15036 9364 15088
rect 10968 15036 11020 15088
rect 10416 14968 10468 15020
rect 11244 14968 11296 15020
rect 11336 14968 11388 15020
rect 2596 14900 2648 14909
rect 6460 14900 6512 14952
rect 8116 14900 8168 14952
rect 8300 14943 8352 14952
rect 8300 14909 8309 14943
rect 8309 14909 8343 14943
rect 8343 14909 8352 14943
rect 8300 14900 8352 14909
rect 9588 14900 9640 14952
rect 9772 14900 9824 14952
rect 10324 14900 10376 14952
rect 12440 14968 12492 15020
rect 13820 15011 13872 15020
rect 13820 14977 13829 15011
rect 13829 14977 13863 15011
rect 13863 14977 13872 15011
rect 13820 14968 13872 14977
rect 12532 14900 12584 14952
rect 13084 14900 13136 14952
rect 2964 14764 3016 14816
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 3608 14764 3660 14773
rect 3792 14764 3844 14816
rect 5632 14764 5684 14816
rect 10140 14764 10192 14816
rect 10968 14764 11020 14816
rect 11152 14764 11204 14816
rect 11796 14807 11848 14816
rect 11796 14773 11805 14807
rect 11805 14773 11839 14807
rect 11839 14773 11848 14807
rect 11796 14764 11848 14773
rect 12348 14764 12400 14816
rect 12624 14764 12676 14816
rect 15108 14764 15160 14816
rect 2916 14662 2968 14714
rect 2980 14662 3032 14714
rect 3044 14662 3096 14714
rect 3108 14662 3160 14714
rect 3172 14662 3224 14714
rect 6849 14662 6901 14714
rect 6913 14662 6965 14714
rect 6977 14662 7029 14714
rect 7041 14662 7093 14714
rect 7105 14662 7157 14714
rect 10782 14662 10834 14714
rect 10846 14662 10898 14714
rect 10910 14662 10962 14714
rect 10974 14662 11026 14714
rect 11038 14662 11090 14714
rect 14715 14662 14767 14714
rect 14779 14662 14831 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 2320 14560 2372 14612
rect 4252 14560 4304 14612
rect 8116 14603 8168 14612
rect 8116 14569 8125 14603
rect 8125 14569 8159 14603
rect 8159 14569 8168 14603
rect 8116 14560 8168 14569
rect 9588 14603 9640 14612
rect 9588 14569 9597 14603
rect 9597 14569 9631 14603
rect 9631 14569 9640 14603
rect 9588 14560 9640 14569
rect 11612 14560 11664 14612
rect 10140 14492 10192 14544
rect 5816 14424 5868 14476
rect 8300 14399 8352 14408
rect 8300 14365 8309 14399
rect 8309 14365 8343 14399
rect 8343 14365 8352 14399
rect 8300 14356 8352 14365
rect 9772 14399 9824 14408
rect 9772 14365 9781 14399
rect 9781 14365 9815 14399
rect 9815 14365 9824 14399
rect 9772 14356 9824 14365
rect 10232 14399 10284 14408
rect 10232 14365 10241 14399
rect 10241 14365 10275 14399
rect 10275 14365 10284 14399
rect 10232 14356 10284 14365
rect 3608 14288 3660 14340
rect 4712 14288 4764 14340
rect 5448 14288 5500 14340
rect 6460 14288 6512 14340
rect 11796 14288 11848 14340
rect 3332 14220 3384 14272
rect 6552 14263 6604 14272
rect 6552 14229 6561 14263
rect 6561 14229 6595 14263
rect 6595 14229 6604 14263
rect 6552 14220 6604 14229
rect 7380 14220 7432 14272
rect 10416 14220 10468 14272
rect 10876 14220 10928 14272
rect 11244 14220 11296 14272
rect 13084 14399 13136 14408
rect 13084 14365 13093 14399
rect 13093 14365 13127 14399
rect 13127 14365 13136 14399
rect 13084 14356 13136 14365
rect 11980 14263 12032 14272
rect 11980 14229 11989 14263
rect 11989 14229 12023 14263
rect 12023 14229 12032 14263
rect 12532 14263 12584 14272
rect 11980 14220 12032 14229
rect 12532 14229 12541 14263
rect 12541 14229 12575 14263
rect 12575 14229 12584 14263
rect 12532 14220 12584 14229
rect 13176 14263 13228 14272
rect 13176 14229 13185 14263
rect 13185 14229 13219 14263
rect 13219 14229 13228 14263
rect 13176 14220 13228 14229
rect 15108 14220 15160 14272
rect 4882 14118 4934 14170
rect 4946 14118 4998 14170
rect 5010 14118 5062 14170
rect 5074 14118 5126 14170
rect 5138 14118 5190 14170
rect 8815 14118 8867 14170
rect 8879 14118 8931 14170
rect 8943 14118 8995 14170
rect 9007 14118 9059 14170
rect 9071 14118 9123 14170
rect 12748 14118 12800 14170
rect 12812 14118 12864 14170
rect 12876 14118 12928 14170
rect 12940 14118 12992 14170
rect 13004 14118 13056 14170
rect 16681 14118 16733 14170
rect 16745 14118 16797 14170
rect 16809 14118 16861 14170
rect 16873 14118 16925 14170
rect 16937 14118 16989 14170
rect 1676 14059 1728 14068
rect 1676 14025 1685 14059
rect 1685 14025 1719 14059
rect 1719 14025 1728 14059
rect 1676 14016 1728 14025
rect 2780 14016 2832 14068
rect 3332 14016 3384 14068
rect 5356 14016 5408 14068
rect 5448 14016 5500 14068
rect 6736 14016 6788 14068
rect 11336 14016 11388 14068
rect 11612 14016 11664 14068
rect 11888 14016 11940 14068
rect 14556 14016 14608 14068
rect 4068 13948 4120 14000
rect 13176 13948 13228 14000
rect 3792 13923 3844 13932
rect 3792 13889 3801 13923
rect 3801 13889 3835 13923
rect 3835 13889 3844 13923
rect 3792 13880 3844 13889
rect 6092 13880 6144 13932
rect 7380 13923 7432 13932
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 9680 13880 9732 13932
rect 9772 13880 9824 13932
rect 7840 13812 7892 13864
rect 10324 13812 10376 13864
rect 11244 13880 11296 13932
rect 11796 13923 11848 13932
rect 11796 13889 11805 13923
rect 11805 13889 11839 13923
rect 11839 13889 11848 13923
rect 11796 13880 11848 13889
rect 12716 13923 12768 13932
rect 12716 13889 12725 13923
rect 12725 13889 12759 13923
rect 12759 13889 12768 13923
rect 12716 13880 12768 13889
rect 13636 13923 13688 13932
rect 13636 13889 13645 13923
rect 13645 13889 13679 13923
rect 13679 13889 13688 13923
rect 13636 13880 13688 13889
rect 10692 13812 10744 13864
rect 4620 13676 4672 13728
rect 6092 13676 6144 13728
rect 6736 13676 6788 13728
rect 7748 13676 7800 13728
rect 10416 13676 10468 13728
rect 13268 13744 13320 13796
rect 11060 13676 11112 13728
rect 12348 13676 12400 13728
rect 13084 13676 13136 13728
rect 13176 13676 13228 13728
rect 13820 13676 13872 13728
rect 2916 13574 2968 13626
rect 2980 13574 3032 13626
rect 3044 13574 3096 13626
rect 3108 13574 3160 13626
rect 3172 13574 3224 13626
rect 6849 13574 6901 13626
rect 6913 13574 6965 13626
rect 6977 13574 7029 13626
rect 7041 13574 7093 13626
rect 7105 13574 7157 13626
rect 10782 13574 10834 13626
rect 10846 13574 10898 13626
rect 10910 13574 10962 13626
rect 10974 13574 11026 13626
rect 11038 13574 11090 13626
rect 14715 13574 14767 13626
rect 14779 13574 14831 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 4804 13472 4856 13524
rect 10600 13472 10652 13524
rect 11060 13472 11112 13524
rect 11796 13472 11848 13524
rect 14556 13472 14608 13524
rect 4620 13447 4672 13456
rect 4620 13413 4629 13447
rect 4629 13413 4663 13447
rect 4663 13413 4672 13447
rect 4620 13404 4672 13413
rect 2320 13336 2372 13388
rect 2596 13379 2648 13388
rect 2596 13345 2605 13379
rect 2605 13345 2639 13379
rect 2639 13345 2648 13379
rect 2596 13336 2648 13345
rect 5724 13336 5776 13388
rect 7840 13336 7892 13388
rect 2044 13268 2096 13320
rect 2780 13311 2832 13320
rect 2780 13277 2789 13311
rect 2789 13277 2823 13311
rect 2823 13277 2832 13311
rect 2780 13268 2832 13277
rect 3332 13268 3384 13320
rect 4804 13268 4856 13320
rect 6736 13268 6788 13320
rect 11152 13404 11204 13456
rect 1676 13175 1728 13184
rect 1676 13141 1685 13175
rect 1685 13141 1719 13175
rect 1719 13141 1728 13175
rect 1676 13132 1728 13141
rect 3148 13175 3200 13184
rect 3148 13141 3157 13175
rect 3157 13141 3191 13175
rect 3191 13141 3200 13175
rect 3148 13132 3200 13141
rect 5632 13200 5684 13252
rect 7104 13243 7156 13252
rect 6736 13132 6788 13184
rect 7104 13209 7113 13243
rect 7113 13209 7147 13243
rect 7147 13209 7156 13243
rect 7104 13200 7156 13209
rect 7748 13132 7800 13184
rect 7840 13132 7892 13184
rect 12440 13336 12492 13388
rect 13912 13336 13964 13388
rect 8484 13132 8536 13184
rect 10968 13268 11020 13320
rect 9312 13175 9364 13184
rect 9312 13141 9321 13175
rect 9321 13141 9355 13175
rect 9355 13141 9364 13175
rect 9312 13132 9364 13141
rect 12532 13268 12584 13320
rect 13636 13311 13688 13320
rect 13636 13277 13645 13311
rect 13645 13277 13679 13311
rect 13679 13277 13688 13311
rect 13636 13268 13688 13277
rect 14464 13311 14516 13320
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 11428 13243 11480 13252
rect 11428 13209 11437 13243
rect 11437 13209 11471 13243
rect 11471 13209 11480 13243
rect 11428 13200 11480 13209
rect 12440 13132 12492 13184
rect 12716 13132 12768 13184
rect 14188 13132 14240 13184
rect 14280 13132 14332 13184
rect 4882 13030 4934 13082
rect 4946 13030 4998 13082
rect 5010 13030 5062 13082
rect 5074 13030 5126 13082
rect 5138 13030 5190 13082
rect 8815 13030 8867 13082
rect 8879 13030 8931 13082
rect 8943 13030 8995 13082
rect 9007 13030 9059 13082
rect 9071 13030 9123 13082
rect 12748 13030 12800 13082
rect 12812 13030 12864 13082
rect 12876 13030 12928 13082
rect 12940 13030 12992 13082
rect 13004 13030 13056 13082
rect 16681 13030 16733 13082
rect 16745 13030 16797 13082
rect 16809 13030 16861 13082
rect 16873 13030 16925 13082
rect 16937 13030 16989 13082
rect 2412 12928 2464 12980
rect 3240 12860 3292 12912
rect 2044 12835 2096 12844
rect 2044 12801 2053 12835
rect 2053 12801 2087 12835
rect 2087 12801 2096 12835
rect 2044 12792 2096 12801
rect 4068 12835 4120 12844
rect 4068 12801 4077 12835
rect 4077 12801 4111 12835
rect 4111 12801 4120 12835
rect 4068 12792 4120 12801
rect 13820 12928 13872 12980
rect 14096 12928 14148 12980
rect 5816 12860 5868 12912
rect 7104 12860 7156 12912
rect 4804 12835 4856 12844
rect 4804 12801 4838 12835
rect 4838 12801 4856 12835
rect 4804 12792 4856 12801
rect 5080 12792 5132 12844
rect 2320 12767 2372 12776
rect 2320 12733 2329 12767
rect 2329 12733 2363 12767
rect 2363 12733 2372 12767
rect 2320 12724 2372 12733
rect 3148 12699 3200 12708
rect 3148 12665 3157 12699
rect 3157 12665 3191 12699
rect 3191 12665 3200 12699
rect 3148 12656 3200 12665
rect 4528 12656 4580 12708
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 5632 12588 5684 12640
rect 6736 12792 6788 12844
rect 8024 12792 8076 12844
rect 8484 12835 8536 12844
rect 8484 12801 8493 12835
rect 8493 12801 8527 12835
rect 8527 12801 8536 12835
rect 8484 12792 8536 12801
rect 9312 12860 9364 12912
rect 10692 12860 10744 12912
rect 11428 12860 11480 12912
rect 12440 12792 12492 12844
rect 13084 12860 13136 12912
rect 13176 12903 13228 12912
rect 13176 12869 13185 12903
rect 13185 12869 13219 12903
rect 13219 12869 13228 12903
rect 13176 12860 13228 12869
rect 14280 12792 14332 12844
rect 10600 12724 10652 12776
rect 13636 12724 13688 12776
rect 7196 12588 7248 12640
rect 2916 12486 2968 12538
rect 2980 12486 3032 12538
rect 3044 12486 3096 12538
rect 3108 12486 3160 12538
rect 3172 12486 3224 12538
rect 6849 12486 6901 12538
rect 6913 12486 6965 12538
rect 6977 12486 7029 12538
rect 7041 12486 7093 12538
rect 7105 12486 7157 12538
rect 10782 12486 10834 12538
rect 10846 12486 10898 12538
rect 10910 12486 10962 12538
rect 10974 12486 11026 12538
rect 11038 12486 11090 12538
rect 14715 12486 14767 12538
rect 14779 12486 14831 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 2044 12384 2096 12436
rect 12532 12316 12584 12368
rect 5908 12180 5960 12232
rect 10600 12180 10652 12232
rect 3240 12112 3292 12164
rect 4252 12155 4304 12164
rect 4252 12121 4261 12155
rect 4261 12121 4295 12155
rect 4295 12121 4304 12155
rect 4252 12112 4304 12121
rect 7288 12112 7340 12164
rect 10232 12112 10284 12164
rect 11244 12112 11296 12164
rect 13360 12180 13412 12232
rect 14464 12223 14516 12232
rect 14464 12189 14473 12223
rect 14473 12189 14507 12223
rect 14507 12189 14516 12223
rect 14464 12180 14516 12189
rect 15108 12223 15160 12232
rect 15108 12189 15117 12223
rect 15117 12189 15151 12223
rect 15151 12189 15160 12223
rect 15108 12180 15160 12189
rect 12624 12112 12676 12164
rect 7196 12044 7248 12096
rect 8024 12087 8076 12096
rect 8024 12053 8033 12087
rect 8033 12053 8067 12087
rect 8067 12053 8076 12087
rect 8024 12044 8076 12053
rect 9680 12044 9732 12096
rect 12440 12044 12492 12096
rect 13912 12044 13964 12096
rect 14372 12087 14424 12096
rect 14372 12053 14381 12087
rect 14381 12053 14415 12087
rect 14415 12053 14424 12087
rect 14372 12044 14424 12053
rect 4882 11942 4934 11994
rect 4946 11942 4998 11994
rect 5010 11942 5062 11994
rect 5074 11942 5126 11994
rect 5138 11942 5190 11994
rect 8815 11942 8867 11994
rect 8879 11942 8931 11994
rect 8943 11942 8995 11994
rect 9007 11942 9059 11994
rect 9071 11942 9123 11994
rect 12748 11942 12800 11994
rect 12812 11942 12864 11994
rect 12876 11942 12928 11994
rect 12940 11942 12992 11994
rect 13004 11942 13056 11994
rect 16681 11942 16733 11994
rect 16745 11942 16797 11994
rect 16809 11942 16861 11994
rect 16873 11942 16925 11994
rect 16937 11942 16989 11994
rect 1676 11772 1728 11824
rect 5264 11840 5316 11892
rect 5908 11883 5960 11892
rect 5908 11849 5917 11883
rect 5917 11849 5951 11883
rect 5951 11849 5960 11883
rect 5908 11840 5960 11849
rect 7288 11883 7340 11892
rect 4436 11772 4488 11824
rect 7288 11849 7297 11883
rect 7297 11849 7331 11883
rect 7331 11849 7340 11883
rect 7288 11840 7340 11849
rect 8116 11840 8168 11892
rect 13360 11840 13412 11892
rect 2136 11500 2188 11552
rect 2688 11636 2740 11688
rect 4068 11636 4120 11688
rect 5908 11704 5960 11756
rect 3148 11500 3200 11552
rect 5264 11500 5316 11552
rect 6736 11568 6788 11620
rect 7656 11704 7708 11756
rect 8024 11747 8076 11756
rect 8024 11713 8033 11747
rect 8033 11713 8067 11747
rect 8067 11713 8076 11747
rect 8024 11704 8076 11713
rect 9220 11747 9272 11756
rect 9220 11713 9229 11747
rect 9229 11713 9263 11747
rect 9263 11713 9272 11747
rect 9220 11704 9272 11713
rect 9588 11704 9640 11756
rect 14004 11772 14056 11824
rect 14372 11772 14424 11824
rect 9496 11636 9548 11688
rect 14188 11636 14240 11688
rect 8300 11568 8352 11620
rect 13268 11568 13320 11620
rect 9588 11500 9640 11552
rect 10416 11500 10468 11552
rect 13636 11543 13688 11552
rect 13636 11509 13645 11543
rect 13645 11509 13679 11543
rect 13679 11509 13688 11543
rect 13636 11500 13688 11509
rect 2916 11398 2968 11450
rect 2980 11398 3032 11450
rect 3044 11398 3096 11450
rect 3108 11398 3160 11450
rect 3172 11398 3224 11450
rect 6849 11398 6901 11450
rect 6913 11398 6965 11450
rect 6977 11398 7029 11450
rect 7041 11398 7093 11450
rect 7105 11398 7157 11450
rect 10782 11398 10834 11450
rect 10846 11398 10898 11450
rect 10910 11398 10962 11450
rect 10974 11398 11026 11450
rect 11038 11398 11090 11450
rect 14715 11398 14767 11450
rect 14779 11398 14831 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 2688 11339 2740 11348
rect 2688 11305 2697 11339
rect 2697 11305 2731 11339
rect 2731 11305 2740 11339
rect 2688 11296 2740 11305
rect 5632 11339 5684 11348
rect 5632 11305 5662 11339
rect 5662 11305 5684 11339
rect 9220 11339 9272 11348
rect 5632 11296 5684 11305
rect 1676 11271 1728 11280
rect 1676 11237 1685 11271
rect 1685 11237 1719 11271
rect 1719 11237 1728 11271
rect 1676 11228 1728 11237
rect 4436 11228 4488 11280
rect 6736 11228 6788 11280
rect 7288 11228 7340 11280
rect 3332 11160 3384 11212
rect 6276 11160 6328 11212
rect 4068 11024 4120 11076
rect 4344 11092 4396 11144
rect 7656 11092 7708 11144
rect 9220 11305 9229 11339
rect 9229 11305 9263 11339
rect 9263 11305 9272 11339
rect 9220 11296 9272 11305
rect 10232 11339 10284 11348
rect 10232 11305 10241 11339
rect 10241 11305 10275 11339
rect 10275 11305 10284 11339
rect 10232 11296 10284 11305
rect 13452 11296 13504 11348
rect 13268 11271 13320 11280
rect 13268 11237 13277 11271
rect 13277 11237 13311 11271
rect 13311 11237 13320 11271
rect 13268 11228 13320 11237
rect 9312 11092 9364 11144
rect 9772 11160 9824 11212
rect 11244 11160 11296 11212
rect 11428 11160 11480 11212
rect 14464 11228 14516 11280
rect 9588 11135 9640 11144
rect 9588 11101 9597 11135
rect 9597 11101 9631 11135
rect 9631 11101 9640 11135
rect 9588 11092 9640 11101
rect 11152 11092 11204 11144
rect 12716 11135 12768 11144
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 13360 11135 13412 11144
rect 12716 11092 12768 11101
rect 13360 11101 13369 11135
rect 13369 11101 13403 11135
rect 13403 11101 13412 11135
rect 13360 11092 13412 11101
rect 13452 11092 13504 11144
rect 16120 11092 16172 11144
rect 4620 11024 4672 11076
rect 6368 11024 6420 11076
rect 4528 10956 4580 11008
rect 7748 10956 7800 11008
rect 7932 11024 7984 11076
rect 11060 10956 11112 11008
rect 12440 11067 12492 11076
rect 12440 11033 12449 11067
rect 12449 11033 12483 11067
rect 12483 11033 12492 11067
rect 12440 11024 12492 11033
rect 15660 11067 15712 11076
rect 15660 11033 15669 11067
rect 15669 11033 15703 11067
rect 15703 11033 15712 11067
rect 15660 11024 15712 11033
rect 13820 10956 13872 11008
rect 4882 10854 4934 10906
rect 4946 10854 4998 10906
rect 5010 10854 5062 10906
rect 5074 10854 5126 10906
rect 5138 10854 5190 10906
rect 8815 10854 8867 10906
rect 8879 10854 8931 10906
rect 8943 10854 8995 10906
rect 9007 10854 9059 10906
rect 9071 10854 9123 10906
rect 12748 10854 12800 10906
rect 12812 10854 12864 10906
rect 12876 10854 12928 10906
rect 12940 10854 12992 10906
rect 13004 10854 13056 10906
rect 16681 10854 16733 10906
rect 16745 10854 16797 10906
rect 16809 10854 16861 10906
rect 16873 10854 16925 10906
rect 16937 10854 16989 10906
rect 4068 10752 4120 10804
rect 7840 10795 7892 10804
rect 7840 10761 7849 10795
rect 7849 10761 7883 10795
rect 7883 10761 7892 10795
rect 7840 10752 7892 10761
rect 10324 10752 10376 10804
rect 4252 10727 4304 10736
rect 4252 10693 4261 10727
rect 4261 10693 4295 10727
rect 4295 10693 4304 10727
rect 4252 10684 4304 10693
rect 6552 10727 6604 10736
rect 6552 10693 6561 10727
rect 6561 10693 6595 10727
rect 6595 10693 6604 10727
rect 6552 10684 6604 10693
rect 10416 10684 10468 10736
rect 15660 10684 15712 10736
rect 9312 10548 9364 10600
rect 11060 10616 11112 10668
rect 11796 10616 11848 10668
rect 13912 10659 13964 10668
rect 13912 10625 13921 10659
rect 13921 10625 13955 10659
rect 13955 10625 13964 10659
rect 13912 10616 13964 10625
rect 16120 10659 16172 10668
rect 16120 10625 16129 10659
rect 16129 10625 16163 10659
rect 16163 10625 16172 10659
rect 16120 10616 16172 10625
rect 14188 10591 14240 10600
rect 14188 10557 14197 10591
rect 14197 10557 14231 10591
rect 14231 10557 14240 10591
rect 14188 10548 14240 10557
rect 13820 10480 13872 10532
rect 8300 10412 8352 10464
rect 9404 10412 9456 10464
rect 10324 10412 10376 10464
rect 11152 10412 11204 10464
rect 13544 10412 13596 10464
rect 16212 10455 16264 10464
rect 16212 10421 16221 10455
rect 16221 10421 16255 10455
rect 16255 10421 16264 10455
rect 16212 10412 16264 10421
rect 2916 10310 2968 10362
rect 2980 10310 3032 10362
rect 3044 10310 3096 10362
rect 3108 10310 3160 10362
rect 3172 10310 3224 10362
rect 6849 10310 6901 10362
rect 6913 10310 6965 10362
rect 6977 10310 7029 10362
rect 7041 10310 7093 10362
rect 7105 10310 7157 10362
rect 10782 10310 10834 10362
rect 10846 10310 10898 10362
rect 10910 10310 10962 10362
rect 10974 10310 11026 10362
rect 11038 10310 11090 10362
rect 14715 10310 14767 10362
rect 14779 10310 14831 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 4620 10208 4672 10260
rect 5356 10208 5408 10260
rect 5724 10251 5776 10260
rect 5724 10217 5733 10251
rect 5733 10217 5767 10251
rect 5767 10217 5776 10251
rect 5724 10208 5776 10217
rect 5908 10208 5960 10260
rect 11428 10208 11480 10260
rect 14188 10208 14240 10260
rect 4068 10140 4120 10192
rect 15108 10140 15160 10192
rect 7564 10115 7616 10124
rect 7564 10081 7573 10115
rect 7573 10081 7607 10115
rect 7607 10081 7616 10115
rect 7564 10072 7616 10081
rect 7748 10115 7800 10124
rect 7748 10081 7757 10115
rect 7757 10081 7791 10115
rect 7791 10081 7800 10115
rect 7748 10072 7800 10081
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 5264 10004 5316 10056
rect 9496 10072 9548 10124
rect 16120 10072 16172 10124
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 13636 10004 13688 10056
rect 1952 9936 2004 9988
rect 3332 9936 3384 9988
rect 4620 9936 4672 9988
rect 10416 9936 10468 9988
rect 3976 9911 4028 9920
rect 3976 9877 3985 9911
rect 3985 9877 4019 9911
rect 4019 9877 4028 9911
rect 3976 9868 4028 9877
rect 4528 9868 4580 9920
rect 8392 9868 8444 9920
rect 9404 9911 9456 9920
rect 9404 9877 9413 9911
rect 9413 9877 9447 9911
rect 9447 9877 9456 9911
rect 9404 9868 9456 9877
rect 14188 9868 14240 9920
rect 4882 9766 4934 9818
rect 4946 9766 4998 9818
rect 5010 9766 5062 9818
rect 5074 9766 5126 9818
rect 5138 9766 5190 9818
rect 8815 9766 8867 9818
rect 8879 9766 8931 9818
rect 8943 9766 8995 9818
rect 9007 9766 9059 9818
rect 9071 9766 9123 9818
rect 12748 9766 12800 9818
rect 12812 9766 12864 9818
rect 12876 9766 12928 9818
rect 12940 9766 12992 9818
rect 13004 9766 13056 9818
rect 16681 9766 16733 9818
rect 16745 9766 16797 9818
rect 16809 9766 16861 9818
rect 16873 9766 16925 9818
rect 16937 9766 16989 9818
rect 3332 9596 3384 9648
rect 4436 9596 4488 9648
rect 6368 9596 6420 9648
rect 5356 9528 5408 9580
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 5816 9528 5868 9537
rect 8300 9596 8352 9648
rect 9404 9596 9456 9648
rect 8116 9571 8168 9580
rect 4160 9460 4212 9512
rect 5080 9460 5132 9512
rect 5908 9435 5960 9444
rect 5908 9401 5917 9435
rect 5917 9401 5951 9435
rect 5951 9401 5960 9435
rect 5908 9392 5960 9401
rect 8116 9537 8125 9571
rect 8125 9537 8159 9571
rect 8159 9537 8168 9571
rect 8116 9528 8168 9537
rect 16212 9664 16264 9716
rect 15476 9596 15528 9648
rect 14188 9571 14240 9580
rect 7932 9460 7984 9512
rect 9588 9460 9640 9512
rect 14188 9537 14197 9571
rect 14197 9537 14231 9571
rect 14231 9537 14240 9571
rect 14188 9528 14240 9537
rect 13452 9503 13504 9512
rect 4528 9324 4580 9376
rect 4804 9324 4856 9376
rect 5264 9324 5316 9376
rect 11428 9392 11480 9444
rect 13452 9469 13461 9503
rect 13461 9469 13495 9503
rect 13495 9469 13504 9503
rect 13452 9460 13504 9469
rect 13728 9503 13780 9512
rect 13728 9469 13737 9503
rect 13737 9469 13771 9503
rect 13771 9469 13780 9503
rect 13728 9460 13780 9469
rect 15108 9460 15160 9512
rect 12348 9392 12400 9444
rect 6644 9324 6696 9376
rect 9864 9367 9916 9376
rect 9864 9333 9873 9367
rect 9873 9333 9907 9367
rect 9907 9333 9916 9367
rect 9864 9324 9916 9333
rect 15568 9324 15620 9376
rect 2916 9222 2968 9274
rect 2980 9222 3032 9274
rect 3044 9222 3096 9274
rect 3108 9222 3160 9274
rect 3172 9222 3224 9274
rect 6849 9222 6901 9274
rect 6913 9222 6965 9274
rect 6977 9222 7029 9274
rect 7041 9222 7093 9274
rect 7105 9222 7157 9274
rect 10782 9222 10834 9274
rect 10846 9222 10898 9274
rect 10910 9222 10962 9274
rect 10974 9222 11026 9274
rect 11038 9222 11090 9274
rect 14715 9222 14767 9274
rect 14779 9222 14831 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 7564 9120 7616 9172
rect 11796 9163 11848 9172
rect 3516 8916 3568 8968
rect 4252 9052 4304 9104
rect 5356 9052 5408 9104
rect 11796 9129 11805 9163
rect 11805 9129 11839 9163
rect 11839 9129 11848 9163
rect 11796 9120 11848 9129
rect 13452 9120 13504 9172
rect 15108 9163 15160 9172
rect 15108 9129 15117 9163
rect 15117 9129 15151 9163
rect 15151 9129 15160 9163
rect 15108 9120 15160 9129
rect 13728 9052 13780 9104
rect 4436 9027 4488 9036
rect 4436 8993 4445 9027
rect 4445 8993 4479 9027
rect 4479 8993 4488 9027
rect 4436 8984 4488 8993
rect 6276 8984 6328 9036
rect 6644 9027 6696 9036
rect 6644 8993 6653 9027
rect 6653 8993 6687 9027
rect 6687 8993 6696 9027
rect 6644 8984 6696 8993
rect 4344 8959 4396 8968
rect 4344 8925 4353 8959
rect 4353 8925 4387 8959
rect 4387 8925 4396 8959
rect 4344 8916 4396 8925
rect 5080 8916 5132 8968
rect 7472 8916 7524 8968
rect 9220 8916 9272 8968
rect 9864 8984 9916 9036
rect 10324 9027 10376 9036
rect 10324 8993 10333 9027
rect 10333 8993 10367 9027
rect 10367 8993 10376 9027
rect 10324 8984 10376 8993
rect 11336 8984 11388 9036
rect 11428 8916 11480 8968
rect 3700 8848 3752 8900
rect 5908 8848 5960 8900
rect 10232 8848 10284 8900
rect 12348 8916 12400 8968
rect 15568 8916 15620 8968
rect 16120 8916 16172 8968
rect 13268 8848 13320 8900
rect 2596 8780 2648 8832
rect 4528 8780 4580 8832
rect 5448 8780 5500 8832
rect 6092 8780 6144 8832
rect 14648 8780 14700 8832
rect 15844 8823 15896 8832
rect 15844 8789 15853 8823
rect 15853 8789 15887 8823
rect 15887 8789 15896 8823
rect 15844 8780 15896 8789
rect 4882 8678 4934 8730
rect 4946 8678 4998 8730
rect 5010 8678 5062 8730
rect 5074 8678 5126 8730
rect 5138 8678 5190 8730
rect 8815 8678 8867 8730
rect 8879 8678 8931 8730
rect 8943 8678 8995 8730
rect 9007 8678 9059 8730
rect 9071 8678 9123 8730
rect 12748 8678 12800 8730
rect 12812 8678 12864 8730
rect 12876 8678 12928 8730
rect 12940 8678 12992 8730
rect 13004 8678 13056 8730
rect 16681 8678 16733 8730
rect 16745 8678 16797 8730
rect 16809 8678 16861 8730
rect 16873 8678 16925 8730
rect 16937 8678 16989 8730
rect 1768 8619 1820 8628
rect 1768 8585 1777 8619
rect 1777 8585 1811 8619
rect 1811 8585 1820 8619
rect 1768 8576 1820 8585
rect 1492 8440 1544 8492
rect 2596 8440 2648 8492
rect 7932 8576 7984 8628
rect 15476 8619 15528 8628
rect 15476 8585 15485 8619
rect 15485 8585 15519 8619
rect 15519 8585 15528 8619
rect 15476 8576 15528 8585
rect 7564 8508 7616 8560
rect 9496 8508 9548 8560
rect 4160 8440 4212 8492
rect 4620 8372 4672 8424
rect 5356 8440 5408 8492
rect 5816 8440 5868 8492
rect 9772 8483 9824 8492
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 11244 8440 11296 8492
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 15844 8508 15896 8560
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 16120 8440 16172 8492
rect 7288 8415 7340 8424
rect 4436 8304 4488 8356
rect 5264 8304 5316 8356
rect 5816 8304 5868 8356
rect 7288 8381 7297 8415
rect 7297 8381 7331 8415
rect 7331 8381 7340 8415
rect 7288 8372 7340 8381
rect 14372 8415 14424 8424
rect 14372 8381 14381 8415
rect 14381 8381 14415 8415
rect 14415 8381 14424 8415
rect 14372 8372 14424 8381
rect 7472 8304 7524 8356
rect 6000 8236 6052 8288
rect 8300 8279 8352 8288
rect 8300 8245 8309 8279
rect 8309 8245 8343 8279
rect 8343 8245 8352 8279
rect 8300 8236 8352 8245
rect 11336 8304 11388 8356
rect 8484 8236 8536 8288
rect 12072 8236 12124 8288
rect 12900 8279 12952 8288
rect 12900 8245 12909 8279
rect 12909 8245 12943 8279
rect 12943 8245 12952 8279
rect 12900 8236 12952 8245
rect 2916 8134 2968 8186
rect 2980 8134 3032 8186
rect 3044 8134 3096 8186
rect 3108 8134 3160 8186
rect 3172 8134 3224 8186
rect 6849 8134 6901 8186
rect 6913 8134 6965 8186
rect 6977 8134 7029 8186
rect 7041 8134 7093 8186
rect 7105 8134 7157 8186
rect 10782 8134 10834 8186
rect 10846 8134 10898 8186
rect 10910 8134 10962 8186
rect 10974 8134 11026 8186
rect 11038 8134 11090 8186
rect 14715 8134 14767 8186
rect 14779 8134 14831 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 1768 8075 1820 8084
rect 1768 8041 1777 8075
rect 1777 8041 1811 8075
rect 1811 8041 1820 8075
rect 1768 8032 1820 8041
rect 9772 8032 9824 8084
rect 3792 7964 3844 8016
rect 4160 7964 4212 8016
rect 5724 7964 5776 8016
rect 9128 7964 9180 8016
rect 1676 7828 1728 7880
rect 3148 7828 3200 7880
rect 3884 7828 3936 7880
rect 4252 7871 4304 7880
rect 4252 7837 4261 7871
rect 4261 7837 4295 7871
rect 4295 7837 4304 7871
rect 4252 7828 4304 7837
rect 5448 7828 5500 7880
rect 8300 7896 8352 7948
rect 12348 8032 12400 8084
rect 14372 8032 14424 8084
rect 12072 7939 12124 7948
rect 4344 7760 4396 7812
rect 8208 7871 8260 7880
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 8392 7871 8444 7880
rect 8392 7837 8401 7871
rect 8401 7837 8435 7871
rect 8435 7837 8444 7871
rect 8392 7828 8444 7837
rect 8484 7828 8536 7880
rect 12072 7905 12081 7939
rect 12081 7905 12115 7939
rect 12115 7905 12124 7939
rect 12072 7896 12124 7905
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 12900 7828 12952 7880
rect 13084 7871 13136 7880
rect 13084 7837 13093 7871
rect 13093 7837 13127 7871
rect 13127 7837 13136 7871
rect 13084 7828 13136 7837
rect 7748 7760 7800 7812
rect 10048 7760 10100 7812
rect 3976 7692 4028 7744
rect 5540 7735 5592 7744
rect 5540 7701 5549 7735
rect 5549 7701 5583 7735
rect 5583 7701 5592 7735
rect 5540 7692 5592 7701
rect 8024 7735 8076 7744
rect 8024 7701 8033 7735
rect 8033 7701 8067 7735
rect 8067 7701 8076 7735
rect 8024 7692 8076 7701
rect 11336 7760 11388 7812
rect 11888 7760 11940 7812
rect 4882 7590 4934 7642
rect 4946 7590 4998 7642
rect 5010 7590 5062 7642
rect 5074 7590 5126 7642
rect 5138 7590 5190 7642
rect 8815 7590 8867 7642
rect 8879 7590 8931 7642
rect 8943 7590 8995 7642
rect 9007 7590 9059 7642
rect 9071 7590 9123 7642
rect 12748 7590 12800 7642
rect 12812 7590 12864 7642
rect 12876 7590 12928 7642
rect 12940 7590 12992 7642
rect 13004 7590 13056 7642
rect 16681 7590 16733 7642
rect 16745 7590 16797 7642
rect 16809 7590 16861 7642
rect 16873 7590 16925 7642
rect 16937 7590 16989 7642
rect 1492 7488 1544 7540
rect 2780 7488 2832 7540
rect 5448 7488 5500 7540
rect 3148 7420 3200 7472
rect 4712 7420 4764 7472
rect 9496 7488 9548 7540
rect 9772 7488 9824 7540
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 2596 7352 2648 7404
rect 4528 7395 4580 7404
rect 2044 7327 2096 7336
rect 2044 7293 2053 7327
rect 2053 7293 2087 7327
rect 2087 7293 2096 7327
rect 4528 7361 4537 7395
rect 4537 7361 4571 7395
rect 4571 7361 4580 7395
rect 4528 7352 4580 7361
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 8576 7420 8628 7472
rect 9680 7420 9732 7472
rect 10048 7463 10100 7472
rect 10048 7429 10057 7463
rect 10057 7429 10091 7463
rect 10091 7429 10100 7463
rect 10048 7420 10100 7429
rect 6000 7352 6052 7404
rect 6552 7395 6604 7404
rect 6552 7361 6561 7395
rect 6561 7361 6595 7395
rect 6595 7361 6604 7395
rect 6552 7352 6604 7361
rect 8484 7352 8536 7404
rect 9864 7352 9916 7404
rect 10324 7395 10376 7404
rect 10324 7361 10333 7395
rect 10333 7361 10367 7395
rect 10367 7361 10376 7395
rect 12348 7420 12400 7472
rect 10324 7352 10376 7361
rect 2044 7284 2096 7293
rect 3608 7284 3660 7336
rect 5632 7216 5684 7268
rect 7564 7284 7616 7336
rect 13268 7395 13320 7404
rect 13268 7361 13277 7395
rect 13277 7361 13311 7395
rect 13311 7361 13320 7395
rect 13268 7352 13320 7361
rect 6736 7259 6788 7268
rect 6736 7225 6745 7259
rect 6745 7225 6779 7259
rect 6779 7225 6788 7259
rect 6736 7216 6788 7225
rect 8208 7216 8260 7268
rect 2320 7148 2372 7200
rect 3884 7191 3936 7200
rect 3884 7157 3893 7191
rect 3893 7157 3927 7191
rect 3927 7157 3936 7191
rect 3884 7148 3936 7157
rect 4160 7148 4212 7200
rect 5356 7148 5408 7200
rect 10232 7148 10284 7200
rect 2916 7046 2968 7098
rect 2980 7046 3032 7098
rect 3044 7046 3096 7098
rect 3108 7046 3160 7098
rect 3172 7046 3224 7098
rect 6849 7046 6901 7098
rect 6913 7046 6965 7098
rect 6977 7046 7029 7098
rect 7041 7046 7093 7098
rect 7105 7046 7157 7098
rect 10782 7046 10834 7098
rect 10846 7046 10898 7098
rect 10910 7046 10962 7098
rect 10974 7046 11026 7098
rect 11038 7046 11090 7098
rect 14715 7046 14767 7098
rect 14779 7046 14831 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 1676 6944 1728 6996
rect 2044 6944 2096 6996
rect 4528 6944 4580 6996
rect 5172 6944 5224 6996
rect 6552 6944 6604 6996
rect 10324 6944 10376 6996
rect 3976 6876 4028 6928
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 2596 6740 2648 6792
rect 3792 6808 3844 6860
rect 5632 6808 5684 6860
rect 2688 6672 2740 6724
rect 3424 6672 3476 6724
rect 4436 6672 4488 6724
rect 5172 6672 5224 6724
rect 5816 6672 5868 6724
rect 8484 6808 8536 6860
rect 9220 6851 9272 6860
rect 9220 6817 9229 6851
rect 9229 6817 9263 6851
rect 9263 6817 9272 6851
rect 9220 6808 9272 6817
rect 6644 6740 6696 6792
rect 7472 6783 7524 6792
rect 7472 6749 7481 6783
rect 7481 6749 7515 6783
rect 7515 6749 7524 6783
rect 7472 6740 7524 6749
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 9312 6783 9364 6792
rect 7564 6740 7616 6749
rect 9312 6749 9321 6783
rect 9321 6749 9355 6783
rect 9355 6749 9364 6783
rect 9312 6740 9364 6749
rect 13084 6740 13136 6792
rect 1860 6604 1912 6656
rect 4344 6604 4396 6656
rect 10140 6647 10192 6656
rect 10140 6613 10149 6647
rect 10149 6613 10183 6647
rect 10183 6613 10192 6647
rect 10140 6604 10192 6613
rect 11152 6672 11204 6724
rect 11244 6604 11296 6656
rect 4882 6502 4934 6554
rect 4946 6502 4998 6554
rect 5010 6502 5062 6554
rect 5074 6502 5126 6554
rect 5138 6502 5190 6554
rect 8815 6502 8867 6554
rect 8879 6502 8931 6554
rect 8943 6502 8995 6554
rect 9007 6502 9059 6554
rect 9071 6502 9123 6554
rect 12748 6502 12800 6554
rect 12812 6502 12864 6554
rect 12876 6502 12928 6554
rect 12940 6502 12992 6554
rect 13004 6502 13056 6554
rect 16681 6502 16733 6554
rect 16745 6502 16797 6554
rect 16809 6502 16861 6554
rect 16873 6502 16925 6554
rect 16937 6502 16989 6554
rect 1676 6443 1728 6452
rect 1676 6409 1685 6443
rect 1685 6409 1719 6443
rect 1719 6409 1728 6443
rect 1676 6400 1728 6409
rect 2320 6443 2372 6452
rect 2320 6409 2329 6443
rect 2329 6409 2363 6443
rect 2363 6409 2372 6443
rect 2320 6400 2372 6409
rect 3332 6400 3384 6452
rect 1860 6307 1912 6316
rect 1860 6273 1869 6307
rect 1869 6273 1903 6307
rect 1903 6273 1912 6307
rect 1860 6264 1912 6273
rect 2412 6264 2464 6316
rect 2688 6307 2740 6316
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 2688 6264 2740 6273
rect 2780 6307 2832 6316
rect 2780 6273 2789 6307
rect 2789 6273 2823 6307
rect 2823 6273 2832 6307
rect 4804 6400 4856 6452
rect 6644 6400 6696 6452
rect 8576 6443 8628 6452
rect 4436 6332 4488 6384
rect 5448 6375 5500 6384
rect 5448 6341 5457 6375
rect 5457 6341 5491 6375
rect 5491 6341 5500 6375
rect 5448 6332 5500 6341
rect 7656 6375 7708 6384
rect 7656 6341 7665 6375
rect 7665 6341 7699 6375
rect 7699 6341 7708 6375
rect 7656 6332 7708 6341
rect 7748 6332 7800 6384
rect 8576 6409 8585 6443
rect 8585 6409 8619 6443
rect 8619 6409 8628 6443
rect 8576 6400 8628 6409
rect 2780 6264 2832 6273
rect 6092 6264 6144 6316
rect 6644 6264 6696 6316
rect 7196 6307 7248 6316
rect 7196 6273 7205 6307
rect 7205 6273 7239 6307
rect 7239 6273 7248 6307
rect 7196 6264 7248 6273
rect 8484 6264 8536 6316
rect 5356 6196 5408 6248
rect 7656 6196 7708 6248
rect 10140 6400 10192 6452
rect 11152 6400 11204 6452
rect 9588 6332 9640 6384
rect 9312 6264 9364 6316
rect 9864 6307 9916 6316
rect 9864 6273 9873 6307
rect 9873 6273 9907 6307
rect 9907 6273 9916 6307
rect 9864 6264 9916 6273
rect 8392 6128 8444 6180
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 10508 6128 10560 6180
rect 4252 6060 4304 6112
rect 8484 6060 8536 6112
rect 9496 6060 9548 6112
rect 2916 5958 2968 6010
rect 2980 5958 3032 6010
rect 3044 5958 3096 6010
rect 3108 5958 3160 6010
rect 3172 5958 3224 6010
rect 6849 5958 6901 6010
rect 6913 5958 6965 6010
rect 6977 5958 7029 6010
rect 7041 5958 7093 6010
rect 7105 5958 7157 6010
rect 10782 5958 10834 6010
rect 10846 5958 10898 6010
rect 10910 5958 10962 6010
rect 10974 5958 11026 6010
rect 11038 5958 11090 6010
rect 14715 5958 14767 6010
rect 14779 5958 14831 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 4712 5856 4764 5908
rect 7196 5856 7248 5908
rect 11244 5899 11296 5908
rect 11244 5865 11253 5899
rect 11253 5865 11287 5899
rect 11287 5865 11296 5899
rect 11244 5856 11296 5865
rect 2320 5788 2372 5840
rect 2504 5788 2556 5840
rect 2688 5788 2740 5840
rect 2596 5720 2648 5772
rect 2228 5652 2280 5704
rect 2964 5720 3016 5772
rect 2780 5652 2832 5704
rect 1860 5516 1912 5568
rect 2688 5559 2740 5568
rect 2688 5525 2697 5559
rect 2697 5525 2731 5559
rect 2731 5525 2740 5559
rect 2688 5516 2740 5525
rect 6644 5788 6696 5840
rect 4436 5763 4488 5772
rect 4436 5729 4445 5763
rect 4445 5729 4479 5763
rect 4479 5729 4488 5763
rect 4436 5720 4488 5729
rect 3608 5652 3660 5704
rect 5540 5720 5592 5772
rect 6736 5720 6788 5772
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 4252 5584 4304 5636
rect 3332 5516 3384 5568
rect 6644 5652 6696 5704
rect 8392 5788 8444 5840
rect 9496 5763 9548 5772
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 9496 5720 9548 5729
rect 9772 5763 9824 5772
rect 9772 5729 9781 5763
rect 9781 5729 9815 5763
rect 9815 5729 9824 5763
rect 9772 5720 9824 5729
rect 5540 5627 5592 5636
rect 5540 5593 5549 5627
rect 5549 5593 5583 5627
rect 5583 5593 5592 5627
rect 5540 5584 5592 5593
rect 9404 5652 9456 5704
rect 10508 5584 10560 5636
rect 5632 5516 5684 5568
rect 7564 5559 7616 5568
rect 7564 5525 7573 5559
rect 7573 5525 7607 5559
rect 7607 5525 7616 5559
rect 7564 5516 7616 5525
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 10140 5516 10192 5568
rect 4882 5414 4934 5466
rect 4946 5414 4998 5466
rect 5010 5414 5062 5466
rect 5074 5414 5126 5466
rect 5138 5414 5190 5466
rect 8815 5414 8867 5466
rect 8879 5414 8931 5466
rect 8943 5414 8995 5466
rect 9007 5414 9059 5466
rect 9071 5414 9123 5466
rect 12748 5414 12800 5466
rect 12812 5414 12864 5466
rect 12876 5414 12928 5466
rect 12940 5414 12992 5466
rect 13004 5414 13056 5466
rect 16681 5414 16733 5466
rect 16745 5414 16797 5466
rect 16809 5414 16861 5466
rect 16873 5414 16925 5466
rect 16937 5414 16989 5466
rect 2228 5312 2280 5364
rect 3240 5312 3292 5364
rect 4620 5312 4672 5364
rect 5632 5355 5684 5364
rect 5632 5321 5641 5355
rect 5641 5321 5675 5355
rect 5675 5321 5684 5355
rect 5632 5312 5684 5321
rect 6644 5355 6696 5364
rect 6644 5321 6653 5355
rect 6653 5321 6687 5355
rect 6687 5321 6696 5355
rect 6644 5312 6696 5321
rect 10324 5312 10376 5364
rect 2136 5244 2188 5296
rect 1768 5219 1820 5228
rect 1768 5185 1777 5219
rect 1777 5185 1811 5219
rect 1811 5185 1820 5219
rect 1768 5176 1820 5185
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2504 5219 2556 5228
rect 2044 5176 2096 5185
rect 2504 5185 2513 5219
rect 2513 5185 2547 5219
rect 2547 5185 2556 5219
rect 2504 5176 2556 5185
rect 2780 5176 2832 5228
rect 4252 5244 4304 5296
rect 4344 5287 4396 5296
rect 4344 5253 4353 5287
rect 4353 5253 4387 5287
rect 4387 5253 4396 5287
rect 4344 5244 4396 5253
rect 4804 5244 4856 5296
rect 5264 5244 5316 5296
rect 2320 5108 2372 5160
rect 4528 5176 4580 5228
rect 5356 5176 5408 5228
rect 8300 5244 8352 5296
rect 9588 5287 9640 5296
rect 9588 5253 9597 5287
rect 9597 5253 9631 5287
rect 9631 5253 9640 5287
rect 9588 5244 9640 5253
rect 6736 5219 6788 5228
rect 6736 5185 6745 5219
rect 6745 5185 6779 5219
rect 6779 5185 6788 5219
rect 6736 5176 6788 5185
rect 10140 5176 10192 5228
rect 4252 5108 4304 5160
rect 8024 5108 8076 5160
rect 1676 4972 1728 5024
rect 2688 4972 2740 5024
rect 3976 5015 4028 5024
rect 3976 4981 3985 5015
rect 3985 4981 4019 5015
rect 4019 4981 4028 5015
rect 3976 4972 4028 4981
rect 2916 4870 2968 4922
rect 2980 4870 3032 4922
rect 3044 4870 3096 4922
rect 3108 4870 3160 4922
rect 3172 4870 3224 4922
rect 6849 4870 6901 4922
rect 6913 4870 6965 4922
rect 6977 4870 7029 4922
rect 7041 4870 7093 4922
rect 7105 4870 7157 4922
rect 10782 4870 10834 4922
rect 10846 4870 10898 4922
rect 10910 4870 10962 4922
rect 10974 4870 11026 4922
rect 11038 4870 11090 4922
rect 14715 4870 14767 4922
rect 14779 4870 14831 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 1584 4768 1636 4820
rect 3700 4768 3752 4820
rect 5540 4811 5592 4820
rect 5540 4777 5549 4811
rect 5549 4777 5583 4811
rect 5583 4777 5592 4811
rect 5540 4768 5592 4777
rect 9772 4768 9824 4820
rect 1492 4700 1544 4752
rect 2596 4743 2648 4752
rect 2596 4709 2605 4743
rect 2605 4709 2639 4743
rect 2639 4709 2648 4743
rect 2596 4700 2648 4709
rect 3792 4700 3844 4752
rect 5448 4700 5500 4752
rect 3056 4632 3108 4684
rect 1860 4607 1912 4616
rect 1860 4573 1869 4607
rect 1869 4573 1903 4607
rect 1903 4573 1912 4607
rect 1860 4564 1912 4573
rect 2320 4496 2372 4548
rect 4068 4564 4120 4616
rect 4160 4607 4212 4616
rect 4160 4573 4169 4607
rect 4169 4573 4203 4607
rect 4203 4573 4212 4607
rect 4160 4564 4212 4573
rect 5264 4564 5316 4616
rect 4712 4496 4764 4548
rect 9312 4564 9364 4616
rect 11244 4564 11296 4616
rect 7748 4539 7800 4548
rect 7748 4505 7757 4539
rect 7757 4505 7791 4539
rect 7791 4505 7800 4539
rect 7748 4496 7800 4505
rect 1860 4428 1912 4480
rect 4882 4326 4934 4378
rect 4946 4326 4998 4378
rect 5010 4326 5062 4378
rect 5074 4326 5126 4378
rect 5138 4326 5190 4378
rect 8815 4326 8867 4378
rect 8879 4326 8931 4378
rect 8943 4326 8995 4378
rect 9007 4326 9059 4378
rect 9071 4326 9123 4378
rect 12748 4326 12800 4378
rect 12812 4326 12864 4378
rect 12876 4326 12928 4378
rect 12940 4326 12992 4378
rect 13004 4326 13056 4378
rect 16681 4326 16733 4378
rect 16745 4326 16797 4378
rect 16809 4326 16861 4378
rect 16873 4326 16925 4378
rect 16937 4326 16989 4378
rect 4068 4267 4120 4276
rect 4068 4233 4077 4267
rect 4077 4233 4111 4267
rect 4111 4233 4120 4267
rect 4068 4224 4120 4233
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 3056 4088 3108 4140
rect 3976 4156 4028 4208
rect 3516 4131 3568 4140
rect 3516 4097 3525 4131
rect 3525 4097 3559 4131
rect 3559 4097 3568 4131
rect 3516 4088 3568 4097
rect 2504 4020 2556 4072
rect 2964 4020 3016 4072
rect 7748 4156 7800 4208
rect 8484 4156 8536 4208
rect 7564 4131 7616 4140
rect 2688 3952 2740 4004
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 1400 3884 1452 3936
rect 1860 3884 1912 3936
rect 3240 3884 3292 3936
rect 2916 3782 2968 3834
rect 2980 3782 3032 3834
rect 3044 3782 3096 3834
rect 3108 3782 3160 3834
rect 3172 3782 3224 3834
rect 6849 3782 6901 3834
rect 6913 3782 6965 3834
rect 6977 3782 7029 3834
rect 7041 3782 7093 3834
rect 7105 3782 7157 3834
rect 10782 3782 10834 3834
rect 10846 3782 10898 3834
rect 10910 3782 10962 3834
rect 10974 3782 11026 3834
rect 11038 3782 11090 3834
rect 14715 3782 14767 3834
rect 14779 3782 14831 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 1952 3680 2004 3732
rect 2780 3723 2832 3732
rect 2780 3689 2789 3723
rect 2789 3689 2823 3723
rect 2823 3689 2832 3723
rect 2780 3680 2832 3689
rect 3792 3680 3844 3732
rect 4068 3680 4120 3732
rect 3332 3655 3384 3664
rect 3332 3621 3341 3655
rect 3341 3621 3375 3655
rect 3375 3621 3384 3655
rect 3332 3612 3384 3621
rect 2044 3519 2096 3528
rect 2044 3485 2053 3519
rect 2053 3485 2087 3519
rect 2087 3485 2096 3519
rect 2044 3476 2096 3485
rect 2412 3476 2464 3528
rect 3608 3408 3660 3460
rect 4344 3476 4396 3528
rect 4882 3238 4934 3290
rect 4946 3238 4998 3290
rect 5010 3238 5062 3290
rect 5074 3238 5126 3290
rect 5138 3238 5190 3290
rect 8815 3238 8867 3290
rect 8879 3238 8931 3290
rect 8943 3238 8995 3290
rect 9007 3238 9059 3290
rect 9071 3238 9123 3290
rect 12748 3238 12800 3290
rect 12812 3238 12864 3290
rect 12876 3238 12928 3290
rect 12940 3238 12992 3290
rect 13004 3238 13056 3290
rect 16681 3238 16733 3290
rect 16745 3238 16797 3290
rect 16809 3238 16861 3290
rect 16873 3238 16925 3290
rect 16937 3238 16989 3290
rect 3424 3179 3476 3188
rect 3424 3145 3433 3179
rect 3433 3145 3467 3179
rect 3467 3145 3476 3179
rect 3424 3136 3476 3145
rect 1768 3068 1820 3120
rect 1860 3043 1912 3052
rect 1860 3009 1869 3043
rect 1869 3009 1903 3043
rect 1903 3009 1912 3043
rect 1860 3000 1912 3009
rect 3608 3000 3660 3052
rect 3976 3043 4028 3052
rect 3976 3009 3985 3043
rect 3985 3009 4019 3043
rect 4019 3009 4028 3043
rect 3976 3000 4028 3009
rect 4252 3000 4304 3052
rect 1400 2796 1452 2848
rect 2916 2694 2968 2746
rect 2980 2694 3032 2746
rect 3044 2694 3096 2746
rect 3108 2694 3160 2746
rect 3172 2694 3224 2746
rect 6849 2694 6901 2746
rect 6913 2694 6965 2746
rect 6977 2694 7029 2746
rect 7041 2694 7093 2746
rect 7105 2694 7157 2746
rect 10782 2694 10834 2746
rect 10846 2694 10898 2746
rect 10910 2694 10962 2746
rect 10974 2694 11026 2746
rect 11038 2694 11090 2746
rect 14715 2694 14767 2746
rect 14779 2694 14831 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 1676 2388 1728 2440
rect 1768 2295 1820 2304
rect 1768 2261 1777 2295
rect 1777 2261 1811 2295
rect 1811 2261 1820 2295
rect 1768 2252 1820 2261
rect 4882 2150 4934 2202
rect 4946 2150 4998 2202
rect 5010 2150 5062 2202
rect 5074 2150 5126 2202
rect 5138 2150 5190 2202
rect 8815 2150 8867 2202
rect 8879 2150 8931 2202
rect 8943 2150 8995 2202
rect 9007 2150 9059 2202
rect 9071 2150 9123 2202
rect 12748 2150 12800 2202
rect 12812 2150 12864 2202
rect 12876 2150 12928 2202
rect 12940 2150 12992 2202
rect 13004 2150 13056 2202
rect 16681 2150 16733 2202
rect 16745 2150 16797 2202
rect 16809 2150 16861 2202
rect 16873 2150 16925 2202
rect 16937 2150 16989 2202
<< metal2 >>
rect 4434 17354 4490 18000
rect 13450 17354 13506 18000
rect 4434 17326 4752 17354
rect 4158 17232 4214 17241
rect 4434 17200 4490 17326
rect 4158 17167 4214 17176
rect 2916 15804 3224 15813
rect 2916 15802 2922 15804
rect 2978 15802 3002 15804
rect 3058 15802 3082 15804
rect 3138 15802 3162 15804
rect 3218 15802 3224 15804
rect 2978 15750 2980 15802
rect 3160 15750 3162 15802
rect 2916 15748 2922 15750
rect 2978 15748 3002 15750
rect 3058 15748 3082 15750
rect 3138 15748 3162 15750
rect 3218 15748 3224 15750
rect 2778 15736 2834 15745
rect 2916 15739 3224 15748
rect 4172 15706 4200 17167
rect 4436 15904 4488 15910
rect 4436 15846 4488 15852
rect 2778 15671 2780 15680
rect 2832 15671 2834 15680
rect 4160 15700 4212 15706
rect 2780 15642 2832 15648
rect 4160 15642 4212 15648
rect 4448 15638 4476 15846
rect 2044 15632 2096 15638
rect 2044 15574 2096 15580
rect 4252 15632 4304 15638
rect 4252 15574 4304 15580
rect 4436 15632 4488 15638
rect 4436 15574 4488 15580
rect 2056 15162 2084 15574
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2412 15428 2464 15434
rect 2412 15370 2464 15376
rect 2424 15162 2452 15370
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 2412 15156 2464 15162
rect 2412 15098 2464 15104
rect 2424 14634 2452 15098
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2332 14618 2452 14634
rect 2320 14612 2452 14618
rect 2372 14606 2452 14612
rect 2320 14554 2372 14560
rect 1674 14240 1730 14249
rect 1674 14175 1730 14184
rect 1688 14074 1716 14175
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1688 12753 1716 13126
rect 2056 12850 2084 13262
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1674 12744 1730 12753
rect 1674 12679 1730 12688
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 11830 1716 12582
rect 2056 12442 2084 12786
rect 2332 12782 2360 13330
rect 2424 12986 2452 14606
rect 2608 13394 2636 14894
rect 2976 14822 3004 15438
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 2916 14716 3224 14725
rect 2916 14714 2922 14716
rect 2978 14714 3002 14716
rect 3058 14714 3082 14716
rect 3138 14714 3162 14716
rect 3218 14714 3224 14716
rect 2978 14662 2980 14714
rect 3160 14662 3162 14714
rect 2916 14660 2922 14662
rect 2978 14660 3002 14662
rect 3058 14660 3082 14662
rect 3138 14660 3162 14662
rect 3218 14660 3224 14662
rect 2916 14651 3224 14660
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2792 13326 2820 14010
rect 2916 13628 3224 13637
rect 2916 13626 2922 13628
rect 2978 13626 3002 13628
rect 3058 13626 3082 13628
rect 3138 13626 3162 13628
rect 3218 13626 3224 13628
rect 2978 13574 2980 13626
rect 3160 13574 3162 13626
rect 2916 13572 2922 13574
rect 2978 13572 3002 13574
rect 3058 13572 3082 13574
rect 3138 13572 3162 13574
rect 3218 13572 3224 13574
rect 2916 13563 3224 13572
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 2412 12980 2464 12986
rect 2412 12922 2464 12928
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 3160 12714 3188 13126
rect 3252 12918 3280 15302
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3620 14346 3648 14758
rect 3608 14340 3660 14346
rect 3608 14282 3660 14288
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3344 14074 3372 14214
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3804 13938 3832 14758
rect 4264 14618 4292 15574
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4724 14346 4752 17326
rect 13450 17326 13768 17354
rect 13450 17200 13506 17326
rect 13740 16574 13768 17326
rect 13740 16546 13860 16574
rect 6849 15804 7157 15813
rect 6849 15802 6855 15804
rect 6911 15802 6935 15804
rect 6991 15802 7015 15804
rect 7071 15802 7095 15804
rect 7151 15802 7157 15804
rect 6911 15750 6913 15802
rect 7093 15750 7095 15802
rect 6849 15748 6855 15750
rect 6911 15748 6935 15750
rect 6991 15748 7015 15750
rect 7071 15748 7095 15750
rect 7151 15748 7157 15750
rect 6849 15739 7157 15748
rect 10782 15804 11090 15813
rect 10782 15802 10788 15804
rect 10844 15802 10868 15804
rect 10924 15802 10948 15804
rect 11004 15802 11028 15804
rect 11084 15802 11090 15804
rect 10844 15750 10846 15802
rect 11026 15750 11028 15802
rect 10782 15748 10788 15750
rect 10844 15748 10868 15750
rect 10924 15748 10948 15750
rect 11004 15748 11028 15750
rect 11084 15748 11090 15750
rect 10782 15739 11090 15748
rect 5908 15632 5960 15638
rect 5908 15574 5960 15580
rect 5920 15502 5948 15574
rect 13832 15570 13860 16546
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 4882 15260 5190 15269
rect 4882 15258 4888 15260
rect 4944 15258 4968 15260
rect 5024 15258 5048 15260
rect 5104 15258 5128 15260
rect 5184 15258 5190 15260
rect 4944 15206 4946 15258
rect 5126 15206 5128 15258
rect 4882 15204 4888 15206
rect 4944 15204 4968 15206
rect 5024 15204 5048 15206
rect 5104 15204 5128 15206
rect 5184 15204 5190 15206
rect 4882 15195 5190 15204
rect 4712 14340 4764 14346
rect 4712 14282 4764 14288
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 4882 14172 5190 14181
rect 4882 14170 4888 14172
rect 4944 14170 4968 14172
rect 5024 14170 5048 14172
rect 5104 14170 5128 14172
rect 5184 14170 5190 14172
rect 4944 14118 4946 14170
rect 5126 14118 5128 14170
rect 4882 14116 4888 14118
rect 4944 14116 4968 14118
rect 5024 14116 5048 14118
rect 5104 14116 5128 14118
rect 5184 14116 5190 14118
rect 4882 14107 5190 14116
rect 5460 14074 5488 14282
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 4068 14000 4120 14006
rect 4066 13968 4068 13977
rect 4120 13968 4122 13977
rect 3792 13932 3844 13938
rect 5368 13954 5396 14010
rect 5552 13954 5580 15438
rect 6368 15428 6420 15434
rect 6368 15370 6420 15376
rect 6552 15428 6604 15434
rect 6552 15370 6604 15376
rect 6380 15026 6408 15370
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5368 13926 5580 13954
rect 4066 13903 4122 13912
rect 3792 13874 3844 13880
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4632 13462 4660 13670
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4620 13456 4672 13462
rect 4620 13398 4672 13404
rect 4816 13326 4844 13466
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 3240 12912 3292 12918
rect 3240 12854 3292 12860
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 2916 12540 3224 12549
rect 2916 12538 2922 12540
rect 2978 12538 3002 12540
rect 3058 12538 3082 12540
rect 3138 12538 3162 12540
rect 3218 12538 3224 12540
rect 2978 12486 2980 12538
rect 3160 12486 3162 12538
rect 2916 12484 2922 12486
rect 2978 12484 3002 12486
rect 3058 12484 3082 12486
rect 3138 12484 3162 12486
rect 3218 12484 3224 12486
rect 2916 12475 3224 12484
rect 2044 12436 2096 12442
rect 3252 12434 3280 12854
rect 2044 12378 2096 12384
rect 3160 12406 3280 12434
rect 1676 11824 1728 11830
rect 1676 11766 1728 11772
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 1676 11280 1728 11286
rect 1674 11248 1676 11257
rect 1728 11248 1730 11257
rect 1674 11183 1730 11192
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1504 7546 1532 8434
rect 1492 7540 1544 7546
rect 1492 7482 1544 7488
rect 1490 5264 1546 5273
rect 1490 5199 1546 5208
rect 1504 4758 1532 5199
rect 1596 4826 1624 9998
rect 1952 9988 2004 9994
rect 1952 9930 2004 9936
rect 1766 9752 1822 9761
rect 1766 9687 1822 9696
rect 1780 8634 1808 9687
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1766 8256 1822 8265
rect 1766 8191 1822 8200
rect 1780 8090 1808 8191
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1688 7002 1716 7822
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1780 6798 1808 7346
rect 1768 6792 1820 6798
rect 1674 6760 1730 6769
rect 1768 6734 1820 6740
rect 1674 6695 1730 6704
rect 1688 6458 1716 6695
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1780 5234 1808 6734
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1872 6322 1900 6598
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1492 4752 1544 4758
rect 1492 4694 1544 4700
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 1412 3777 1440 3878
rect 1398 3768 1454 3777
rect 1398 3703 1454 3712
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1412 785 1440 2790
rect 1688 2446 1716 4966
rect 1780 3126 1808 5170
rect 1872 4622 1900 5510
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1872 4146 1900 4422
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1768 3120 1820 3126
rect 1768 3062 1820 3068
rect 1872 3058 1900 3878
rect 1964 3738 1992 9930
rect 2044 7336 2096 7342
rect 2044 7278 2096 7284
rect 2056 7002 2084 7278
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 2056 5234 2084 6734
rect 2148 5302 2176 11494
rect 2700 11354 2728 11630
rect 3160 11558 3188 12406
rect 3240 12164 3292 12170
rect 3240 12106 3292 12112
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 2916 11452 3224 11461
rect 2916 11450 2922 11452
rect 2978 11450 3002 11452
rect 3058 11450 3082 11452
rect 3138 11450 3162 11452
rect 3218 11450 3224 11452
rect 2978 11398 2980 11450
rect 3160 11398 3162 11450
rect 2916 11396 2922 11398
rect 2978 11396 3002 11398
rect 3058 11396 3082 11398
rect 3138 11396 3162 11398
rect 3218 11396 3224 11398
rect 2916 11387 3224 11396
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2916 10364 3224 10373
rect 2916 10362 2922 10364
rect 2978 10362 3002 10364
rect 3058 10362 3082 10364
rect 3138 10362 3162 10364
rect 3218 10362 3224 10364
rect 2978 10310 2980 10362
rect 3160 10310 3162 10362
rect 2916 10308 2922 10310
rect 2978 10308 3002 10310
rect 3058 10308 3082 10310
rect 3138 10308 3162 10310
rect 3218 10308 3224 10310
rect 2916 10299 3224 10308
rect 2916 9276 3224 9285
rect 2916 9274 2922 9276
rect 2978 9274 3002 9276
rect 3058 9274 3082 9276
rect 3138 9274 3162 9276
rect 3218 9274 3224 9276
rect 2978 9222 2980 9274
rect 3160 9222 3162 9274
rect 2916 9220 2922 9222
rect 2978 9220 3002 9222
rect 3058 9220 3082 9222
rect 3138 9220 3162 9222
rect 3218 9220 3224 9222
rect 2916 9211 3224 9220
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2608 8498 2636 8774
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2916 8188 3224 8197
rect 2916 8186 2922 8188
rect 2978 8186 3002 8188
rect 3058 8186 3082 8188
rect 3138 8186 3162 8188
rect 3218 8186 3224 8188
rect 2978 8134 2980 8186
rect 3160 8134 3162 8186
rect 2916 8132 2922 8134
rect 2978 8132 3002 8134
rect 3058 8132 3082 8134
rect 3138 8132 3162 8134
rect 3218 8132 3224 8134
rect 2916 8123 3224 8132
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2332 6458 2360 7142
rect 2608 6798 2636 7346
rect 2792 7018 2820 7482
rect 3160 7478 3188 7822
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 2916 7100 3224 7109
rect 2916 7098 2922 7100
rect 2978 7098 3002 7100
rect 3058 7098 3082 7100
rect 3138 7098 3162 7100
rect 3218 7098 3224 7100
rect 2978 7046 2980 7098
rect 3160 7046 3162 7098
rect 2916 7044 2922 7046
rect 2978 7044 3002 7046
rect 3058 7044 3082 7046
rect 3138 7044 3162 7046
rect 3218 7044 3224 7046
rect 2916 7035 3224 7044
rect 2700 6990 2820 7018
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2332 5846 2360 6394
rect 2412 6316 2464 6322
rect 2608 6304 2636 6734
rect 2700 6730 2728 6990
rect 2688 6724 2740 6730
rect 2688 6666 2740 6672
rect 2700 6474 2728 6666
rect 2700 6446 2820 6474
rect 2792 6322 2820 6446
rect 2688 6316 2740 6322
rect 2608 6276 2688 6304
rect 2412 6258 2464 6264
rect 2688 6258 2740 6264
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2320 5840 2372 5846
rect 2320 5782 2372 5788
rect 2228 5704 2280 5710
rect 2424 5658 2452 6258
rect 2700 5846 2728 6258
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2228 5646 2280 5652
rect 2240 5370 2268 5646
rect 2332 5630 2452 5658
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2136 5296 2188 5302
rect 2136 5238 2188 5244
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 2332 5166 2360 5630
rect 2516 5386 2544 5782
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2424 5358 2544 5386
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 2332 4554 2360 5102
rect 2320 4548 2372 4554
rect 2320 4490 2372 4496
rect 2042 4040 2098 4049
rect 2042 3975 2098 3984
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 2056 3534 2084 3975
rect 2424 3534 2452 5358
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2516 4078 2544 5170
rect 2608 4758 2636 5714
rect 2792 5710 2820 6258
rect 2916 6012 3224 6021
rect 2916 6010 2922 6012
rect 2978 6010 3002 6012
rect 3058 6010 3082 6012
rect 3138 6010 3162 6012
rect 3218 6010 3224 6012
rect 2978 5958 2980 6010
rect 3160 5958 3162 6010
rect 2916 5956 2922 5958
rect 2978 5956 3002 5958
rect 3058 5956 3082 5958
rect 3138 5956 3162 5958
rect 3218 5956 3224 5958
rect 2916 5947 3224 5956
rect 2964 5772 3016 5778
rect 3016 5732 3188 5760
rect 2964 5714 3016 5720
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2700 5030 2728 5510
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 2596 4752 2648 4758
rect 2596 4694 2648 4700
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2700 4010 2728 4966
rect 2792 4060 2820 5170
rect 3160 5114 3188 5732
rect 3252 5370 3280 12106
rect 3344 11218 3372 13262
rect 4816 12850 4844 13262
rect 5644 13258 5672 14758
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 5724 13388 5776 13394
rect 5828 13376 5856 14418
rect 6472 14346 6500 14894
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 6564 14278 6592 15370
rect 7840 15360 7892 15366
rect 7840 15302 7892 15308
rect 6736 15088 6788 15094
rect 6736 15030 6788 15036
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 6104 13734 6132 13874
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 5776 13348 5856 13376
rect 5724 13330 5776 13336
rect 5632 13252 5684 13258
rect 5632 13194 5684 13200
rect 4882 13084 5190 13093
rect 4882 13082 4888 13084
rect 4944 13082 4968 13084
rect 5024 13082 5048 13084
rect 5104 13082 5128 13084
rect 5184 13082 5190 13084
rect 4944 13030 4946 13082
rect 5126 13030 5128 13082
rect 4882 13028 4888 13030
rect 4944 13028 4968 13030
rect 5024 13028 5048 13030
rect 5104 13028 5128 13030
rect 5184 13028 5190 13030
rect 4882 13019 5190 13028
rect 5828 12918 5856 13348
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 4080 11694 4108 12786
rect 5092 12730 5120 12786
rect 4540 12714 5120 12730
rect 4528 12708 5120 12714
rect 4580 12702 5120 12708
rect 4528 12650 4580 12656
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 4068 11076 4120 11082
rect 4120 11036 4200 11064
rect 4068 11018 4120 11024
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4080 10198 4108 10746
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 3332 9988 3384 9994
rect 3332 9930 3384 9936
rect 3344 9654 3372 9930
rect 3976 9920 4028 9926
rect 3976 9862 4028 9868
rect 3988 9761 4016 9862
rect 3974 9752 4030 9761
rect 3974 9687 4030 9696
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 3344 6458 3372 9590
rect 3516 8968 3568 8974
rect 4080 8922 4108 10134
rect 4172 9518 4200 11036
rect 4264 10742 4292 12106
rect 4882 11996 5190 12005
rect 4882 11994 4888 11996
rect 4944 11994 4968 11996
rect 5024 11994 5048 11996
rect 5104 11994 5128 11996
rect 5184 11994 5190 11996
rect 4944 11942 4946 11994
rect 5126 11942 5128 11994
rect 4882 11940 4888 11942
rect 4944 11940 4968 11942
rect 5024 11940 5048 11942
rect 5104 11940 5128 11942
rect 5184 11940 5190 11942
rect 4882 11931 5190 11940
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 4436 11824 4488 11830
rect 4436 11766 4488 11772
rect 4448 11286 4476 11766
rect 5276 11558 5304 11834
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4252 9104 4304 9110
rect 4252 9046 4304 9052
rect 3516 8910 3568 8916
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3160 5086 3280 5114
rect 2916 4924 3224 4933
rect 2916 4922 2922 4924
rect 2978 4922 3002 4924
rect 3058 4922 3082 4924
rect 3138 4922 3162 4924
rect 3218 4922 3224 4924
rect 2978 4870 2980 4922
rect 3160 4870 3162 4922
rect 2916 4868 2922 4870
rect 2978 4868 3002 4870
rect 3058 4868 3082 4870
rect 3138 4868 3162 4870
rect 3218 4868 3224 4870
rect 2916 4859 3224 4868
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 3068 4146 3096 4626
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 2964 4072 3016 4078
rect 2792 4032 2964 4060
rect 2688 4004 2740 4010
rect 2688 3946 2740 3952
rect 2792 3738 2820 4032
rect 2964 4014 3016 4020
rect 3252 3942 3280 5086
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 2916 3836 3224 3845
rect 2916 3834 2922 3836
rect 2978 3834 3002 3836
rect 3058 3834 3082 3836
rect 3138 3834 3162 3836
rect 3218 3834 3224 3836
rect 2978 3782 2980 3834
rect 3160 3782 3162 3834
rect 2916 3780 2922 3782
rect 2978 3780 3002 3782
rect 3058 3780 3082 3782
rect 3138 3780 3162 3782
rect 3218 3780 3224 3782
rect 2916 3771 3224 3780
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 3344 3670 3372 5510
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 3436 3194 3464 6666
rect 3528 4146 3556 8910
rect 3700 8900 3752 8906
rect 3700 8842 3752 8848
rect 3896 8894 4108 8922
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3620 5710 3648 7278
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3620 3466 3648 5646
rect 3712 4826 3740 8842
rect 3792 8016 3844 8022
rect 3792 7958 3844 7964
rect 3896 7970 3924 8894
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4172 8022 4200 8434
rect 4160 8016 4212 8022
rect 3804 6866 3832 7958
rect 3896 7942 4108 7970
rect 4160 7958 4212 7964
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3896 7206 3924 7822
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3988 6934 4016 7686
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 3804 3738 3832 4694
rect 3988 4214 4016 4966
rect 4080 4622 4108 7942
rect 4264 7886 4292 9046
rect 4356 8974 4384 11086
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4540 9926 4568 10950
rect 4632 10266 4660 11018
rect 4882 10908 5190 10917
rect 4882 10906 4888 10908
rect 4944 10906 4968 10908
rect 5024 10906 5048 10908
rect 5104 10906 5128 10908
rect 5184 10906 5190 10908
rect 4944 10854 4946 10906
rect 5126 10854 5128 10906
rect 4882 10852 4888 10854
rect 4944 10852 4968 10854
rect 5024 10852 5048 10854
rect 5104 10852 5128 10854
rect 5184 10852 5190 10854
rect 4882 10843 5190 10852
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 5276 10062 5304 11494
rect 5644 11354 5672 12582
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5920 11898 5948 12174
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5920 10266 5948 11698
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 4448 9042 4476 9590
rect 4540 9382 4568 9862
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4356 7818 4384 8910
rect 4540 8838 4568 9318
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4632 8430 4660 9930
rect 4882 9820 5190 9829
rect 4882 9818 4888 9820
rect 4944 9818 4968 9820
rect 5024 9818 5048 9820
rect 5104 9818 5128 9820
rect 5184 9818 5190 9820
rect 4944 9766 4946 9818
rect 5126 9766 5128 9818
rect 4882 9764 4888 9766
rect 4944 9764 4968 9766
rect 5024 9764 5048 9766
rect 5104 9764 5128 9766
rect 5184 9764 5190 9766
rect 4882 9755 5190 9764
rect 5368 9586 5396 10202
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4172 4622 4200 7142
rect 4448 6730 4476 8298
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4540 7002 4568 7346
rect 4528 6996 4580 7002
rect 4528 6938 4580 6944
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4264 5642 4292 6054
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 4264 5302 4292 5578
rect 4356 5302 4384 6598
rect 4448 6474 4476 6666
rect 4448 6446 4568 6474
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4448 5778 4476 6326
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4252 5296 4304 5302
rect 4252 5238 4304 5244
rect 4344 5296 4396 5302
rect 4344 5238 4396 5244
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4080 4282 4108 4558
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3608 3460 3660 3466
rect 3608 3402 3660 3408
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3620 3058 3648 3402
rect 3988 3058 4016 4150
rect 4080 3738 4108 4218
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4264 3058 4292 5102
rect 4356 3534 4384 5238
rect 4540 5234 4568 6446
rect 4632 5370 4660 8366
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4724 5914 4752 7414
rect 4816 6458 4844 9318
rect 5092 8974 5120 9454
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 4882 8732 5190 8741
rect 4882 8730 4888 8732
rect 4944 8730 4968 8732
rect 5024 8730 5048 8732
rect 5104 8730 5128 8732
rect 5184 8730 5190 8732
rect 4944 8678 4946 8730
rect 5126 8678 5128 8730
rect 4882 8676 4888 8678
rect 4944 8676 4968 8678
rect 5024 8676 5048 8678
rect 5104 8676 5128 8678
rect 5184 8676 5190 8678
rect 4882 8667 5190 8676
rect 5276 8362 5304 9318
rect 5368 9110 5396 9522
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5368 8242 5396 8434
rect 5276 8214 5396 8242
rect 4882 7644 5190 7653
rect 4882 7642 4888 7644
rect 4944 7642 4968 7644
rect 5024 7642 5048 7644
rect 5104 7642 5128 7644
rect 5184 7642 5190 7644
rect 4944 7590 4946 7642
rect 5126 7590 5128 7642
rect 4882 7588 4888 7590
rect 4944 7588 4968 7590
rect 5024 7588 5048 7590
rect 5104 7588 5128 7590
rect 5184 7588 5190 7590
rect 4882 7579 5190 7588
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5184 7313 5212 7346
rect 5170 7304 5226 7313
rect 5170 7239 5226 7248
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5184 6730 5212 6938
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 4882 6556 5190 6565
rect 4882 6554 4888 6556
rect 4944 6554 4968 6556
rect 5024 6554 5048 6556
rect 5104 6554 5128 6556
rect 5184 6554 5190 6556
rect 4944 6502 4946 6554
rect 5126 6502 5128 6554
rect 4882 6500 4888 6502
rect 4944 6500 4968 6502
rect 5024 6500 5048 6502
rect 5104 6500 5128 6502
rect 5184 6500 5190 6502
rect 4882 6491 5190 6500
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4724 4554 4752 5850
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4816 5302 4844 5646
rect 4882 5468 5190 5477
rect 4882 5466 4888 5468
rect 4944 5466 4968 5468
rect 5024 5466 5048 5468
rect 5104 5466 5128 5468
rect 5184 5466 5190 5468
rect 4944 5414 4946 5466
rect 5126 5414 5128 5466
rect 4882 5412 4888 5414
rect 4944 5412 4968 5414
rect 5024 5412 5048 5414
rect 5104 5412 5128 5414
rect 5184 5412 5190 5414
rect 4882 5403 5190 5412
rect 5276 5302 5304 8214
rect 5460 7886 5488 8774
rect 5736 8022 5764 10202
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5828 8498 5856 9522
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5920 8906 5948 9386
rect 6288 9042 6316 11154
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6380 9654 6408 11018
rect 6564 10742 6592 14214
rect 6748 14074 6776 15030
rect 6849 14716 7157 14725
rect 6849 14714 6855 14716
rect 6911 14714 6935 14716
rect 6991 14714 7015 14716
rect 7071 14714 7095 14716
rect 7151 14714 7157 14716
rect 6911 14662 6913 14714
rect 7093 14662 7095 14714
rect 6849 14660 6855 14662
rect 6911 14660 6935 14662
rect 6991 14660 7015 14662
rect 7071 14660 7095 14662
rect 7151 14660 7157 14662
rect 6849 14651 7157 14660
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 7392 13938 7420 14214
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7852 13870 7880 15302
rect 8312 14958 8340 15438
rect 8668 15428 8720 15434
rect 8668 15370 8720 15376
rect 8680 15094 8708 15370
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 8815 15260 9123 15269
rect 8815 15258 8821 15260
rect 8877 15258 8901 15260
rect 8957 15258 8981 15260
rect 9037 15258 9061 15260
rect 9117 15258 9123 15260
rect 8877 15206 8879 15258
rect 9059 15206 9061 15258
rect 8815 15204 8821 15206
rect 8877 15204 8901 15206
rect 8957 15204 8981 15206
rect 9037 15204 9061 15206
rect 9117 15204 9123 15206
rect 8815 15195 9123 15204
rect 9324 15094 9352 15302
rect 8668 15088 8720 15094
rect 8668 15030 8720 15036
rect 9312 15088 9364 15094
rect 9312 15030 9364 15036
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 8128 14618 8156 14894
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8312 14414 8340 14894
rect 9600 14618 9628 14894
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9784 14414 9812 14894
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10152 14550 10180 14758
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 10244 14414 10272 15302
rect 10336 14958 10364 15438
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10980 15094 11008 15302
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10428 14278 10456 14962
rect 10968 14816 11020 14822
rect 11072 14804 11100 15302
rect 11348 15026 11376 15438
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 11020 14776 11100 14804
rect 11152 14816 11204 14822
rect 10968 14758 11020 14764
rect 11152 14758 11204 14764
rect 10782 14716 11090 14725
rect 10782 14714 10788 14716
rect 10844 14714 10868 14716
rect 10924 14714 10948 14716
rect 11004 14714 11028 14716
rect 11084 14714 11090 14716
rect 10844 14662 10846 14714
rect 11026 14662 11028 14714
rect 10782 14660 10788 14662
rect 10844 14660 10868 14662
rect 10924 14660 10948 14662
rect 11004 14660 11028 14662
rect 11084 14660 11090 14662
rect 10782 14651 11090 14660
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 8815 14172 9123 14181
rect 8815 14170 8821 14172
rect 8877 14170 8901 14172
rect 8957 14170 8981 14172
rect 9037 14170 9061 14172
rect 9117 14170 9123 14172
rect 8877 14118 8879 14170
rect 9059 14118 9061 14170
rect 8815 14116 8821 14118
rect 8877 14116 8901 14118
rect 8957 14116 8981 14118
rect 9037 14116 9061 14118
rect 9117 14116 9123 14118
rect 8815 14107 9123 14116
rect 10888 14113 10916 14214
rect 10874 14104 10930 14113
rect 10874 14039 10930 14048
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9772 13932 9824 13938
rect 10612 13926 11008 13954
rect 10612 13920 10640 13926
rect 9772 13874 9824 13880
rect 10428 13892 10640 13920
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 7748 13728 7800 13734
rect 7748 13670 7800 13676
rect 6748 13326 6776 13670
rect 6849 13628 7157 13637
rect 6849 13626 6855 13628
rect 6911 13626 6935 13628
rect 6991 13626 7015 13628
rect 7071 13626 7095 13628
rect 7151 13626 7157 13628
rect 6911 13574 6913 13626
rect 7093 13574 7095 13626
rect 6849 13572 6855 13574
rect 6911 13572 6935 13574
rect 6991 13572 7015 13574
rect 7071 13572 7095 13574
rect 7151 13572 7157 13574
rect 6849 13563 7157 13572
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6748 12850 6776 13126
rect 7116 12918 7144 13194
rect 7760 13190 7788 13670
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7852 13190 7880 13330
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 6849 12540 7157 12549
rect 6849 12538 6855 12540
rect 6911 12538 6935 12540
rect 6991 12538 7015 12540
rect 7071 12538 7095 12540
rect 7151 12538 7157 12540
rect 6911 12486 6913 12538
rect 7093 12486 7095 12538
rect 6849 12484 6855 12486
rect 6911 12484 6935 12486
rect 6991 12484 7015 12486
rect 7071 12484 7095 12486
rect 7151 12484 7157 12486
rect 6849 12475 7157 12484
rect 7208 12102 7236 12582
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7300 11898 7328 12106
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6748 11286 6776 11562
rect 6849 11452 7157 11461
rect 6849 11450 6855 11452
rect 6911 11450 6935 11452
rect 6991 11450 7015 11452
rect 7071 11450 7095 11452
rect 7151 11450 7157 11452
rect 6911 11398 6913 11450
rect 7093 11398 7095 11450
rect 6849 11396 6855 11398
rect 6911 11396 6935 11398
rect 6991 11396 7015 11398
rect 7071 11396 7095 11398
rect 7151 11396 7157 11398
rect 6849 11387 7157 11396
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 7288 11280 7340 11286
rect 7288 11222 7340 11228
rect 6552 10736 6604 10742
rect 6552 10678 6604 10684
rect 6849 10364 7157 10373
rect 6849 10362 6855 10364
rect 6911 10362 6935 10364
rect 6991 10362 7015 10364
rect 7071 10362 7095 10364
rect 7151 10362 7157 10364
rect 6911 10310 6913 10362
rect 7093 10310 7095 10362
rect 6849 10308 6855 10310
rect 6911 10308 6935 10310
rect 6991 10308 7015 10310
rect 7071 10308 7095 10310
rect 7151 10308 7157 10310
rect 6849 10299 7157 10308
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6656 9042 6684 9318
rect 6849 9276 7157 9285
rect 6849 9274 6855 9276
rect 6911 9274 6935 9276
rect 6991 9274 7015 9276
rect 7071 9274 7095 9276
rect 7151 9274 7157 9276
rect 6911 9222 6913 9274
rect 7093 9222 7095 9274
rect 6849 9220 6855 9222
rect 6911 9220 6935 9222
rect 6991 9220 7015 9222
rect 7071 9220 7095 9222
rect 7151 9220 7157 9222
rect 6849 9211 7157 9220
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5724 8016 5776 8022
rect 5724 7958 5776 7964
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5368 6254 5396 7142
rect 5460 6390 5488 7482
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 5264 5296 5316 5302
rect 5264 5238 5316 5244
rect 5368 5234 5396 6190
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5264 4616 5316 4622
rect 5368 4604 5396 5170
rect 5460 4758 5488 6326
rect 5552 5778 5580 7686
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 5644 6866 5672 7210
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5828 6730 5856 8298
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 6012 7410 6040 8230
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 6104 6322 6132 8774
rect 7300 8430 7328 11222
rect 7668 11150 7696 11698
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7576 9178 7604 10066
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7484 8362 7512 8910
rect 7576 8566 7604 9114
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 6849 8188 7157 8197
rect 6849 8186 6855 8188
rect 6911 8186 6935 8188
rect 6991 8186 7015 8188
rect 7071 8186 7095 8188
rect 7151 8186 7157 8188
rect 6911 8134 6913 8186
rect 7093 8134 7095 8186
rect 6849 8132 6855 8134
rect 6911 8132 6935 8134
rect 6991 8132 7015 8134
rect 7071 8132 7095 8134
rect 7151 8132 7157 8134
rect 6849 8123 7157 8132
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6564 7002 6592 7346
rect 6734 7304 6790 7313
rect 6734 7239 6736 7248
rect 6788 7239 6790 7248
rect 6736 7210 6788 7216
rect 6849 7100 7157 7109
rect 6849 7098 6855 7100
rect 6911 7098 6935 7100
rect 6991 7098 7015 7100
rect 7071 7098 7095 7100
rect 7151 7098 7157 7100
rect 6911 7046 6913 7098
rect 7093 7046 7095 7098
rect 6849 7044 6855 7046
rect 6911 7044 6935 7046
rect 6991 7044 7015 7046
rect 7071 7044 7095 7046
rect 7151 7044 7157 7046
rect 6849 7035 7157 7044
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 7484 6798 7512 8298
rect 7576 7342 7604 8502
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7576 6798 7604 7278
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 6656 6458 6684 6734
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 6656 5846 6684 6258
rect 6849 6012 7157 6021
rect 6849 6010 6855 6012
rect 6911 6010 6935 6012
rect 6991 6010 7015 6012
rect 7071 6010 7095 6012
rect 7151 6010 7157 6012
rect 6911 5958 6913 6010
rect 7093 5958 7095 6010
rect 6849 5956 6855 5958
rect 6911 5956 6935 5958
rect 6991 5956 7015 5958
rect 7071 5956 7095 5958
rect 7151 5956 7157 5958
rect 6849 5947 7157 5956
rect 7208 5914 7236 6258
rect 7576 6202 7604 6734
rect 7668 6390 7696 11086
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7760 10130 7788 10950
rect 7852 10810 7880 13126
rect 8496 12850 8524 13126
rect 8815 13084 9123 13093
rect 8815 13082 8821 13084
rect 8877 13082 8901 13084
rect 8957 13082 8981 13084
rect 9037 13082 9061 13084
rect 9117 13082 9123 13084
rect 8877 13030 8879 13082
rect 9059 13030 9061 13082
rect 8815 13028 8821 13030
rect 8877 13028 8901 13030
rect 8957 13028 8981 13030
rect 9037 13028 9061 13030
rect 9117 13028 9123 13030
rect 8815 13019 9123 13028
rect 9324 12918 9352 13126
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8036 12102 8064 12786
rect 9692 12102 9720 13874
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 8036 11762 8064 12038
rect 8815 11996 9123 12005
rect 8815 11994 8821 11996
rect 8877 11994 8901 11996
rect 8957 11994 8981 11996
rect 9037 11994 9061 11996
rect 9117 11994 9123 11996
rect 8877 11942 8879 11994
rect 9059 11942 9061 11994
rect 8815 11940 8821 11942
rect 8877 11940 8901 11942
rect 8957 11940 8981 11942
rect 9037 11940 9061 11942
rect 9117 11940 9123 11942
rect 8815 11931 9123 11940
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7944 9518 7972 11018
rect 8128 9586 8156 11834
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 8312 10470 8340 11562
rect 9232 11354 9260 11698
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 8815 10908 9123 10917
rect 8815 10906 8821 10908
rect 8877 10906 8901 10908
rect 8957 10906 8981 10908
rect 9037 10906 9061 10908
rect 9117 10906 9123 10908
rect 8877 10854 8879 10906
rect 9059 10854 9061 10906
rect 8815 10852 8821 10854
rect 8877 10852 8901 10854
rect 8957 10852 8981 10854
rect 9037 10852 9061 10854
rect 9117 10852 9123 10854
rect 8815 10843 9123 10852
rect 9324 10606 9352 11086
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8312 9654 8340 10406
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7944 8634 7972 9454
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8312 7954 8340 8230
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 7748 7812 7800 7818
rect 7748 7754 7800 7760
rect 7760 6390 7788 7754
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7656 6248 7708 6254
rect 7576 6196 7656 6202
rect 7576 6190 7708 6196
rect 7576 6174 7696 6190
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 6644 5840 6696 5846
rect 6644 5782 6696 5788
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5552 4826 5580 5578
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5644 5370 5672 5510
rect 6656 5370 6684 5646
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6748 5234 6776 5714
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6849 4924 7157 4933
rect 6849 4922 6855 4924
rect 6911 4922 6935 4924
rect 6991 4922 7015 4924
rect 7071 4922 7095 4924
rect 7151 4922 7157 4924
rect 6911 4870 6913 4922
rect 7093 4870 7095 4922
rect 6849 4868 6855 4870
rect 6911 4868 6935 4870
rect 6991 4868 7015 4870
rect 7071 4868 7095 4870
rect 7151 4868 7157 4870
rect 6849 4859 7157 4868
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 5316 4576 5396 4604
rect 5264 4558 5316 4564
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4882 4380 5190 4389
rect 4882 4378 4888 4380
rect 4944 4378 4968 4380
rect 5024 4378 5048 4380
rect 5104 4378 5128 4380
rect 5184 4378 5190 4380
rect 4944 4326 4946 4378
rect 5126 4326 5128 4378
rect 4882 4324 4888 4326
rect 4944 4324 4968 4326
rect 5024 4324 5048 4326
rect 5104 4324 5128 4326
rect 5184 4324 5190 4326
rect 4882 4315 5190 4324
rect 7576 4146 7604 5510
rect 8036 5166 8064 7686
rect 8220 7274 8248 7822
rect 8208 7268 8260 7274
rect 8208 7210 8260 7216
rect 8312 5302 8340 7890
rect 8404 7886 8432 9862
rect 8815 9820 9123 9829
rect 8815 9818 8821 9820
rect 8877 9818 8901 9820
rect 8957 9818 8981 9820
rect 9037 9818 9061 9820
rect 9117 9818 9123 9820
rect 8877 9766 8879 9818
rect 9059 9766 9061 9818
rect 8815 9764 8821 9766
rect 8877 9764 8901 9766
rect 8957 9764 8981 9766
rect 9037 9764 9061 9766
rect 9117 9764 9123 9766
rect 8815 9755 9123 9764
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 8815 8732 9123 8741
rect 8815 8730 8821 8732
rect 8877 8730 8901 8732
rect 8957 8730 8981 8732
rect 9037 8730 9061 8732
rect 9117 8730 9123 8732
rect 8877 8678 8879 8730
rect 9059 8678 9061 8730
rect 8815 8676 8821 8678
rect 8877 8676 8901 8678
rect 8957 8676 8981 8678
rect 9037 8676 9061 8678
rect 9117 8676 9123 8678
rect 8815 8667 9123 8676
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8496 7886 8524 8230
rect 9128 8016 9180 8022
rect 9128 7958 9180 7964
rect 9140 7886 9168 7958
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 8496 7410 8524 7822
rect 8815 7644 9123 7653
rect 8815 7642 8821 7644
rect 8877 7642 8901 7644
rect 8957 7642 8981 7644
rect 9037 7642 9061 7644
rect 9117 7642 9123 7644
rect 8877 7590 8879 7642
rect 9059 7590 9061 7642
rect 8815 7588 8821 7590
rect 8877 7588 8901 7590
rect 8957 7588 8981 7590
rect 9037 7588 9061 7590
rect 9117 7588 9123 7590
rect 8815 7579 9123 7588
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8496 6866 8524 7346
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8496 6322 8524 6802
rect 8588 6458 8616 7414
rect 9232 6866 9260 8910
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9324 6798 9352 10542
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9416 10062 9444 10406
rect 9508 10130 9536 11630
rect 9600 11558 9628 11698
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9600 11150 9628 11494
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9416 9654 9444 9862
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9508 8566 9536 10066
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9508 7546 9536 8502
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 8815 6556 9123 6565
rect 8815 6554 8821 6556
rect 8877 6554 8901 6556
rect 8957 6554 8981 6556
rect 9037 6554 9061 6556
rect 9117 6554 9123 6556
rect 8877 6502 8879 6554
rect 9059 6502 9061 6554
rect 8815 6500 8821 6502
rect 8877 6500 8901 6502
rect 8957 6500 8981 6502
rect 9037 6500 9061 6502
rect 9117 6500 9123 6502
rect 8815 6491 9123 6500
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 9600 6390 9628 9454
rect 9692 7478 9720 12038
rect 9784 11218 9812 13874
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10232 12164 10284 12170
rect 10232 12106 10284 12112
rect 10244 11354 10272 12106
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 10336 10810 10364 13806
rect 10428 13734 10456 13892
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10980 13818 11008 13926
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10600 13524 10652 13530
rect 10600 13466 10652 13472
rect 10612 12782 10640 13466
rect 10704 12918 10732 13806
rect 10980 13790 11100 13818
rect 11072 13734 11100 13790
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 10782 13628 11090 13637
rect 10782 13626 10788 13628
rect 10844 13626 10868 13628
rect 10924 13626 10948 13628
rect 11004 13626 11028 13628
rect 11084 13626 11090 13628
rect 10844 13574 10846 13626
rect 11026 13574 11028 13626
rect 10782 13572 10788 13574
rect 10844 13572 10868 13574
rect 10924 13572 10948 13574
rect 11004 13572 11028 13574
rect 11084 13572 11090 13574
rect 10782 13563 11090 13572
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 10968 13320 11020 13326
rect 11072 13308 11100 13466
rect 11164 13462 11192 14758
rect 11256 14278 11284 14962
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11256 13938 11284 14214
rect 11348 14074 11376 14962
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11624 14074 11652 14554
rect 11808 14346 11836 14758
rect 11796 14340 11848 14346
rect 11796 14282 11848 14288
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11886 14104 11942 14113
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11612 14068 11664 14074
rect 11886 14039 11888 14048
rect 11612 14010 11664 14016
rect 11940 14039 11942 14048
rect 11888 14010 11940 14016
rect 11244 13932 11296 13938
rect 11244 13874 11296 13880
rect 11796 13932 11848 13938
rect 11992 13920 12020 14214
rect 11848 13892 12020 13920
rect 11796 13874 11848 13880
rect 11152 13456 11204 13462
rect 11152 13398 11204 13404
rect 11020 13280 11100 13308
rect 10968 13262 11020 13268
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10612 12238 10640 12718
rect 10782 12540 11090 12549
rect 10782 12538 10788 12540
rect 10844 12538 10868 12540
rect 10924 12538 10948 12540
rect 11004 12538 11028 12540
rect 11084 12538 11090 12540
rect 10844 12486 10846 12538
rect 11026 12486 11028 12538
rect 10782 12484 10788 12486
rect 10844 12484 10868 12486
rect 10924 12484 10948 12486
rect 11004 12484 11028 12486
rect 11084 12484 11090 12486
rect 10782 12475 11090 12484
rect 11256 12434 11284 13874
rect 11808 13530 11836 13874
rect 12360 13734 12388 14758
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 12452 13394 12480 14962
rect 12544 14958 12572 15438
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 12748 15260 13056 15269
rect 12748 15258 12754 15260
rect 12810 15258 12834 15260
rect 12890 15258 12914 15260
rect 12970 15258 12994 15260
rect 13050 15258 13056 15260
rect 12810 15206 12812 15258
rect 12992 15206 12994 15258
rect 12748 15204 12754 15206
rect 12810 15204 12834 15206
rect 12890 15204 12914 15206
rect 12970 15204 12994 15206
rect 13050 15204 13056 15206
rect 12748 15195 13056 15204
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12544 13326 12572 14214
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 11428 13252 11480 13258
rect 11428 13194 11480 13200
rect 11440 12918 11468 13194
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 11428 12912 11480 12918
rect 11428 12854 11480 12860
rect 12452 12850 12480 13126
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 11256 12406 11468 12434
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10428 10742 10456 11494
rect 10782 11452 11090 11461
rect 10782 11450 10788 11452
rect 10844 11450 10868 11452
rect 10924 11450 10948 11452
rect 11004 11450 11028 11452
rect 11084 11450 11090 11452
rect 10844 11398 10846 11450
rect 11026 11398 11028 11450
rect 10782 11396 10788 11398
rect 10844 11396 10868 11398
rect 10924 11396 10948 11398
rect 11004 11396 11028 11398
rect 11084 11396 11090 11398
rect 10782 11387 11090 11396
rect 11256 11218 11284 12106
rect 11440 11218 11468 12406
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 10416 10736 10468 10742
rect 10416 10678 10468 10684
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9876 9042 9904 9318
rect 10336 9042 10364 10406
rect 10428 9994 10456 10678
rect 11072 10674 11100 10950
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11164 10470 11192 11086
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 10782 10364 11090 10373
rect 10782 10362 10788 10364
rect 10844 10362 10868 10364
rect 10924 10362 10948 10364
rect 11004 10362 11028 10364
rect 11084 10362 11090 10364
rect 10844 10310 10846 10362
rect 11026 10310 11028 10362
rect 10782 10308 10788 10310
rect 10844 10308 10868 10310
rect 10924 10308 10948 10310
rect 11004 10308 11028 10310
rect 11084 10308 11090 10310
rect 10782 10299 11090 10308
rect 10416 9988 10468 9994
rect 10416 9930 10468 9936
rect 10782 9276 11090 9285
rect 10782 9274 10788 9276
rect 10844 9274 10868 9276
rect 10924 9274 10948 9276
rect 11004 9274 11028 9276
rect 11084 9274 11090 9276
rect 10844 9222 10846 9274
rect 11026 9222 11028 9274
rect 10782 9220 10788 9222
rect 10844 9220 10868 9222
rect 10924 9220 10948 9222
rect 11004 9220 11028 9222
rect 11084 9220 11090 9222
rect 10782 9211 11090 9220
rect 11256 9058 11284 11154
rect 11440 10266 11468 11154
rect 12452 11082 12480 12038
rect 12544 11778 12572 12310
rect 12636 12170 12664 14758
rect 13096 14414 13124 14894
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 12748 14172 13056 14181
rect 12748 14170 12754 14172
rect 12810 14170 12834 14172
rect 12890 14170 12914 14172
rect 12970 14170 12994 14172
rect 13050 14170 13056 14172
rect 12810 14118 12812 14170
rect 12992 14118 12994 14170
rect 12748 14116 12754 14118
rect 12810 14116 12834 14118
rect 12890 14116 12914 14118
rect 12970 14116 12994 14118
rect 13050 14116 13056 14118
rect 12748 14107 13056 14116
rect 13188 14006 13216 14214
rect 13176 14000 13228 14006
rect 13176 13942 13228 13948
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12728 13190 12756 13874
rect 13280 13802 13308 15302
rect 13832 15026 13860 15302
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 13268 13796 13320 13802
rect 13268 13738 13320 13744
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12748 13084 13056 13093
rect 12748 13082 12754 13084
rect 12810 13082 12834 13084
rect 12890 13082 12914 13084
rect 12970 13082 12994 13084
rect 13050 13082 13056 13084
rect 12810 13030 12812 13082
rect 12992 13030 12994 13082
rect 12748 13028 12754 13030
rect 12810 13028 12834 13030
rect 12890 13028 12914 13030
rect 12970 13028 12994 13030
rect 13050 13028 13056 13030
rect 12748 13019 13056 13028
rect 13096 12918 13124 13670
rect 13188 12918 13216 13670
rect 13648 13326 13676 13874
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 13176 12912 13228 12918
rect 13176 12854 13228 12860
rect 13648 12782 13676 13262
rect 13832 12986 13860 13670
rect 13924 13394 13952 15846
rect 14715 15804 15023 15813
rect 14715 15802 14721 15804
rect 14777 15802 14801 15804
rect 14857 15802 14881 15804
rect 14937 15802 14961 15804
rect 15017 15802 15023 15804
rect 14777 15750 14779 15802
rect 14959 15750 14961 15802
rect 14715 15748 14721 15750
rect 14777 15748 14801 15750
rect 14857 15748 14881 15750
rect 14937 15748 14961 15750
rect 15017 15748 15023 15750
rect 14715 15739 15023 15748
rect 14004 15496 14056 15502
rect 14004 15438 14056 15444
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12748 11996 13056 12005
rect 12748 11994 12754 11996
rect 12810 11994 12834 11996
rect 12890 11994 12914 11996
rect 12970 11994 12994 11996
rect 13050 11994 13056 11996
rect 12810 11942 12812 11994
rect 12992 11942 12994 11994
rect 12748 11940 12754 11942
rect 12810 11940 12834 11942
rect 12890 11940 12914 11942
rect 12970 11940 12994 11942
rect 13050 11940 13056 11942
rect 12748 11931 13056 11940
rect 13372 11898 13400 12174
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 12544 11750 12756 11778
rect 12728 11150 12756 11750
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13280 11286 13308 11562
rect 13268 11280 13320 11286
rect 13268 11222 13320 11228
rect 13372 11150 13400 11834
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13464 11150 13492 11290
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12748 10908 13056 10917
rect 12748 10906 12754 10908
rect 12810 10906 12834 10908
rect 12890 10906 12914 10908
rect 12970 10906 12994 10908
rect 13050 10906 13056 10908
rect 12810 10854 12812 10906
rect 12992 10854 12994 10906
rect 12748 10852 12754 10854
rect 12810 10852 12834 10854
rect 12890 10852 12914 10854
rect 12970 10852 12994 10854
rect 13050 10852 13056 10854
rect 12748 10843 13056 10852
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11428 9444 11480 9450
rect 11428 9386 11480 9392
rect 11256 9042 11376 9058
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 10324 9036 10376 9042
rect 11256 9036 11388 9042
rect 11256 9030 11336 9036
rect 10324 8978 10376 8984
rect 11336 8978 11388 8984
rect 11440 8974 11468 9386
rect 11808 9178 11836 10610
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13556 10062 13584 10406
rect 13648 10062 13676 11494
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13832 10538 13860 10950
rect 13924 10674 13952 12038
rect 14016 11830 14044 15438
rect 16681 15260 16989 15269
rect 16681 15258 16687 15260
rect 16743 15258 16767 15260
rect 16823 15258 16847 15260
rect 16903 15258 16927 15260
rect 16983 15258 16989 15260
rect 16743 15206 16745 15258
rect 16925 15206 16927 15258
rect 16681 15204 16687 15206
rect 16743 15204 16767 15206
rect 16823 15204 16847 15206
rect 16903 15204 16927 15206
rect 16983 15204 16989 15206
rect 16681 15195 16989 15204
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 14715 14716 15023 14725
rect 14715 14714 14721 14716
rect 14777 14714 14801 14716
rect 14857 14714 14881 14716
rect 14937 14714 14961 14716
rect 15017 14714 15023 14716
rect 14777 14662 14779 14714
rect 14959 14662 14961 14714
rect 14715 14660 14721 14662
rect 14777 14660 14801 14662
rect 14857 14660 14881 14662
rect 14937 14660 14961 14662
rect 15017 14660 15023 14662
rect 14715 14651 15023 14660
rect 15120 14278 15148 14758
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14094 13968 14150 13977
rect 14094 13903 14150 13912
rect 14108 12986 14136 13903
rect 14568 13530 14596 14010
rect 14715 13628 15023 13637
rect 14715 13626 14721 13628
rect 14777 13626 14801 13628
rect 14857 13626 14881 13628
rect 14937 13626 14961 13628
rect 15017 13626 15023 13628
rect 14777 13574 14779 13626
rect 14959 13574 14961 13626
rect 14715 13572 14721 13574
rect 14777 13572 14801 13574
rect 14857 13572 14881 13574
rect 14937 13572 14961 13574
rect 15017 13572 15023 13574
rect 14715 13563 15023 13572
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 14200 11694 14228 13126
rect 14292 12850 14320 13126
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14476 12238 14504 13262
rect 14715 12540 15023 12549
rect 14715 12538 14721 12540
rect 14777 12538 14801 12540
rect 14857 12538 14881 12540
rect 14937 12538 14961 12540
rect 15017 12538 15023 12540
rect 14777 12486 14779 12538
rect 14959 12486 14961 12538
rect 14715 12484 14721 12486
rect 14777 12484 14801 12486
rect 14857 12484 14881 12486
rect 14937 12484 14961 12486
rect 15017 12484 15023 12486
rect 14715 12475 15023 12484
rect 15120 12238 15148 14214
rect 16681 14172 16989 14181
rect 16681 14170 16687 14172
rect 16743 14170 16767 14172
rect 16823 14170 16847 14172
rect 16903 14170 16927 14172
rect 16983 14170 16989 14172
rect 16743 14118 16745 14170
rect 16925 14118 16927 14170
rect 16681 14116 16687 14118
rect 16743 14116 16767 14118
rect 16823 14116 16847 14118
rect 16903 14116 16927 14118
rect 16983 14116 16989 14118
rect 16681 14107 16989 14116
rect 16681 13084 16989 13093
rect 16681 13082 16687 13084
rect 16743 13082 16767 13084
rect 16823 13082 16847 13084
rect 16903 13082 16927 13084
rect 16983 13082 16989 13084
rect 16743 13030 16745 13082
rect 16925 13030 16927 13082
rect 16681 13028 16687 13030
rect 16743 13028 16767 13030
rect 16823 13028 16847 13030
rect 16903 13028 16927 13030
rect 16983 13028 16989 13030
rect 16681 13019 16989 13028
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14384 11830 14412 12038
rect 14372 11824 14424 11830
rect 14372 11766 14424 11772
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 14476 11286 14504 12174
rect 14715 11452 15023 11461
rect 14715 11450 14721 11452
rect 14777 11450 14801 11452
rect 14857 11450 14881 11452
rect 14937 11450 14961 11452
rect 15017 11450 15023 11452
rect 14777 11398 14779 11450
rect 14959 11398 14961 11450
rect 14715 11396 14721 11398
rect 14777 11396 14801 11398
rect 14857 11396 14881 11398
rect 14937 11396 14961 11398
rect 15017 11396 15023 11398
rect 14715 11387 15023 11396
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 13820 10532 13872 10538
rect 13820 10474 13872 10480
rect 14200 10266 14228 10542
rect 14715 10364 15023 10373
rect 14715 10362 14721 10364
rect 14777 10362 14801 10364
rect 14857 10362 14881 10364
rect 14937 10362 14961 10364
rect 15017 10362 15023 10364
rect 14777 10310 14779 10362
rect 14959 10310 14961 10362
rect 14715 10308 14721 10310
rect 14777 10308 14801 10310
rect 14857 10308 14881 10310
rect 14937 10308 14961 10310
rect 15017 10308 15023 10310
rect 14715 10299 15023 10308
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 15120 10198 15148 12174
rect 16681 11996 16989 12005
rect 16681 11994 16687 11996
rect 16743 11994 16767 11996
rect 16823 11994 16847 11996
rect 16903 11994 16927 11996
rect 16983 11994 16989 11996
rect 16743 11942 16745 11994
rect 16925 11942 16927 11994
rect 16681 11940 16687 11942
rect 16743 11940 16767 11942
rect 16823 11940 16847 11942
rect 16903 11940 16927 11942
rect 16983 11940 16989 11942
rect 16681 11931 16989 11940
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 15672 10742 15700 11018
rect 15660 10736 15712 10742
rect 15660 10678 15712 10684
rect 16132 10674 16160 11086
rect 16681 10908 16989 10917
rect 16681 10906 16687 10908
rect 16743 10906 16767 10908
rect 16823 10906 16847 10908
rect 16903 10906 16927 10908
rect 16983 10906 16989 10908
rect 16743 10854 16745 10906
rect 16925 10854 16927 10906
rect 16681 10852 16687 10854
rect 16743 10852 16767 10854
rect 16823 10852 16847 10854
rect 16903 10852 16927 10854
rect 16983 10852 16989 10854
rect 16681 10843 16989 10852
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 15108 10192 15160 10198
rect 15108 10134 15160 10140
rect 16132 10130 16160 10610
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 12748 9820 13056 9829
rect 12748 9818 12754 9820
rect 12810 9818 12834 9820
rect 12890 9818 12914 9820
rect 12970 9818 12994 9820
rect 13050 9818 13056 9820
rect 12810 9766 12812 9818
rect 12992 9766 12994 9818
rect 12748 9764 12754 9766
rect 12810 9764 12834 9766
rect 12890 9764 12914 9766
rect 12970 9764 12994 9766
rect 13050 9764 13056 9766
rect 12748 9755 13056 9764
rect 14200 9586 14228 9862
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 12360 8974 12388 9386
rect 13464 9178 13492 9454
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13740 9110 13768 9454
rect 14715 9276 15023 9285
rect 14715 9274 14721 9276
rect 14777 9274 14801 9276
rect 14857 9274 14881 9276
rect 14937 9274 14961 9276
rect 15017 9274 15023 9276
rect 14777 9222 14779 9274
rect 14959 9222 14961 9274
rect 14715 9220 14721 9222
rect 14777 9220 14801 9222
rect 14857 9220 14881 9222
rect 14937 9220 14961 9222
rect 15017 9220 15023 9222
rect 14715 9211 15023 9220
rect 15120 9178 15148 9454
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 13728 9104 13780 9110
rect 13728 9046 13780 9052
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9784 8090 9812 8434
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8404 5846 8432 6122
rect 8496 6118 8524 6258
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 7760 4214 7788 4490
rect 8496 4214 8524 5510
rect 8815 5468 9123 5477
rect 8815 5466 8821 5468
rect 8877 5466 8901 5468
rect 8957 5466 8981 5468
rect 9037 5466 9061 5468
rect 9117 5466 9123 5468
rect 8877 5414 8879 5466
rect 9059 5414 9061 5466
rect 8815 5412 8821 5414
rect 8877 5412 8901 5414
rect 8957 5412 8981 5414
rect 9037 5412 9061 5414
rect 9117 5412 9123 5414
rect 8815 5403 9123 5412
rect 9324 4622 9352 6258
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5778 9536 6054
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9404 5704 9456 5710
rect 9600 5658 9628 6326
rect 9784 5778 9812 7482
rect 10060 7478 10088 7754
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9876 6322 9904 7346
rect 10244 7206 10272 8842
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 10782 8188 11090 8197
rect 10782 8186 10788 8188
rect 10844 8186 10868 8188
rect 10924 8186 10948 8188
rect 11004 8186 11028 8188
rect 11084 8186 11090 8188
rect 10844 8134 10846 8186
rect 11026 8134 11028 8186
rect 10782 8132 10788 8134
rect 10844 8132 10868 8134
rect 10924 8132 10948 8134
rect 11004 8132 11028 8134
rect 11084 8132 11090 8134
rect 10782 8123 11090 8132
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10336 7002 10364 7346
rect 10782 7100 11090 7109
rect 10782 7098 10788 7100
rect 10844 7098 10868 7100
rect 10924 7098 10948 7100
rect 11004 7098 11028 7100
rect 11084 7098 11090 7100
rect 10844 7046 10846 7098
rect 11026 7046 11028 7098
rect 10782 7044 10788 7046
rect 10844 7044 10868 7046
rect 10924 7044 10948 7046
rect 11004 7044 11028 7046
rect 11084 7044 11090 7046
rect 10782 7035 11090 7044
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10152 6458 10180 6598
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9456 5652 9628 5658
rect 9404 5646 9628 5652
rect 9416 5630 9628 5646
rect 9600 5302 9628 5630
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9784 4826 9812 5714
rect 10152 5574 10180 6394
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10152 5234 10180 5510
rect 10336 5370 10364 6938
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11164 6458 11192 6666
rect 11256 6662 11284 8434
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11348 7818 11376 8298
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10520 5642 10548 6122
rect 10782 6012 11090 6021
rect 10782 6010 10788 6012
rect 10844 6010 10868 6012
rect 10924 6010 10948 6012
rect 11004 6010 11028 6012
rect 11084 6010 11090 6012
rect 10844 5958 10846 6010
rect 11026 5958 11028 6010
rect 10782 5956 10788 5958
rect 10844 5956 10868 5958
rect 10924 5956 10948 5958
rect 11004 5956 11028 5958
rect 11084 5956 11090 5958
rect 10782 5947 11090 5956
rect 11256 5914 11284 6598
rect 11716 6322 11744 8434
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 12084 7954 12112 8230
rect 12360 8090 12388 8910
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 12748 8732 13056 8741
rect 12748 8730 12754 8732
rect 12810 8730 12834 8732
rect 12890 8730 12914 8732
rect 12970 8730 12994 8732
rect 13050 8730 13056 8732
rect 12810 8678 12812 8730
rect 12992 8678 12994 8730
rect 12748 8676 12754 8678
rect 12810 8676 12834 8678
rect 12890 8676 12914 8678
rect 12970 8676 12994 8678
rect 13050 8676 13056 8678
rect 12748 8667 13056 8676
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 11900 7546 11928 7754
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 12360 7478 12388 8026
rect 12912 7886 12940 8230
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 12748 7644 13056 7653
rect 12748 7642 12754 7644
rect 12810 7642 12834 7644
rect 12890 7642 12914 7644
rect 12970 7642 12994 7644
rect 13050 7642 13056 7644
rect 12810 7590 12812 7642
rect 12992 7590 12994 7642
rect 12748 7588 12754 7590
rect 12810 7588 12834 7590
rect 12890 7588 12914 7590
rect 12970 7588 12994 7590
rect 13050 7588 13056 7590
rect 12748 7579 13056 7588
rect 12348 7472 12400 7478
rect 12348 7414 12400 7420
rect 13096 6798 13124 7822
rect 13280 7410 13308 8842
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14660 8498 14688 8774
rect 15488 8634 15516 9590
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15580 8974 15608 9318
rect 16132 8974 16160 10066
rect 16224 9722 16252 10406
rect 16681 9820 16989 9829
rect 16681 9818 16687 9820
rect 16743 9818 16767 9820
rect 16823 9818 16847 9820
rect 16903 9818 16927 9820
rect 16983 9818 16989 9820
rect 16743 9766 16745 9818
rect 16925 9766 16927 9818
rect 16681 9764 16687 9766
rect 16743 9764 16767 9766
rect 16823 9764 16847 9766
rect 16903 9764 16927 9766
rect 16983 9764 16989 9766
rect 16681 9755 16989 9764
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15856 8566 15884 8774
rect 15844 8560 15896 8566
rect 15844 8502 15896 8508
rect 16132 8498 16160 8910
rect 16681 8732 16989 8741
rect 16681 8730 16687 8732
rect 16743 8730 16767 8732
rect 16823 8730 16847 8732
rect 16903 8730 16927 8732
rect 16983 8730 16989 8732
rect 16743 8678 16745 8730
rect 16925 8678 16927 8730
rect 16681 8676 16687 8678
rect 16743 8676 16767 8678
rect 16823 8676 16847 8678
rect 16903 8676 16927 8678
rect 16983 8676 16989 8678
rect 16681 8667 16989 8676
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14384 8090 14412 8366
rect 14715 8188 15023 8197
rect 14715 8186 14721 8188
rect 14777 8186 14801 8188
rect 14857 8186 14881 8188
rect 14937 8186 14961 8188
rect 15017 8186 15023 8188
rect 14777 8134 14779 8186
rect 14959 8134 14961 8186
rect 14715 8132 14721 8134
rect 14777 8132 14801 8134
rect 14857 8132 14881 8134
rect 14937 8132 14961 8134
rect 15017 8132 15023 8134
rect 14715 8123 15023 8132
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 16681 7644 16989 7653
rect 16681 7642 16687 7644
rect 16743 7642 16767 7644
rect 16823 7642 16847 7644
rect 16903 7642 16927 7644
rect 16983 7642 16989 7644
rect 16743 7590 16745 7642
rect 16925 7590 16927 7642
rect 16681 7588 16687 7590
rect 16743 7588 16767 7590
rect 16823 7588 16847 7590
rect 16903 7588 16927 7590
rect 16983 7588 16989 7590
rect 16681 7579 16989 7588
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 14715 7100 15023 7109
rect 14715 7098 14721 7100
rect 14777 7098 14801 7100
rect 14857 7098 14881 7100
rect 14937 7098 14961 7100
rect 15017 7098 15023 7100
rect 14777 7046 14779 7098
rect 14959 7046 14961 7098
rect 14715 7044 14721 7046
rect 14777 7044 14801 7046
rect 14857 7044 14881 7046
rect 14937 7044 14961 7046
rect 15017 7044 15023 7046
rect 14715 7035 15023 7044
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12748 6556 13056 6565
rect 12748 6554 12754 6556
rect 12810 6554 12834 6556
rect 12890 6554 12914 6556
rect 12970 6554 12994 6556
rect 13050 6554 13056 6556
rect 12810 6502 12812 6554
rect 12992 6502 12994 6554
rect 12748 6500 12754 6502
rect 12810 6500 12834 6502
rect 12890 6500 12914 6502
rect 12970 6500 12994 6502
rect 13050 6500 13056 6502
rect 12748 6491 13056 6500
rect 16681 6556 16989 6565
rect 16681 6554 16687 6556
rect 16743 6554 16767 6556
rect 16823 6554 16847 6556
rect 16903 6554 16927 6556
rect 16983 6554 16989 6556
rect 16743 6502 16745 6554
rect 16925 6502 16927 6554
rect 16681 6500 16687 6502
rect 16743 6500 16767 6502
rect 16823 6500 16847 6502
rect 16903 6500 16927 6502
rect 16983 6500 16989 6502
rect 16681 6491 16989 6500
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 14715 6012 15023 6021
rect 14715 6010 14721 6012
rect 14777 6010 14801 6012
rect 14857 6010 14881 6012
rect 14937 6010 14961 6012
rect 15017 6010 15023 6012
rect 14777 5958 14779 6010
rect 14959 5958 14961 6010
rect 14715 5956 14721 5958
rect 14777 5956 14801 5958
rect 14857 5956 14881 5958
rect 14937 5956 14961 5958
rect 15017 5956 15023 5958
rect 14715 5947 15023 5956
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10782 4924 11090 4933
rect 10782 4922 10788 4924
rect 10844 4922 10868 4924
rect 10924 4922 10948 4924
rect 11004 4922 11028 4924
rect 11084 4922 11090 4924
rect 10844 4870 10846 4922
rect 11026 4870 11028 4922
rect 10782 4868 10788 4870
rect 10844 4868 10868 4870
rect 10924 4868 10948 4870
rect 11004 4868 11028 4870
rect 11084 4868 11090 4870
rect 10782 4859 11090 4868
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 11256 4622 11284 5850
rect 12748 5468 13056 5477
rect 12748 5466 12754 5468
rect 12810 5466 12834 5468
rect 12890 5466 12914 5468
rect 12970 5466 12994 5468
rect 13050 5466 13056 5468
rect 12810 5414 12812 5466
rect 12992 5414 12994 5466
rect 12748 5412 12754 5414
rect 12810 5412 12834 5414
rect 12890 5412 12914 5414
rect 12970 5412 12994 5414
rect 13050 5412 13056 5414
rect 12748 5403 13056 5412
rect 16681 5468 16989 5477
rect 16681 5466 16687 5468
rect 16743 5466 16767 5468
rect 16823 5466 16847 5468
rect 16903 5466 16927 5468
rect 16983 5466 16989 5468
rect 16743 5414 16745 5466
rect 16925 5414 16927 5466
rect 16681 5412 16687 5414
rect 16743 5412 16767 5414
rect 16823 5412 16847 5414
rect 16903 5412 16927 5414
rect 16983 5412 16989 5414
rect 16681 5403 16989 5412
rect 14715 4924 15023 4933
rect 14715 4922 14721 4924
rect 14777 4922 14801 4924
rect 14857 4922 14881 4924
rect 14937 4922 14961 4924
rect 15017 4922 15023 4924
rect 14777 4870 14779 4922
rect 14959 4870 14961 4922
rect 14715 4868 14721 4870
rect 14777 4868 14801 4870
rect 14857 4868 14881 4870
rect 14937 4868 14961 4870
rect 15017 4868 15023 4870
rect 14715 4859 15023 4868
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 8815 4380 9123 4389
rect 8815 4378 8821 4380
rect 8877 4378 8901 4380
rect 8957 4378 8981 4380
rect 9037 4378 9061 4380
rect 9117 4378 9123 4380
rect 8877 4326 8879 4378
rect 9059 4326 9061 4378
rect 8815 4324 8821 4326
rect 8877 4324 8901 4326
rect 8957 4324 8981 4326
rect 9037 4324 9061 4326
rect 9117 4324 9123 4326
rect 8815 4315 9123 4324
rect 7748 4208 7800 4214
rect 7748 4150 7800 4156
rect 8484 4208 8536 4214
rect 8484 4150 8536 4156
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 9324 4078 9352 4558
rect 12748 4380 13056 4389
rect 12748 4378 12754 4380
rect 12810 4378 12834 4380
rect 12890 4378 12914 4380
rect 12970 4378 12994 4380
rect 13050 4378 13056 4380
rect 12810 4326 12812 4378
rect 12992 4326 12994 4378
rect 12748 4324 12754 4326
rect 12810 4324 12834 4326
rect 12890 4324 12914 4326
rect 12970 4324 12994 4326
rect 13050 4324 13056 4326
rect 12748 4315 13056 4324
rect 16681 4380 16989 4389
rect 16681 4378 16687 4380
rect 16743 4378 16767 4380
rect 16823 4378 16847 4380
rect 16903 4378 16927 4380
rect 16983 4378 16989 4380
rect 16743 4326 16745 4378
rect 16925 4326 16927 4378
rect 16681 4324 16687 4326
rect 16743 4324 16767 4326
rect 16823 4324 16847 4326
rect 16903 4324 16927 4326
rect 16983 4324 16989 4326
rect 16681 4315 16989 4324
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 6849 3836 7157 3845
rect 6849 3834 6855 3836
rect 6911 3834 6935 3836
rect 6991 3834 7015 3836
rect 7071 3834 7095 3836
rect 7151 3834 7157 3836
rect 6911 3782 6913 3834
rect 7093 3782 7095 3834
rect 6849 3780 6855 3782
rect 6911 3780 6935 3782
rect 6991 3780 7015 3782
rect 7071 3780 7095 3782
rect 7151 3780 7157 3782
rect 6849 3771 7157 3780
rect 10782 3836 11090 3845
rect 10782 3834 10788 3836
rect 10844 3834 10868 3836
rect 10924 3834 10948 3836
rect 11004 3834 11028 3836
rect 11084 3834 11090 3836
rect 10844 3782 10846 3834
rect 11026 3782 11028 3834
rect 10782 3780 10788 3782
rect 10844 3780 10868 3782
rect 10924 3780 10948 3782
rect 11004 3780 11028 3782
rect 11084 3780 11090 3782
rect 10782 3771 11090 3780
rect 14715 3836 15023 3845
rect 14715 3834 14721 3836
rect 14777 3834 14801 3836
rect 14857 3834 14881 3836
rect 14937 3834 14961 3836
rect 15017 3834 15023 3836
rect 14777 3782 14779 3834
rect 14959 3782 14961 3834
rect 14715 3780 14721 3782
rect 14777 3780 14801 3782
rect 14857 3780 14881 3782
rect 14937 3780 14961 3782
rect 15017 3780 15023 3782
rect 14715 3771 15023 3780
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4882 3292 5190 3301
rect 4882 3290 4888 3292
rect 4944 3290 4968 3292
rect 5024 3290 5048 3292
rect 5104 3290 5128 3292
rect 5184 3290 5190 3292
rect 4944 3238 4946 3290
rect 5126 3238 5128 3290
rect 4882 3236 4888 3238
rect 4944 3236 4968 3238
rect 5024 3236 5048 3238
rect 5104 3236 5128 3238
rect 5184 3236 5190 3238
rect 4882 3227 5190 3236
rect 8815 3292 9123 3301
rect 8815 3290 8821 3292
rect 8877 3290 8901 3292
rect 8957 3290 8981 3292
rect 9037 3290 9061 3292
rect 9117 3290 9123 3292
rect 8877 3238 8879 3290
rect 9059 3238 9061 3290
rect 8815 3236 8821 3238
rect 8877 3236 8901 3238
rect 8957 3236 8981 3238
rect 9037 3236 9061 3238
rect 9117 3236 9123 3238
rect 8815 3227 9123 3236
rect 12748 3292 13056 3301
rect 12748 3290 12754 3292
rect 12810 3290 12834 3292
rect 12890 3290 12914 3292
rect 12970 3290 12994 3292
rect 13050 3290 13056 3292
rect 12810 3238 12812 3290
rect 12992 3238 12994 3290
rect 12748 3236 12754 3238
rect 12810 3236 12834 3238
rect 12890 3236 12914 3238
rect 12970 3236 12994 3238
rect 13050 3236 13056 3238
rect 12748 3227 13056 3236
rect 16681 3292 16989 3301
rect 16681 3290 16687 3292
rect 16743 3290 16767 3292
rect 16823 3290 16847 3292
rect 16903 3290 16927 3292
rect 16983 3290 16989 3292
rect 16743 3238 16745 3290
rect 16925 3238 16927 3290
rect 16681 3236 16687 3238
rect 16743 3236 16767 3238
rect 16823 3236 16847 3238
rect 16903 3236 16927 3238
rect 16983 3236 16989 3238
rect 16681 3227 16989 3236
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 2916 2748 3224 2757
rect 2916 2746 2922 2748
rect 2978 2746 3002 2748
rect 3058 2746 3082 2748
rect 3138 2746 3162 2748
rect 3218 2746 3224 2748
rect 2978 2694 2980 2746
rect 3160 2694 3162 2746
rect 2916 2692 2922 2694
rect 2978 2692 3002 2694
rect 3058 2692 3082 2694
rect 3138 2692 3162 2694
rect 3218 2692 3224 2694
rect 2916 2683 3224 2692
rect 6849 2748 7157 2757
rect 6849 2746 6855 2748
rect 6911 2746 6935 2748
rect 6991 2746 7015 2748
rect 7071 2746 7095 2748
rect 7151 2746 7157 2748
rect 6911 2694 6913 2746
rect 7093 2694 7095 2746
rect 6849 2692 6855 2694
rect 6911 2692 6935 2694
rect 6991 2692 7015 2694
rect 7071 2692 7095 2694
rect 7151 2692 7157 2694
rect 6849 2683 7157 2692
rect 10782 2748 11090 2757
rect 10782 2746 10788 2748
rect 10844 2746 10868 2748
rect 10924 2746 10948 2748
rect 11004 2746 11028 2748
rect 11084 2746 11090 2748
rect 10844 2694 10846 2746
rect 11026 2694 11028 2746
rect 10782 2692 10788 2694
rect 10844 2692 10868 2694
rect 10924 2692 10948 2694
rect 11004 2692 11028 2694
rect 11084 2692 11090 2694
rect 10782 2683 11090 2692
rect 14715 2748 15023 2757
rect 14715 2746 14721 2748
rect 14777 2746 14801 2748
rect 14857 2746 14881 2748
rect 14937 2746 14961 2748
rect 15017 2746 15023 2748
rect 14777 2694 14779 2746
rect 14959 2694 14961 2746
rect 14715 2692 14721 2694
rect 14777 2692 14801 2694
rect 14857 2692 14881 2694
rect 14937 2692 14961 2694
rect 15017 2692 15023 2694
rect 14715 2683 15023 2692
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1768 2304 1820 2310
rect 1766 2272 1768 2281
rect 1820 2272 1822 2281
rect 1766 2207 1822 2216
rect 4882 2204 5190 2213
rect 4882 2202 4888 2204
rect 4944 2202 4968 2204
rect 5024 2202 5048 2204
rect 5104 2202 5128 2204
rect 5184 2202 5190 2204
rect 4944 2150 4946 2202
rect 5126 2150 5128 2202
rect 4882 2148 4888 2150
rect 4944 2148 4968 2150
rect 5024 2148 5048 2150
rect 5104 2148 5128 2150
rect 5184 2148 5190 2150
rect 4882 2139 5190 2148
rect 8815 2204 9123 2213
rect 8815 2202 8821 2204
rect 8877 2202 8901 2204
rect 8957 2202 8981 2204
rect 9037 2202 9061 2204
rect 9117 2202 9123 2204
rect 8877 2150 8879 2202
rect 9059 2150 9061 2202
rect 8815 2148 8821 2150
rect 8877 2148 8901 2150
rect 8957 2148 8981 2150
rect 9037 2148 9061 2150
rect 9117 2148 9123 2150
rect 8815 2139 9123 2148
rect 12748 2204 13056 2213
rect 12748 2202 12754 2204
rect 12810 2202 12834 2204
rect 12890 2202 12914 2204
rect 12970 2202 12994 2204
rect 13050 2202 13056 2204
rect 12810 2150 12812 2202
rect 12992 2150 12994 2202
rect 12748 2148 12754 2150
rect 12810 2148 12834 2150
rect 12890 2148 12914 2150
rect 12970 2148 12994 2150
rect 13050 2148 13056 2150
rect 12748 2139 13056 2148
rect 16681 2204 16989 2213
rect 16681 2202 16687 2204
rect 16743 2202 16767 2204
rect 16823 2202 16847 2204
rect 16903 2202 16927 2204
rect 16983 2202 16989 2204
rect 16743 2150 16745 2202
rect 16925 2150 16927 2202
rect 16681 2148 16687 2150
rect 16743 2148 16767 2150
rect 16823 2148 16847 2150
rect 16903 2148 16927 2150
rect 16983 2148 16989 2150
rect 16681 2139 16989 2148
rect 1398 776 1454 785
rect 1398 711 1454 720
<< via2 >>
rect 4158 17176 4214 17232
rect 2922 15802 2978 15804
rect 3002 15802 3058 15804
rect 3082 15802 3138 15804
rect 3162 15802 3218 15804
rect 2922 15750 2968 15802
rect 2968 15750 2978 15802
rect 3002 15750 3032 15802
rect 3032 15750 3044 15802
rect 3044 15750 3058 15802
rect 3082 15750 3096 15802
rect 3096 15750 3108 15802
rect 3108 15750 3138 15802
rect 3162 15750 3172 15802
rect 3172 15750 3218 15802
rect 2922 15748 2978 15750
rect 3002 15748 3058 15750
rect 3082 15748 3138 15750
rect 3162 15748 3218 15750
rect 2778 15700 2834 15736
rect 2778 15680 2780 15700
rect 2780 15680 2832 15700
rect 2832 15680 2834 15700
rect 1674 14184 1730 14240
rect 1674 12688 1730 12744
rect 2922 14714 2978 14716
rect 3002 14714 3058 14716
rect 3082 14714 3138 14716
rect 3162 14714 3218 14716
rect 2922 14662 2968 14714
rect 2968 14662 2978 14714
rect 3002 14662 3032 14714
rect 3032 14662 3044 14714
rect 3044 14662 3058 14714
rect 3082 14662 3096 14714
rect 3096 14662 3108 14714
rect 3108 14662 3138 14714
rect 3162 14662 3172 14714
rect 3172 14662 3218 14714
rect 2922 14660 2978 14662
rect 3002 14660 3058 14662
rect 3082 14660 3138 14662
rect 3162 14660 3218 14662
rect 2922 13626 2978 13628
rect 3002 13626 3058 13628
rect 3082 13626 3138 13628
rect 3162 13626 3218 13628
rect 2922 13574 2968 13626
rect 2968 13574 2978 13626
rect 3002 13574 3032 13626
rect 3032 13574 3044 13626
rect 3044 13574 3058 13626
rect 3082 13574 3096 13626
rect 3096 13574 3108 13626
rect 3108 13574 3138 13626
rect 3162 13574 3172 13626
rect 3172 13574 3218 13626
rect 2922 13572 2978 13574
rect 3002 13572 3058 13574
rect 3082 13572 3138 13574
rect 3162 13572 3218 13574
rect 6855 15802 6911 15804
rect 6935 15802 6991 15804
rect 7015 15802 7071 15804
rect 7095 15802 7151 15804
rect 6855 15750 6901 15802
rect 6901 15750 6911 15802
rect 6935 15750 6965 15802
rect 6965 15750 6977 15802
rect 6977 15750 6991 15802
rect 7015 15750 7029 15802
rect 7029 15750 7041 15802
rect 7041 15750 7071 15802
rect 7095 15750 7105 15802
rect 7105 15750 7151 15802
rect 6855 15748 6911 15750
rect 6935 15748 6991 15750
rect 7015 15748 7071 15750
rect 7095 15748 7151 15750
rect 10788 15802 10844 15804
rect 10868 15802 10924 15804
rect 10948 15802 11004 15804
rect 11028 15802 11084 15804
rect 10788 15750 10834 15802
rect 10834 15750 10844 15802
rect 10868 15750 10898 15802
rect 10898 15750 10910 15802
rect 10910 15750 10924 15802
rect 10948 15750 10962 15802
rect 10962 15750 10974 15802
rect 10974 15750 11004 15802
rect 11028 15750 11038 15802
rect 11038 15750 11084 15802
rect 10788 15748 10844 15750
rect 10868 15748 10924 15750
rect 10948 15748 11004 15750
rect 11028 15748 11084 15750
rect 4888 15258 4944 15260
rect 4968 15258 5024 15260
rect 5048 15258 5104 15260
rect 5128 15258 5184 15260
rect 4888 15206 4934 15258
rect 4934 15206 4944 15258
rect 4968 15206 4998 15258
rect 4998 15206 5010 15258
rect 5010 15206 5024 15258
rect 5048 15206 5062 15258
rect 5062 15206 5074 15258
rect 5074 15206 5104 15258
rect 5128 15206 5138 15258
rect 5138 15206 5184 15258
rect 4888 15204 4944 15206
rect 4968 15204 5024 15206
rect 5048 15204 5104 15206
rect 5128 15204 5184 15206
rect 4888 14170 4944 14172
rect 4968 14170 5024 14172
rect 5048 14170 5104 14172
rect 5128 14170 5184 14172
rect 4888 14118 4934 14170
rect 4934 14118 4944 14170
rect 4968 14118 4998 14170
rect 4998 14118 5010 14170
rect 5010 14118 5024 14170
rect 5048 14118 5062 14170
rect 5062 14118 5074 14170
rect 5074 14118 5104 14170
rect 5128 14118 5138 14170
rect 5138 14118 5184 14170
rect 4888 14116 4944 14118
rect 4968 14116 5024 14118
rect 5048 14116 5104 14118
rect 5128 14116 5184 14118
rect 4066 13948 4068 13968
rect 4068 13948 4120 13968
rect 4120 13948 4122 13968
rect 4066 13912 4122 13948
rect 2922 12538 2978 12540
rect 3002 12538 3058 12540
rect 3082 12538 3138 12540
rect 3162 12538 3218 12540
rect 2922 12486 2968 12538
rect 2968 12486 2978 12538
rect 3002 12486 3032 12538
rect 3032 12486 3044 12538
rect 3044 12486 3058 12538
rect 3082 12486 3096 12538
rect 3096 12486 3108 12538
rect 3108 12486 3138 12538
rect 3162 12486 3172 12538
rect 3172 12486 3218 12538
rect 2922 12484 2978 12486
rect 3002 12484 3058 12486
rect 3082 12484 3138 12486
rect 3162 12484 3218 12486
rect 1674 11228 1676 11248
rect 1676 11228 1728 11248
rect 1728 11228 1730 11248
rect 1674 11192 1730 11228
rect 1490 5208 1546 5264
rect 1766 9696 1822 9752
rect 1766 8200 1822 8256
rect 1674 6704 1730 6760
rect 1398 3712 1454 3768
rect 2922 11450 2978 11452
rect 3002 11450 3058 11452
rect 3082 11450 3138 11452
rect 3162 11450 3218 11452
rect 2922 11398 2968 11450
rect 2968 11398 2978 11450
rect 3002 11398 3032 11450
rect 3032 11398 3044 11450
rect 3044 11398 3058 11450
rect 3082 11398 3096 11450
rect 3096 11398 3108 11450
rect 3108 11398 3138 11450
rect 3162 11398 3172 11450
rect 3172 11398 3218 11450
rect 2922 11396 2978 11398
rect 3002 11396 3058 11398
rect 3082 11396 3138 11398
rect 3162 11396 3218 11398
rect 2922 10362 2978 10364
rect 3002 10362 3058 10364
rect 3082 10362 3138 10364
rect 3162 10362 3218 10364
rect 2922 10310 2968 10362
rect 2968 10310 2978 10362
rect 3002 10310 3032 10362
rect 3032 10310 3044 10362
rect 3044 10310 3058 10362
rect 3082 10310 3096 10362
rect 3096 10310 3108 10362
rect 3108 10310 3138 10362
rect 3162 10310 3172 10362
rect 3172 10310 3218 10362
rect 2922 10308 2978 10310
rect 3002 10308 3058 10310
rect 3082 10308 3138 10310
rect 3162 10308 3218 10310
rect 2922 9274 2978 9276
rect 3002 9274 3058 9276
rect 3082 9274 3138 9276
rect 3162 9274 3218 9276
rect 2922 9222 2968 9274
rect 2968 9222 2978 9274
rect 3002 9222 3032 9274
rect 3032 9222 3044 9274
rect 3044 9222 3058 9274
rect 3082 9222 3096 9274
rect 3096 9222 3108 9274
rect 3108 9222 3138 9274
rect 3162 9222 3172 9274
rect 3172 9222 3218 9274
rect 2922 9220 2978 9222
rect 3002 9220 3058 9222
rect 3082 9220 3138 9222
rect 3162 9220 3218 9222
rect 2922 8186 2978 8188
rect 3002 8186 3058 8188
rect 3082 8186 3138 8188
rect 3162 8186 3218 8188
rect 2922 8134 2968 8186
rect 2968 8134 2978 8186
rect 3002 8134 3032 8186
rect 3032 8134 3044 8186
rect 3044 8134 3058 8186
rect 3082 8134 3096 8186
rect 3096 8134 3108 8186
rect 3108 8134 3138 8186
rect 3162 8134 3172 8186
rect 3172 8134 3218 8186
rect 2922 8132 2978 8134
rect 3002 8132 3058 8134
rect 3082 8132 3138 8134
rect 3162 8132 3218 8134
rect 2922 7098 2978 7100
rect 3002 7098 3058 7100
rect 3082 7098 3138 7100
rect 3162 7098 3218 7100
rect 2922 7046 2968 7098
rect 2968 7046 2978 7098
rect 3002 7046 3032 7098
rect 3032 7046 3044 7098
rect 3044 7046 3058 7098
rect 3082 7046 3096 7098
rect 3096 7046 3108 7098
rect 3108 7046 3138 7098
rect 3162 7046 3172 7098
rect 3172 7046 3218 7098
rect 2922 7044 2978 7046
rect 3002 7044 3058 7046
rect 3082 7044 3138 7046
rect 3162 7044 3218 7046
rect 2042 3984 2098 4040
rect 2922 6010 2978 6012
rect 3002 6010 3058 6012
rect 3082 6010 3138 6012
rect 3162 6010 3218 6012
rect 2922 5958 2968 6010
rect 2968 5958 2978 6010
rect 3002 5958 3032 6010
rect 3032 5958 3044 6010
rect 3044 5958 3058 6010
rect 3082 5958 3096 6010
rect 3096 5958 3108 6010
rect 3108 5958 3138 6010
rect 3162 5958 3172 6010
rect 3172 5958 3218 6010
rect 2922 5956 2978 5958
rect 3002 5956 3058 5958
rect 3082 5956 3138 5958
rect 3162 5956 3218 5958
rect 4888 13082 4944 13084
rect 4968 13082 5024 13084
rect 5048 13082 5104 13084
rect 5128 13082 5184 13084
rect 4888 13030 4934 13082
rect 4934 13030 4944 13082
rect 4968 13030 4998 13082
rect 4998 13030 5010 13082
rect 5010 13030 5024 13082
rect 5048 13030 5062 13082
rect 5062 13030 5074 13082
rect 5074 13030 5104 13082
rect 5128 13030 5138 13082
rect 5138 13030 5184 13082
rect 4888 13028 4944 13030
rect 4968 13028 5024 13030
rect 5048 13028 5104 13030
rect 5128 13028 5184 13030
rect 3974 9696 4030 9752
rect 4888 11994 4944 11996
rect 4968 11994 5024 11996
rect 5048 11994 5104 11996
rect 5128 11994 5184 11996
rect 4888 11942 4934 11994
rect 4934 11942 4944 11994
rect 4968 11942 4998 11994
rect 4998 11942 5010 11994
rect 5010 11942 5024 11994
rect 5048 11942 5062 11994
rect 5062 11942 5074 11994
rect 5074 11942 5104 11994
rect 5128 11942 5138 11994
rect 5138 11942 5184 11994
rect 4888 11940 4944 11942
rect 4968 11940 5024 11942
rect 5048 11940 5104 11942
rect 5128 11940 5184 11942
rect 2922 4922 2978 4924
rect 3002 4922 3058 4924
rect 3082 4922 3138 4924
rect 3162 4922 3218 4924
rect 2922 4870 2968 4922
rect 2968 4870 2978 4922
rect 3002 4870 3032 4922
rect 3032 4870 3044 4922
rect 3044 4870 3058 4922
rect 3082 4870 3096 4922
rect 3096 4870 3108 4922
rect 3108 4870 3138 4922
rect 3162 4870 3172 4922
rect 3172 4870 3218 4922
rect 2922 4868 2978 4870
rect 3002 4868 3058 4870
rect 3082 4868 3138 4870
rect 3162 4868 3218 4870
rect 2922 3834 2978 3836
rect 3002 3834 3058 3836
rect 3082 3834 3138 3836
rect 3162 3834 3218 3836
rect 2922 3782 2968 3834
rect 2968 3782 2978 3834
rect 3002 3782 3032 3834
rect 3032 3782 3044 3834
rect 3044 3782 3058 3834
rect 3082 3782 3096 3834
rect 3096 3782 3108 3834
rect 3108 3782 3138 3834
rect 3162 3782 3172 3834
rect 3172 3782 3218 3834
rect 2922 3780 2978 3782
rect 3002 3780 3058 3782
rect 3082 3780 3138 3782
rect 3162 3780 3218 3782
rect 4888 10906 4944 10908
rect 4968 10906 5024 10908
rect 5048 10906 5104 10908
rect 5128 10906 5184 10908
rect 4888 10854 4934 10906
rect 4934 10854 4944 10906
rect 4968 10854 4998 10906
rect 4998 10854 5010 10906
rect 5010 10854 5024 10906
rect 5048 10854 5062 10906
rect 5062 10854 5074 10906
rect 5074 10854 5104 10906
rect 5128 10854 5138 10906
rect 5138 10854 5184 10906
rect 4888 10852 4944 10854
rect 4968 10852 5024 10854
rect 5048 10852 5104 10854
rect 5128 10852 5184 10854
rect 4888 9818 4944 9820
rect 4968 9818 5024 9820
rect 5048 9818 5104 9820
rect 5128 9818 5184 9820
rect 4888 9766 4934 9818
rect 4934 9766 4944 9818
rect 4968 9766 4998 9818
rect 4998 9766 5010 9818
rect 5010 9766 5024 9818
rect 5048 9766 5062 9818
rect 5062 9766 5074 9818
rect 5074 9766 5104 9818
rect 5128 9766 5138 9818
rect 5138 9766 5184 9818
rect 4888 9764 4944 9766
rect 4968 9764 5024 9766
rect 5048 9764 5104 9766
rect 5128 9764 5184 9766
rect 4888 8730 4944 8732
rect 4968 8730 5024 8732
rect 5048 8730 5104 8732
rect 5128 8730 5184 8732
rect 4888 8678 4934 8730
rect 4934 8678 4944 8730
rect 4968 8678 4998 8730
rect 4998 8678 5010 8730
rect 5010 8678 5024 8730
rect 5048 8678 5062 8730
rect 5062 8678 5074 8730
rect 5074 8678 5104 8730
rect 5128 8678 5138 8730
rect 5138 8678 5184 8730
rect 4888 8676 4944 8678
rect 4968 8676 5024 8678
rect 5048 8676 5104 8678
rect 5128 8676 5184 8678
rect 4888 7642 4944 7644
rect 4968 7642 5024 7644
rect 5048 7642 5104 7644
rect 5128 7642 5184 7644
rect 4888 7590 4934 7642
rect 4934 7590 4944 7642
rect 4968 7590 4998 7642
rect 4998 7590 5010 7642
rect 5010 7590 5024 7642
rect 5048 7590 5062 7642
rect 5062 7590 5074 7642
rect 5074 7590 5104 7642
rect 5128 7590 5138 7642
rect 5138 7590 5184 7642
rect 4888 7588 4944 7590
rect 4968 7588 5024 7590
rect 5048 7588 5104 7590
rect 5128 7588 5184 7590
rect 5170 7248 5226 7304
rect 4888 6554 4944 6556
rect 4968 6554 5024 6556
rect 5048 6554 5104 6556
rect 5128 6554 5184 6556
rect 4888 6502 4934 6554
rect 4934 6502 4944 6554
rect 4968 6502 4998 6554
rect 4998 6502 5010 6554
rect 5010 6502 5024 6554
rect 5048 6502 5062 6554
rect 5062 6502 5074 6554
rect 5074 6502 5104 6554
rect 5128 6502 5138 6554
rect 5138 6502 5184 6554
rect 4888 6500 4944 6502
rect 4968 6500 5024 6502
rect 5048 6500 5104 6502
rect 5128 6500 5184 6502
rect 4888 5466 4944 5468
rect 4968 5466 5024 5468
rect 5048 5466 5104 5468
rect 5128 5466 5184 5468
rect 4888 5414 4934 5466
rect 4934 5414 4944 5466
rect 4968 5414 4998 5466
rect 4998 5414 5010 5466
rect 5010 5414 5024 5466
rect 5048 5414 5062 5466
rect 5062 5414 5074 5466
rect 5074 5414 5104 5466
rect 5128 5414 5138 5466
rect 5138 5414 5184 5466
rect 4888 5412 4944 5414
rect 4968 5412 5024 5414
rect 5048 5412 5104 5414
rect 5128 5412 5184 5414
rect 6855 14714 6911 14716
rect 6935 14714 6991 14716
rect 7015 14714 7071 14716
rect 7095 14714 7151 14716
rect 6855 14662 6901 14714
rect 6901 14662 6911 14714
rect 6935 14662 6965 14714
rect 6965 14662 6977 14714
rect 6977 14662 6991 14714
rect 7015 14662 7029 14714
rect 7029 14662 7041 14714
rect 7041 14662 7071 14714
rect 7095 14662 7105 14714
rect 7105 14662 7151 14714
rect 6855 14660 6911 14662
rect 6935 14660 6991 14662
rect 7015 14660 7071 14662
rect 7095 14660 7151 14662
rect 8821 15258 8877 15260
rect 8901 15258 8957 15260
rect 8981 15258 9037 15260
rect 9061 15258 9117 15260
rect 8821 15206 8867 15258
rect 8867 15206 8877 15258
rect 8901 15206 8931 15258
rect 8931 15206 8943 15258
rect 8943 15206 8957 15258
rect 8981 15206 8995 15258
rect 8995 15206 9007 15258
rect 9007 15206 9037 15258
rect 9061 15206 9071 15258
rect 9071 15206 9117 15258
rect 8821 15204 8877 15206
rect 8901 15204 8957 15206
rect 8981 15204 9037 15206
rect 9061 15204 9117 15206
rect 10788 14714 10844 14716
rect 10868 14714 10924 14716
rect 10948 14714 11004 14716
rect 11028 14714 11084 14716
rect 10788 14662 10834 14714
rect 10834 14662 10844 14714
rect 10868 14662 10898 14714
rect 10898 14662 10910 14714
rect 10910 14662 10924 14714
rect 10948 14662 10962 14714
rect 10962 14662 10974 14714
rect 10974 14662 11004 14714
rect 11028 14662 11038 14714
rect 11038 14662 11084 14714
rect 10788 14660 10844 14662
rect 10868 14660 10924 14662
rect 10948 14660 11004 14662
rect 11028 14660 11084 14662
rect 8821 14170 8877 14172
rect 8901 14170 8957 14172
rect 8981 14170 9037 14172
rect 9061 14170 9117 14172
rect 8821 14118 8867 14170
rect 8867 14118 8877 14170
rect 8901 14118 8931 14170
rect 8931 14118 8943 14170
rect 8943 14118 8957 14170
rect 8981 14118 8995 14170
rect 8995 14118 9007 14170
rect 9007 14118 9037 14170
rect 9061 14118 9071 14170
rect 9071 14118 9117 14170
rect 8821 14116 8877 14118
rect 8901 14116 8957 14118
rect 8981 14116 9037 14118
rect 9061 14116 9117 14118
rect 10874 14048 10930 14104
rect 6855 13626 6911 13628
rect 6935 13626 6991 13628
rect 7015 13626 7071 13628
rect 7095 13626 7151 13628
rect 6855 13574 6901 13626
rect 6901 13574 6911 13626
rect 6935 13574 6965 13626
rect 6965 13574 6977 13626
rect 6977 13574 6991 13626
rect 7015 13574 7029 13626
rect 7029 13574 7041 13626
rect 7041 13574 7071 13626
rect 7095 13574 7105 13626
rect 7105 13574 7151 13626
rect 6855 13572 6911 13574
rect 6935 13572 6991 13574
rect 7015 13572 7071 13574
rect 7095 13572 7151 13574
rect 6855 12538 6911 12540
rect 6935 12538 6991 12540
rect 7015 12538 7071 12540
rect 7095 12538 7151 12540
rect 6855 12486 6901 12538
rect 6901 12486 6911 12538
rect 6935 12486 6965 12538
rect 6965 12486 6977 12538
rect 6977 12486 6991 12538
rect 7015 12486 7029 12538
rect 7029 12486 7041 12538
rect 7041 12486 7071 12538
rect 7095 12486 7105 12538
rect 7105 12486 7151 12538
rect 6855 12484 6911 12486
rect 6935 12484 6991 12486
rect 7015 12484 7071 12486
rect 7095 12484 7151 12486
rect 6855 11450 6911 11452
rect 6935 11450 6991 11452
rect 7015 11450 7071 11452
rect 7095 11450 7151 11452
rect 6855 11398 6901 11450
rect 6901 11398 6911 11450
rect 6935 11398 6965 11450
rect 6965 11398 6977 11450
rect 6977 11398 6991 11450
rect 7015 11398 7029 11450
rect 7029 11398 7041 11450
rect 7041 11398 7071 11450
rect 7095 11398 7105 11450
rect 7105 11398 7151 11450
rect 6855 11396 6911 11398
rect 6935 11396 6991 11398
rect 7015 11396 7071 11398
rect 7095 11396 7151 11398
rect 6855 10362 6911 10364
rect 6935 10362 6991 10364
rect 7015 10362 7071 10364
rect 7095 10362 7151 10364
rect 6855 10310 6901 10362
rect 6901 10310 6911 10362
rect 6935 10310 6965 10362
rect 6965 10310 6977 10362
rect 6977 10310 6991 10362
rect 7015 10310 7029 10362
rect 7029 10310 7041 10362
rect 7041 10310 7071 10362
rect 7095 10310 7105 10362
rect 7105 10310 7151 10362
rect 6855 10308 6911 10310
rect 6935 10308 6991 10310
rect 7015 10308 7071 10310
rect 7095 10308 7151 10310
rect 6855 9274 6911 9276
rect 6935 9274 6991 9276
rect 7015 9274 7071 9276
rect 7095 9274 7151 9276
rect 6855 9222 6901 9274
rect 6901 9222 6911 9274
rect 6935 9222 6965 9274
rect 6965 9222 6977 9274
rect 6977 9222 6991 9274
rect 7015 9222 7029 9274
rect 7029 9222 7041 9274
rect 7041 9222 7071 9274
rect 7095 9222 7105 9274
rect 7105 9222 7151 9274
rect 6855 9220 6911 9222
rect 6935 9220 6991 9222
rect 7015 9220 7071 9222
rect 7095 9220 7151 9222
rect 6855 8186 6911 8188
rect 6935 8186 6991 8188
rect 7015 8186 7071 8188
rect 7095 8186 7151 8188
rect 6855 8134 6901 8186
rect 6901 8134 6911 8186
rect 6935 8134 6965 8186
rect 6965 8134 6977 8186
rect 6977 8134 6991 8186
rect 7015 8134 7029 8186
rect 7029 8134 7041 8186
rect 7041 8134 7071 8186
rect 7095 8134 7105 8186
rect 7105 8134 7151 8186
rect 6855 8132 6911 8134
rect 6935 8132 6991 8134
rect 7015 8132 7071 8134
rect 7095 8132 7151 8134
rect 6734 7268 6790 7304
rect 6734 7248 6736 7268
rect 6736 7248 6788 7268
rect 6788 7248 6790 7268
rect 6855 7098 6911 7100
rect 6935 7098 6991 7100
rect 7015 7098 7071 7100
rect 7095 7098 7151 7100
rect 6855 7046 6901 7098
rect 6901 7046 6911 7098
rect 6935 7046 6965 7098
rect 6965 7046 6977 7098
rect 6977 7046 6991 7098
rect 7015 7046 7029 7098
rect 7029 7046 7041 7098
rect 7041 7046 7071 7098
rect 7095 7046 7105 7098
rect 7105 7046 7151 7098
rect 6855 7044 6911 7046
rect 6935 7044 6991 7046
rect 7015 7044 7071 7046
rect 7095 7044 7151 7046
rect 6855 6010 6911 6012
rect 6935 6010 6991 6012
rect 7015 6010 7071 6012
rect 7095 6010 7151 6012
rect 6855 5958 6901 6010
rect 6901 5958 6911 6010
rect 6935 5958 6965 6010
rect 6965 5958 6977 6010
rect 6977 5958 6991 6010
rect 7015 5958 7029 6010
rect 7029 5958 7041 6010
rect 7041 5958 7071 6010
rect 7095 5958 7105 6010
rect 7105 5958 7151 6010
rect 6855 5956 6911 5958
rect 6935 5956 6991 5958
rect 7015 5956 7071 5958
rect 7095 5956 7151 5958
rect 8821 13082 8877 13084
rect 8901 13082 8957 13084
rect 8981 13082 9037 13084
rect 9061 13082 9117 13084
rect 8821 13030 8867 13082
rect 8867 13030 8877 13082
rect 8901 13030 8931 13082
rect 8931 13030 8943 13082
rect 8943 13030 8957 13082
rect 8981 13030 8995 13082
rect 8995 13030 9007 13082
rect 9007 13030 9037 13082
rect 9061 13030 9071 13082
rect 9071 13030 9117 13082
rect 8821 13028 8877 13030
rect 8901 13028 8957 13030
rect 8981 13028 9037 13030
rect 9061 13028 9117 13030
rect 8821 11994 8877 11996
rect 8901 11994 8957 11996
rect 8981 11994 9037 11996
rect 9061 11994 9117 11996
rect 8821 11942 8867 11994
rect 8867 11942 8877 11994
rect 8901 11942 8931 11994
rect 8931 11942 8943 11994
rect 8943 11942 8957 11994
rect 8981 11942 8995 11994
rect 8995 11942 9007 11994
rect 9007 11942 9037 11994
rect 9061 11942 9071 11994
rect 9071 11942 9117 11994
rect 8821 11940 8877 11942
rect 8901 11940 8957 11942
rect 8981 11940 9037 11942
rect 9061 11940 9117 11942
rect 8821 10906 8877 10908
rect 8901 10906 8957 10908
rect 8981 10906 9037 10908
rect 9061 10906 9117 10908
rect 8821 10854 8867 10906
rect 8867 10854 8877 10906
rect 8901 10854 8931 10906
rect 8931 10854 8943 10906
rect 8943 10854 8957 10906
rect 8981 10854 8995 10906
rect 8995 10854 9007 10906
rect 9007 10854 9037 10906
rect 9061 10854 9071 10906
rect 9071 10854 9117 10906
rect 8821 10852 8877 10854
rect 8901 10852 8957 10854
rect 8981 10852 9037 10854
rect 9061 10852 9117 10854
rect 6855 4922 6911 4924
rect 6935 4922 6991 4924
rect 7015 4922 7071 4924
rect 7095 4922 7151 4924
rect 6855 4870 6901 4922
rect 6901 4870 6911 4922
rect 6935 4870 6965 4922
rect 6965 4870 6977 4922
rect 6977 4870 6991 4922
rect 7015 4870 7029 4922
rect 7029 4870 7041 4922
rect 7041 4870 7071 4922
rect 7095 4870 7105 4922
rect 7105 4870 7151 4922
rect 6855 4868 6911 4870
rect 6935 4868 6991 4870
rect 7015 4868 7071 4870
rect 7095 4868 7151 4870
rect 4888 4378 4944 4380
rect 4968 4378 5024 4380
rect 5048 4378 5104 4380
rect 5128 4378 5184 4380
rect 4888 4326 4934 4378
rect 4934 4326 4944 4378
rect 4968 4326 4998 4378
rect 4998 4326 5010 4378
rect 5010 4326 5024 4378
rect 5048 4326 5062 4378
rect 5062 4326 5074 4378
rect 5074 4326 5104 4378
rect 5128 4326 5138 4378
rect 5138 4326 5184 4378
rect 4888 4324 4944 4326
rect 4968 4324 5024 4326
rect 5048 4324 5104 4326
rect 5128 4324 5184 4326
rect 8821 9818 8877 9820
rect 8901 9818 8957 9820
rect 8981 9818 9037 9820
rect 9061 9818 9117 9820
rect 8821 9766 8867 9818
rect 8867 9766 8877 9818
rect 8901 9766 8931 9818
rect 8931 9766 8943 9818
rect 8943 9766 8957 9818
rect 8981 9766 8995 9818
rect 8995 9766 9007 9818
rect 9007 9766 9037 9818
rect 9061 9766 9071 9818
rect 9071 9766 9117 9818
rect 8821 9764 8877 9766
rect 8901 9764 8957 9766
rect 8981 9764 9037 9766
rect 9061 9764 9117 9766
rect 8821 8730 8877 8732
rect 8901 8730 8957 8732
rect 8981 8730 9037 8732
rect 9061 8730 9117 8732
rect 8821 8678 8867 8730
rect 8867 8678 8877 8730
rect 8901 8678 8931 8730
rect 8931 8678 8943 8730
rect 8943 8678 8957 8730
rect 8981 8678 8995 8730
rect 8995 8678 9007 8730
rect 9007 8678 9037 8730
rect 9061 8678 9071 8730
rect 9071 8678 9117 8730
rect 8821 8676 8877 8678
rect 8901 8676 8957 8678
rect 8981 8676 9037 8678
rect 9061 8676 9117 8678
rect 8821 7642 8877 7644
rect 8901 7642 8957 7644
rect 8981 7642 9037 7644
rect 9061 7642 9117 7644
rect 8821 7590 8867 7642
rect 8867 7590 8877 7642
rect 8901 7590 8931 7642
rect 8931 7590 8943 7642
rect 8943 7590 8957 7642
rect 8981 7590 8995 7642
rect 8995 7590 9007 7642
rect 9007 7590 9037 7642
rect 9061 7590 9071 7642
rect 9071 7590 9117 7642
rect 8821 7588 8877 7590
rect 8901 7588 8957 7590
rect 8981 7588 9037 7590
rect 9061 7588 9117 7590
rect 8821 6554 8877 6556
rect 8901 6554 8957 6556
rect 8981 6554 9037 6556
rect 9061 6554 9117 6556
rect 8821 6502 8867 6554
rect 8867 6502 8877 6554
rect 8901 6502 8931 6554
rect 8931 6502 8943 6554
rect 8943 6502 8957 6554
rect 8981 6502 8995 6554
rect 8995 6502 9007 6554
rect 9007 6502 9037 6554
rect 9061 6502 9071 6554
rect 9071 6502 9117 6554
rect 8821 6500 8877 6502
rect 8901 6500 8957 6502
rect 8981 6500 9037 6502
rect 9061 6500 9117 6502
rect 10788 13626 10844 13628
rect 10868 13626 10924 13628
rect 10948 13626 11004 13628
rect 11028 13626 11084 13628
rect 10788 13574 10834 13626
rect 10834 13574 10844 13626
rect 10868 13574 10898 13626
rect 10898 13574 10910 13626
rect 10910 13574 10924 13626
rect 10948 13574 10962 13626
rect 10962 13574 10974 13626
rect 10974 13574 11004 13626
rect 11028 13574 11038 13626
rect 11038 13574 11084 13626
rect 10788 13572 10844 13574
rect 10868 13572 10924 13574
rect 10948 13572 11004 13574
rect 11028 13572 11084 13574
rect 11886 14068 11942 14104
rect 11886 14048 11888 14068
rect 11888 14048 11940 14068
rect 11940 14048 11942 14068
rect 10788 12538 10844 12540
rect 10868 12538 10924 12540
rect 10948 12538 11004 12540
rect 11028 12538 11084 12540
rect 10788 12486 10834 12538
rect 10834 12486 10844 12538
rect 10868 12486 10898 12538
rect 10898 12486 10910 12538
rect 10910 12486 10924 12538
rect 10948 12486 10962 12538
rect 10962 12486 10974 12538
rect 10974 12486 11004 12538
rect 11028 12486 11038 12538
rect 11038 12486 11084 12538
rect 10788 12484 10844 12486
rect 10868 12484 10924 12486
rect 10948 12484 11004 12486
rect 11028 12484 11084 12486
rect 12754 15258 12810 15260
rect 12834 15258 12890 15260
rect 12914 15258 12970 15260
rect 12994 15258 13050 15260
rect 12754 15206 12800 15258
rect 12800 15206 12810 15258
rect 12834 15206 12864 15258
rect 12864 15206 12876 15258
rect 12876 15206 12890 15258
rect 12914 15206 12928 15258
rect 12928 15206 12940 15258
rect 12940 15206 12970 15258
rect 12994 15206 13004 15258
rect 13004 15206 13050 15258
rect 12754 15204 12810 15206
rect 12834 15204 12890 15206
rect 12914 15204 12970 15206
rect 12994 15204 13050 15206
rect 10788 11450 10844 11452
rect 10868 11450 10924 11452
rect 10948 11450 11004 11452
rect 11028 11450 11084 11452
rect 10788 11398 10834 11450
rect 10834 11398 10844 11450
rect 10868 11398 10898 11450
rect 10898 11398 10910 11450
rect 10910 11398 10924 11450
rect 10948 11398 10962 11450
rect 10962 11398 10974 11450
rect 10974 11398 11004 11450
rect 11028 11398 11038 11450
rect 11038 11398 11084 11450
rect 10788 11396 10844 11398
rect 10868 11396 10924 11398
rect 10948 11396 11004 11398
rect 11028 11396 11084 11398
rect 10788 10362 10844 10364
rect 10868 10362 10924 10364
rect 10948 10362 11004 10364
rect 11028 10362 11084 10364
rect 10788 10310 10834 10362
rect 10834 10310 10844 10362
rect 10868 10310 10898 10362
rect 10898 10310 10910 10362
rect 10910 10310 10924 10362
rect 10948 10310 10962 10362
rect 10962 10310 10974 10362
rect 10974 10310 11004 10362
rect 11028 10310 11038 10362
rect 11038 10310 11084 10362
rect 10788 10308 10844 10310
rect 10868 10308 10924 10310
rect 10948 10308 11004 10310
rect 11028 10308 11084 10310
rect 10788 9274 10844 9276
rect 10868 9274 10924 9276
rect 10948 9274 11004 9276
rect 11028 9274 11084 9276
rect 10788 9222 10834 9274
rect 10834 9222 10844 9274
rect 10868 9222 10898 9274
rect 10898 9222 10910 9274
rect 10910 9222 10924 9274
rect 10948 9222 10962 9274
rect 10962 9222 10974 9274
rect 10974 9222 11004 9274
rect 11028 9222 11038 9274
rect 11038 9222 11084 9274
rect 10788 9220 10844 9222
rect 10868 9220 10924 9222
rect 10948 9220 11004 9222
rect 11028 9220 11084 9222
rect 12754 14170 12810 14172
rect 12834 14170 12890 14172
rect 12914 14170 12970 14172
rect 12994 14170 13050 14172
rect 12754 14118 12800 14170
rect 12800 14118 12810 14170
rect 12834 14118 12864 14170
rect 12864 14118 12876 14170
rect 12876 14118 12890 14170
rect 12914 14118 12928 14170
rect 12928 14118 12940 14170
rect 12940 14118 12970 14170
rect 12994 14118 13004 14170
rect 13004 14118 13050 14170
rect 12754 14116 12810 14118
rect 12834 14116 12890 14118
rect 12914 14116 12970 14118
rect 12994 14116 13050 14118
rect 12754 13082 12810 13084
rect 12834 13082 12890 13084
rect 12914 13082 12970 13084
rect 12994 13082 13050 13084
rect 12754 13030 12800 13082
rect 12800 13030 12810 13082
rect 12834 13030 12864 13082
rect 12864 13030 12876 13082
rect 12876 13030 12890 13082
rect 12914 13030 12928 13082
rect 12928 13030 12940 13082
rect 12940 13030 12970 13082
rect 12994 13030 13004 13082
rect 13004 13030 13050 13082
rect 12754 13028 12810 13030
rect 12834 13028 12890 13030
rect 12914 13028 12970 13030
rect 12994 13028 13050 13030
rect 14721 15802 14777 15804
rect 14801 15802 14857 15804
rect 14881 15802 14937 15804
rect 14961 15802 15017 15804
rect 14721 15750 14767 15802
rect 14767 15750 14777 15802
rect 14801 15750 14831 15802
rect 14831 15750 14843 15802
rect 14843 15750 14857 15802
rect 14881 15750 14895 15802
rect 14895 15750 14907 15802
rect 14907 15750 14937 15802
rect 14961 15750 14971 15802
rect 14971 15750 15017 15802
rect 14721 15748 14777 15750
rect 14801 15748 14857 15750
rect 14881 15748 14937 15750
rect 14961 15748 15017 15750
rect 12754 11994 12810 11996
rect 12834 11994 12890 11996
rect 12914 11994 12970 11996
rect 12994 11994 13050 11996
rect 12754 11942 12800 11994
rect 12800 11942 12810 11994
rect 12834 11942 12864 11994
rect 12864 11942 12876 11994
rect 12876 11942 12890 11994
rect 12914 11942 12928 11994
rect 12928 11942 12940 11994
rect 12940 11942 12970 11994
rect 12994 11942 13004 11994
rect 13004 11942 13050 11994
rect 12754 11940 12810 11942
rect 12834 11940 12890 11942
rect 12914 11940 12970 11942
rect 12994 11940 13050 11942
rect 12754 10906 12810 10908
rect 12834 10906 12890 10908
rect 12914 10906 12970 10908
rect 12994 10906 13050 10908
rect 12754 10854 12800 10906
rect 12800 10854 12810 10906
rect 12834 10854 12864 10906
rect 12864 10854 12876 10906
rect 12876 10854 12890 10906
rect 12914 10854 12928 10906
rect 12928 10854 12940 10906
rect 12940 10854 12970 10906
rect 12994 10854 13004 10906
rect 13004 10854 13050 10906
rect 12754 10852 12810 10854
rect 12834 10852 12890 10854
rect 12914 10852 12970 10854
rect 12994 10852 13050 10854
rect 16687 15258 16743 15260
rect 16767 15258 16823 15260
rect 16847 15258 16903 15260
rect 16927 15258 16983 15260
rect 16687 15206 16733 15258
rect 16733 15206 16743 15258
rect 16767 15206 16797 15258
rect 16797 15206 16809 15258
rect 16809 15206 16823 15258
rect 16847 15206 16861 15258
rect 16861 15206 16873 15258
rect 16873 15206 16903 15258
rect 16927 15206 16937 15258
rect 16937 15206 16983 15258
rect 16687 15204 16743 15206
rect 16767 15204 16823 15206
rect 16847 15204 16903 15206
rect 16927 15204 16983 15206
rect 14721 14714 14777 14716
rect 14801 14714 14857 14716
rect 14881 14714 14937 14716
rect 14961 14714 15017 14716
rect 14721 14662 14767 14714
rect 14767 14662 14777 14714
rect 14801 14662 14831 14714
rect 14831 14662 14843 14714
rect 14843 14662 14857 14714
rect 14881 14662 14895 14714
rect 14895 14662 14907 14714
rect 14907 14662 14937 14714
rect 14961 14662 14971 14714
rect 14971 14662 15017 14714
rect 14721 14660 14777 14662
rect 14801 14660 14857 14662
rect 14881 14660 14937 14662
rect 14961 14660 15017 14662
rect 14094 13912 14150 13968
rect 14721 13626 14777 13628
rect 14801 13626 14857 13628
rect 14881 13626 14937 13628
rect 14961 13626 15017 13628
rect 14721 13574 14767 13626
rect 14767 13574 14777 13626
rect 14801 13574 14831 13626
rect 14831 13574 14843 13626
rect 14843 13574 14857 13626
rect 14881 13574 14895 13626
rect 14895 13574 14907 13626
rect 14907 13574 14937 13626
rect 14961 13574 14971 13626
rect 14971 13574 15017 13626
rect 14721 13572 14777 13574
rect 14801 13572 14857 13574
rect 14881 13572 14937 13574
rect 14961 13572 15017 13574
rect 14721 12538 14777 12540
rect 14801 12538 14857 12540
rect 14881 12538 14937 12540
rect 14961 12538 15017 12540
rect 14721 12486 14767 12538
rect 14767 12486 14777 12538
rect 14801 12486 14831 12538
rect 14831 12486 14843 12538
rect 14843 12486 14857 12538
rect 14881 12486 14895 12538
rect 14895 12486 14907 12538
rect 14907 12486 14937 12538
rect 14961 12486 14971 12538
rect 14971 12486 15017 12538
rect 14721 12484 14777 12486
rect 14801 12484 14857 12486
rect 14881 12484 14937 12486
rect 14961 12484 15017 12486
rect 16687 14170 16743 14172
rect 16767 14170 16823 14172
rect 16847 14170 16903 14172
rect 16927 14170 16983 14172
rect 16687 14118 16733 14170
rect 16733 14118 16743 14170
rect 16767 14118 16797 14170
rect 16797 14118 16809 14170
rect 16809 14118 16823 14170
rect 16847 14118 16861 14170
rect 16861 14118 16873 14170
rect 16873 14118 16903 14170
rect 16927 14118 16937 14170
rect 16937 14118 16983 14170
rect 16687 14116 16743 14118
rect 16767 14116 16823 14118
rect 16847 14116 16903 14118
rect 16927 14116 16983 14118
rect 16687 13082 16743 13084
rect 16767 13082 16823 13084
rect 16847 13082 16903 13084
rect 16927 13082 16983 13084
rect 16687 13030 16733 13082
rect 16733 13030 16743 13082
rect 16767 13030 16797 13082
rect 16797 13030 16809 13082
rect 16809 13030 16823 13082
rect 16847 13030 16861 13082
rect 16861 13030 16873 13082
rect 16873 13030 16903 13082
rect 16927 13030 16937 13082
rect 16937 13030 16983 13082
rect 16687 13028 16743 13030
rect 16767 13028 16823 13030
rect 16847 13028 16903 13030
rect 16927 13028 16983 13030
rect 14721 11450 14777 11452
rect 14801 11450 14857 11452
rect 14881 11450 14937 11452
rect 14961 11450 15017 11452
rect 14721 11398 14767 11450
rect 14767 11398 14777 11450
rect 14801 11398 14831 11450
rect 14831 11398 14843 11450
rect 14843 11398 14857 11450
rect 14881 11398 14895 11450
rect 14895 11398 14907 11450
rect 14907 11398 14937 11450
rect 14961 11398 14971 11450
rect 14971 11398 15017 11450
rect 14721 11396 14777 11398
rect 14801 11396 14857 11398
rect 14881 11396 14937 11398
rect 14961 11396 15017 11398
rect 14721 10362 14777 10364
rect 14801 10362 14857 10364
rect 14881 10362 14937 10364
rect 14961 10362 15017 10364
rect 14721 10310 14767 10362
rect 14767 10310 14777 10362
rect 14801 10310 14831 10362
rect 14831 10310 14843 10362
rect 14843 10310 14857 10362
rect 14881 10310 14895 10362
rect 14895 10310 14907 10362
rect 14907 10310 14937 10362
rect 14961 10310 14971 10362
rect 14971 10310 15017 10362
rect 14721 10308 14777 10310
rect 14801 10308 14857 10310
rect 14881 10308 14937 10310
rect 14961 10308 15017 10310
rect 16687 11994 16743 11996
rect 16767 11994 16823 11996
rect 16847 11994 16903 11996
rect 16927 11994 16983 11996
rect 16687 11942 16733 11994
rect 16733 11942 16743 11994
rect 16767 11942 16797 11994
rect 16797 11942 16809 11994
rect 16809 11942 16823 11994
rect 16847 11942 16861 11994
rect 16861 11942 16873 11994
rect 16873 11942 16903 11994
rect 16927 11942 16937 11994
rect 16937 11942 16983 11994
rect 16687 11940 16743 11942
rect 16767 11940 16823 11942
rect 16847 11940 16903 11942
rect 16927 11940 16983 11942
rect 16687 10906 16743 10908
rect 16767 10906 16823 10908
rect 16847 10906 16903 10908
rect 16927 10906 16983 10908
rect 16687 10854 16733 10906
rect 16733 10854 16743 10906
rect 16767 10854 16797 10906
rect 16797 10854 16809 10906
rect 16809 10854 16823 10906
rect 16847 10854 16861 10906
rect 16861 10854 16873 10906
rect 16873 10854 16903 10906
rect 16927 10854 16937 10906
rect 16937 10854 16983 10906
rect 16687 10852 16743 10854
rect 16767 10852 16823 10854
rect 16847 10852 16903 10854
rect 16927 10852 16983 10854
rect 12754 9818 12810 9820
rect 12834 9818 12890 9820
rect 12914 9818 12970 9820
rect 12994 9818 13050 9820
rect 12754 9766 12800 9818
rect 12800 9766 12810 9818
rect 12834 9766 12864 9818
rect 12864 9766 12876 9818
rect 12876 9766 12890 9818
rect 12914 9766 12928 9818
rect 12928 9766 12940 9818
rect 12940 9766 12970 9818
rect 12994 9766 13004 9818
rect 13004 9766 13050 9818
rect 12754 9764 12810 9766
rect 12834 9764 12890 9766
rect 12914 9764 12970 9766
rect 12994 9764 13050 9766
rect 14721 9274 14777 9276
rect 14801 9274 14857 9276
rect 14881 9274 14937 9276
rect 14961 9274 15017 9276
rect 14721 9222 14767 9274
rect 14767 9222 14777 9274
rect 14801 9222 14831 9274
rect 14831 9222 14843 9274
rect 14843 9222 14857 9274
rect 14881 9222 14895 9274
rect 14895 9222 14907 9274
rect 14907 9222 14937 9274
rect 14961 9222 14971 9274
rect 14971 9222 15017 9274
rect 14721 9220 14777 9222
rect 14801 9220 14857 9222
rect 14881 9220 14937 9222
rect 14961 9220 15017 9222
rect 8821 5466 8877 5468
rect 8901 5466 8957 5468
rect 8981 5466 9037 5468
rect 9061 5466 9117 5468
rect 8821 5414 8867 5466
rect 8867 5414 8877 5466
rect 8901 5414 8931 5466
rect 8931 5414 8943 5466
rect 8943 5414 8957 5466
rect 8981 5414 8995 5466
rect 8995 5414 9007 5466
rect 9007 5414 9037 5466
rect 9061 5414 9071 5466
rect 9071 5414 9117 5466
rect 8821 5412 8877 5414
rect 8901 5412 8957 5414
rect 8981 5412 9037 5414
rect 9061 5412 9117 5414
rect 10788 8186 10844 8188
rect 10868 8186 10924 8188
rect 10948 8186 11004 8188
rect 11028 8186 11084 8188
rect 10788 8134 10834 8186
rect 10834 8134 10844 8186
rect 10868 8134 10898 8186
rect 10898 8134 10910 8186
rect 10910 8134 10924 8186
rect 10948 8134 10962 8186
rect 10962 8134 10974 8186
rect 10974 8134 11004 8186
rect 11028 8134 11038 8186
rect 11038 8134 11084 8186
rect 10788 8132 10844 8134
rect 10868 8132 10924 8134
rect 10948 8132 11004 8134
rect 11028 8132 11084 8134
rect 10788 7098 10844 7100
rect 10868 7098 10924 7100
rect 10948 7098 11004 7100
rect 11028 7098 11084 7100
rect 10788 7046 10834 7098
rect 10834 7046 10844 7098
rect 10868 7046 10898 7098
rect 10898 7046 10910 7098
rect 10910 7046 10924 7098
rect 10948 7046 10962 7098
rect 10962 7046 10974 7098
rect 10974 7046 11004 7098
rect 11028 7046 11038 7098
rect 11038 7046 11084 7098
rect 10788 7044 10844 7046
rect 10868 7044 10924 7046
rect 10948 7044 11004 7046
rect 11028 7044 11084 7046
rect 10788 6010 10844 6012
rect 10868 6010 10924 6012
rect 10948 6010 11004 6012
rect 11028 6010 11084 6012
rect 10788 5958 10834 6010
rect 10834 5958 10844 6010
rect 10868 5958 10898 6010
rect 10898 5958 10910 6010
rect 10910 5958 10924 6010
rect 10948 5958 10962 6010
rect 10962 5958 10974 6010
rect 10974 5958 11004 6010
rect 11028 5958 11038 6010
rect 11038 5958 11084 6010
rect 10788 5956 10844 5958
rect 10868 5956 10924 5958
rect 10948 5956 11004 5958
rect 11028 5956 11084 5958
rect 12754 8730 12810 8732
rect 12834 8730 12890 8732
rect 12914 8730 12970 8732
rect 12994 8730 13050 8732
rect 12754 8678 12800 8730
rect 12800 8678 12810 8730
rect 12834 8678 12864 8730
rect 12864 8678 12876 8730
rect 12876 8678 12890 8730
rect 12914 8678 12928 8730
rect 12928 8678 12940 8730
rect 12940 8678 12970 8730
rect 12994 8678 13004 8730
rect 13004 8678 13050 8730
rect 12754 8676 12810 8678
rect 12834 8676 12890 8678
rect 12914 8676 12970 8678
rect 12994 8676 13050 8678
rect 12754 7642 12810 7644
rect 12834 7642 12890 7644
rect 12914 7642 12970 7644
rect 12994 7642 13050 7644
rect 12754 7590 12800 7642
rect 12800 7590 12810 7642
rect 12834 7590 12864 7642
rect 12864 7590 12876 7642
rect 12876 7590 12890 7642
rect 12914 7590 12928 7642
rect 12928 7590 12940 7642
rect 12940 7590 12970 7642
rect 12994 7590 13004 7642
rect 13004 7590 13050 7642
rect 12754 7588 12810 7590
rect 12834 7588 12890 7590
rect 12914 7588 12970 7590
rect 12994 7588 13050 7590
rect 16687 9818 16743 9820
rect 16767 9818 16823 9820
rect 16847 9818 16903 9820
rect 16927 9818 16983 9820
rect 16687 9766 16733 9818
rect 16733 9766 16743 9818
rect 16767 9766 16797 9818
rect 16797 9766 16809 9818
rect 16809 9766 16823 9818
rect 16847 9766 16861 9818
rect 16861 9766 16873 9818
rect 16873 9766 16903 9818
rect 16927 9766 16937 9818
rect 16937 9766 16983 9818
rect 16687 9764 16743 9766
rect 16767 9764 16823 9766
rect 16847 9764 16903 9766
rect 16927 9764 16983 9766
rect 16687 8730 16743 8732
rect 16767 8730 16823 8732
rect 16847 8730 16903 8732
rect 16927 8730 16983 8732
rect 16687 8678 16733 8730
rect 16733 8678 16743 8730
rect 16767 8678 16797 8730
rect 16797 8678 16809 8730
rect 16809 8678 16823 8730
rect 16847 8678 16861 8730
rect 16861 8678 16873 8730
rect 16873 8678 16903 8730
rect 16927 8678 16937 8730
rect 16937 8678 16983 8730
rect 16687 8676 16743 8678
rect 16767 8676 16823 8678
rect 16847 8676 16903 8678
rect 16927 8676 16983 8678
rect 14721 8186 14777 8188
rect 14801 8186 14857 8188
rect 14881 8186 14937 8188
rect 14961 8186 15017 8188
rect 14721 8134 14767 8186
rect 14767 8134 14777 8186
rect 14801 8134 14831 8186
rect 14831 8134 14843 8186
rect 14843 8134 14857 8186
rect 14881 8134 14895 8186
rect 14895 8134 14907 8186
rect 14907 8134 14937 8186
rect 14961 8134 14971 8186
rect 14971 8134 15017 8186
rect 14721 8132 14777 8134
rect 14801 8132 14857 8134
rect 14881 8132 14937 8134
rect 14961 8132 15017 8134
rect 16687 7642 16743 7644
rect 16767 7642 16823 7644
rect 16847 7642 16903 7644
rect 16927 7642 16983 7644
rect 16687 7590 16733 7642
rect 16733 7590 16743 7642
rect 16767 7590 16797 7642
rect 16797 7590 16809 7642
rect 16809 7590 16823 7642
rect 16847 7590 16861 7642
rect 16861 7590 16873 7642
rect 16873 7590 16903 7642
rect 16927 7590 16937 7642
rect 16937 7590 16983 7642
rect 16687 7588 16743 7590
rect 16767 7588 16823 7590
rect 16847 7588 16903 7590
rect 16927 7588 16983 7590
rect 14721 7098 14777 7100
rect 14801 7098 14857 7100
rect 14881 7098 14937 7100
rect 14961 7098 15017 7100
rect 14721 7046 14767 7098
rect 14767 7046 14777 7098
rect 14801 7046 14831 7098
rect 14831 7046 14843 7098
rect 14843 7046 14857 7098
rect 14881 7046 14895 7098
rect 14895 7046 14907 7098
rect 14907 7046 14937 7098
rect 14961 7046 14971 7098
rect 14971 7046 15017 7098
rect 14721 7044 14777 7046
rect 14801 7044 14857 7046
rect 14881 7044 14937 7046
rect 14961 7044 15017 7046
rect 12754 6554 12810 6556
rect 12834 6554 12890 6556
rect 12914 6554 12970 6556
rect 12994 6554 13050 6556
rect 12754 6502 12800 6554
rect 12800 6502 12810 6554
rect 12834 6502 12864 6554
rect 12864 6502 12876 6554
rect 12876 6502 12890 6554
rect 12914 6502 12928 6554
rect 12928 6502 12940 6554
rect 12940 6502 12970 6554
rect 12994 6502 13004 6554
rect 13004 6502 13050 6554
rect 12754 6500 12810 6502
rect 12834 6500 12890 6502
rect 12914 6500 12970 6502
rect 12994 6500 13050 6502
rect 16687 6554 16743 6556
rect 16767 6554 16823 6556
rect 16847 6554 16903 6556
rect 16927 6554 16983 6556
rect 16687 6502 16733 6554
rect 16733 6502 16743 6554
rect 16767 6502 16797 6554
rect 16797 6502 16809 6554
rect 16809 6502 16823 6554
rect 16847 6502 16861 6554
rect 16861 6502 16873 6554
rect 16873 6502 16903 6554
rect 16927 6502 16937 6554
rect 16937 6502 16983 6554
rect 16687 6500 16743 6502
rect 16767 6500 16823 6502
rect 16847 6500 16903 6502
rect 16927 6500 16983 6502
rect 14721 6010 14777 6012
rect 14801 6010 14857 6012
rect 14881 6010 14937 6012
rect 14961 6010 15017 6012
rect 14721 5958 14767 6010
rect 14767 5958 14777 6010
rect 14801 5958 14831 6010
rect 14831 5958 14843 6010
rect 14843 5958 14857 6010
rect 14881 5958 14895 6010
rect 14895 5958 14907 6010
rect 14907 5958 14937 6010
rect 14961 5958 14971 6010
rect 14971 5958 15017 6010
rect 14721 5956 14777 5958
rect 14801 5956 14857 5958
rect 14881 5956 14937 5958
rect 14961 5956 15017 5958
rect 10788 4922 10844 4924
rect 10868 4922 10924 4924
rect 10948 4922 11004 4924
rect 11028 4922 11084 4924
rect 10788 4870 10834 4922
rect 10834 4870 10844 4922
rect 10868 4870 10898 4922
rect 10898 4870 10910 4922
rect 10910 4870 10924 4922
rect 10948 4870 10962 4922
rect 10962 4870 10974 4922
rect 10974 4870 11004 4922
rect 11028 4870 11038 4922
rect 11038 4870 11084 4922
rect 10788 4868 10844 4870
rect 10868 4868 10924 4870
rect 10948 4868 11004 4870
rect 11028 4868 11084 4870
rect 12754 5466 12810 5468
rect 12834 5466 12890 5468
rect 12914 5466 12970 5468
rect 12994 5466 13050 5468
rect 12754 5414 12800 5466
rect 12800 5414 12810 5466
rect 12834 5414 12864 5466
rect 12864 5414 12876 5466
rect 12876 5414 12890 5466
rect 12914 5414 12928 5466
rect 12928 5414 12940 5466
rect 12940 5414 12970 5466
rect 12994 5414 13004 5466
rect 13004 5414 13050 5466
rect 12754 5412 12810 5414
rect 12834 5412 12890 5414
rect 12914 5412 12970 5414
rect 12994 5412 13050 5414
rect 16687 5466 16743 5468
rect 16767 5466 16823 5468
rect 16847 5466 16903 5468
rect 16927 5466 16983 5468
rect 16687 5414 16733 5466
rect 16733 5414 16743 5466
rect 16767 5414 16797 5466
rect 16797 5414 16809 5466
rect 16809 5414 16823 5466
rect 16847 5414 16861 5466
rect 16861 5414 16873 5466
rect 16873 5414 16903 5466
rect 16927 5414 16937 5466
rect 16937 5414 16983 5466
rect 16687 5412 16743 5414
rect 16767 5412 16823 5414
rect 16847 5412 16903 5414
rect 16927 5412 16983 5414
rect 14721 4922 14777 4924
rect 14801 4922 14857 4924
rect 14881 4922 14937 4924
rect 14961 4922 15017 4924
rect 14721 4870 14767 4922
rect 14767 4870 14777 4922
rect 14801 4870 14831 4922
rect 14831 4870 14843 4922
rect 14843 4870 14857 4922
rect 14881 4870 14895 4922
rect 14895 4870 14907 4922
rect 14907 4870 14937 4922
rect 14961 4870 14971 4922
rect 14971 4870 15017 4922
rect 14721 4868 14777 4870
rect 14801 4868 14857 4870
rect 14881 4868 14937 4870
rect 14961 4868 15017 4870
rect 8821 4378 8877 4380
rect 8901 4378 8957 4380
rect 8981 4378 9037 4380
rect 9061 4378 9117 4380
rect 8821 4326 8867 4378
rect 8867 4326 8877 4378
rect 8901 4326 8931 4378
rect 8931 4326 8943 4378
rect 8943 4326 8957 4378
rect 8981 4326 8995 4378
rect 8995 4326 9007 4378
rect 9007 4326 9037 4378
rect 9061 4326 9071 4378
rect 9071 4326 9117 4378
rect 8821 4324 8877 4326
rect 8901 4324 8957 4326
rect 8981 4324 9037 4326
rect 9061 4324 9117 4326
rect 12754 4378 12810 4380
rect 12834 4378 12890 4380
rect 12914 4378 12970 4380
rect 12994 4378 13050 4380
rect 12754 4326 12800 4378
rect 12800 4326 12810 4378
rect 12834 4326 12864 4378
rect 12864 4326 12876 4378
rect 12876 4326 12890 4378
rect 12914 4326 12928 4378
rect 12928 4326 12940 4378
rect 12940 4326 12970 4378
rect 12994 4326 13004 4378
rect 13004 4326 13050 4378
rect 12754 4324 12810 4326
rect 12834 4324 12890 4326
rect 12914 4324 12970 4326
rect 12994 4324 13050 4326
rect 16687 4378 16743 4380
rect 16767 4378 16823 4380
rect 16847 4378 16903 4380
rect 16927 4378 16983 4380
rect 16687 4326 16733 4378
rect 16733 4326 16743 4378
rect 16767 4326 16797 4378
rect 16797 4326 16809 4378
rect 16809 4326 16823 4378
rect 16847 4326 16861 4378
rect 16861 4326 16873 4378
rect 16873 4326 16903 4378
rect 16927 4326 16937 4378
rect 16937 4326 16983 4378
rect 16687 4324 16743 4326
rect 16767 4324 16823 4326
rect 16847 4324 16903 4326
rect 16927 4324 16983 4326
rect 6855 3834 6911 3836
rect 6935 3834 6991 3836
rect 7015 3834 7071 3836
rect 7095 3834 7151 3836
rect 6855 3782 6901 3834
rect 6901 3782 6911 3834
rect 6935 3782 6965 3834
rect 6965 3782 6977 3834
rect 6977 3782 6991 3834
rect 7015 3782 7029 3834
rect 7029 3782 7041 3834
rect 7041 3782 7071 3834
rect 7095 3782 7105 3834
rect 7105 3782 7151 3834
rect 6855 3780 6911 3782
rect 6935 3780 6991 3782
rect 7015 3780 7071 3782
rect 7095 3780 7151 3782
rect 10788 3834 10844 3836
rect 10868 3834 10924 3836
rect 10948 3834 11004 3836
rect 11028 3834 11084 3836
rect 10788 3782 10834 3834
rect 10834 3782 10844 3834
rect 10868 3782 10898 3834
rect 10898 3782 10910 3834
rect 10910 3782 10924 3834
rect 10948 3782 10962 3834
rect 10962 3782 10974 3834
rect 10974 3782 11004 3834
rect 11028 3782 11038 3834
rect 11038 3782 11084 3834
rect 10788 3780 10844 3782
rect 10868 3780 10924 3782
rect 10948 3780 11004 3782
rect 11028 3780 11084 3782
rect 14721 3834 14777 3836
rect 14801 3834 14857 3836
rect 14881 3834 14937 3836
rect 14961 3834 15017 3836
rect 14721 3782 14767 3834
rect 14767 3782 14777 3834
rect 14801 3782 14831 3834
rect 14831 3782 14843 3834
rect 14843 3782 14857 3834
rect 14881 3782 14895 3834
rect 14895 3782 14907 3834
rect 14907 3782 14937 3834
rect 14961 3782 14971 3834
rect 14971 3782 15017 3834
rect 14721 3780 14777 3782
rect 14801 3780 14857 3782
rect 14881 3780 14937 3782
rect 14961 3780 15017 3782
rect 4888 3290 4944 3292
rect 4968 3290 5024 3292
rect 5048 3290 5104 3292
rect 5128 3290 5184 3292
rect 4888 3238 4934 3290
rect 4934 3238 4944 3290
rect 4968 3238 4998 3290
rect 4998 3238 5010 3290
rect 5010 3238 5024 3290
rect 5048 3238 5062 3290
rect 5062 3238 5074 3290
rect 5074 3238 5104 3290
rect 5128 3238 5138 3290
rect 5138 3238 5184 3290
rect 4888 3236 4944 3238
rect 4968 3236 5024 3238
rect 5048 3236 5104 3238
rect 5128 3236 5184 3238
rect 8821 3290 8877 3292
rect 8901 3290 8957 3292
rect 8981 3290 9037 3292
rect 9061 3290 9117 3292
rect 8821 3238 8867 3290
rect 8867 3238 8877 3290
rect 8901 3238 8931 3290
rect 8931 3238 8943 3290
rect 8943 3238 8957 3290
rect 8981 3238 8995 3290
rect 8995 3238 9007 3290
rect 9007 3238 9037 3290
rect 9061 3238 9071 3290
rect 9071 3238 9117 3290
rect 8821 3236 8877 3238
rect 8901 3236 8957 3238
rect 8981 3236 9037 3238
rect 9061 3236 9117 3238
rect 12754 3290 12810 3292
rect 12834 3290 12890 3292
rect 12914 3290 12970 3292
rect 12994 3290 13050 3292
rect 12754 3238 12800 3290
rect 12800 3238 12810 3290
rect 12834 3238 12864 3290
rect 12864 3238 12876 3290
rect 12876 3238 12890 3290
rect 12914 3238 12928 3290
rect 12928 3238 12940 3290
rect 12940 3238 12970 3290
rect 12994 3238 13004 3290
rect 13004 3238 13050 3290
rect 12754 3236 12810 3238
rect 12834 3236 12890 3238
rect 12914 3236 12970 3238
rect 12994 3236 13050 3238
rect 16687 3290 16743 3292
rect 16767 3290 16823 3292
rect 16847 3290 16903 3292
rect 16927 3290 16983 3292
rect 16687 3238 16733 3290
rect 16733 3238 16743 3290
rect 16767 3238 16797 3290
rect 16797 3238 16809 3290
rect 16809 3238 16823 3290
rect 16847 3238 16861 3290
rect 16861 3238 16873 3290
rect 16873 3238 16903 3290
rect 16927 3238 16937 3290
rect 16937 3238 16983 3290
rect 16687 3236 16743 3238
rect 16767 3236 16823 3238
rect 16847 3236 16903 3238
rect 16927 3236 16983 3238
rect 2922 2746 2978 2748
rect 3002 2746 3058 2748
rect 3082 2746 3138 2748
rect 3162 2746 3218 2748
rect 2922 2694 2968 2746
rect 2968 2694 2978 2746
rect 3002 2694 3032 2746
rect 3032 2694 3044 2746
rect 3044 2694 3058 2746
rect 3082 2694 3096 2746
rect 3096 2694 3108 2746
rect 3108 2694 3138 2746
rect 3162 2694 3172 2746
rect 3172 2694 3218 2746
rect 2922 2692 2978 2694
rect 3002 2692 3058 2694
rect 3082 2692 3138 2694
rect 3162 2692 3218 2694
rect 6855 2746 6911 2748
rect 6935 2746 6991 2748
rect 7015 2746 7071 2748
rect 7095 2746 7151 2748
rect 6855 2694 6901 2746
rect 6901 2694 6911 2746
rect 6935 2694 6965 2746
rect 6965 2694 6977 2746
rect 6977 2694 6991 2746
rect 7015 2694 7029 2746
rect 7029 2694 7041 2746
rect 7041 2694 7071 2746
rect 7095 2694 7105 2746
rect 7105 2694 7151 2746
rect 6855 2692 6911 2694
rect 6935 2692 6991 2694
rect 7015 2692 7071 2694
rect 7095 2692 7151 2694
rect 10788 2746 10844 2748
rect 10868 2746 10924 2748
rect 10948 2746 11004 2748
rect 11028 2746 11084 2748
rect 10788 2694 10834 2746
rect 10834 2694 10844 2746
rect 10868 2694 10898 2746
rect 10898 2694 10910 2746
rect 10910 2694 10924 2746
rect 10948 2694 10962 2746
rect 10962 2694 10974 2746
rect 10974 2694 11004 2746
rect 11028 2694 11038 2746
rect 11038 2694 11084 2746
rect 10788 2692 10844 2694
rect 10868 2692 10924 2694
rect 10948 2692 11004 2694
rect 11028 2692 11084 2694
rect 14721 2746 14777 2748
rect 14801 2746 14857 2748
rect 14881 2746 14937 2748
rect 14961 2746 15017 2748
rect 14721 2694 14767 2746
rect 14767 2694 14777 2746
rect 14801 2694 14831 2746
rect 14831 2694 14843 2746
rect 14843 2694 14857 2746
rect 14881 2694 14895 2746
rect 14895 2694 14907 2746
rect 14907 2694 14937 2746
rect 14961 2694 14971 2746
rect 14971 2694 15017 2746
rect 14721 2692 14777 2694
rect 14801 2692 14857 2694
rect 14881 2692 14937 2694
rect 14961 2692 15017 2694
rect 1766 2252 1768 2272
rect 1768 2252 1820 2272
rect 1820 2252 1822 2272
rect 1766 2216 1822 2252
rect 4888 2202 4944 2204
rect 4968 2202 5024 2204
rect 5048 2202 5104 2204
rect 5128 2202 5184 2204
rect 4888 2150 4934 2202
rect 4934 2150 4944 2202
rect 4968 2150 4998 2202
rect 4998 2150 5010 2202
rect 5010 2150 5024 2202
rect 5048 2150 5062 2202
rect 5062 2150 5074 2202
rect 5074 2150 5104 2202
rect 5128 2150 5138 2202
rect 5138 2150 5184 2202
rect 4888 2148 4944 2150
rect 4968 2148 5024 2150
rect 5048 2148 5104 2150
rect 5128 2148 5184 2150
rect 8821 2202 8877 2204
rect 8901 2202 8957 2204
rect 8981 2202 9037 2204
rect 9061 2202 9117 2204
rect 8821 2150 8867 2202
rect 8867 2150 8877 2202
rect 8901 2150 8931 2202
rect 8931 2150 8943 2202
rect 8943 2150 8957 2202
rect 8981 2150 8995 2202
rect 8995 2150 9007 2202
rect 9007 2150 9037 2202
rect 9061 2150 9071 2202
rect 9071 2150 9117 2202
rect 8821 2148 8877 2150
rect 8901 2148 8957 2150
rect 8981 2148 9037 2150
rect 9061 2148 9117 2150
rect 12754 2202 12810 2204
rect 12834 2202 12890 2204
rect 12914 2202 12970 2204
rect 12994 2202 13050 2204
rect 12754 2150 12800 2202
rect 12800 2150 12810 2202
rect 12834 2150 12864 2202
rect 12864 2150 12876 2202
rect 12876 2150 12890 2202
rect 12914 2150 12928 2202
rect 12928 2150 12940 2202
rect 12940 2150 12970 2202
rect 12994 2150 13004 2202
rect 13004 2150 13050 2202
rect 12754 2148 12810 2150
rect 12834 2148 12890 2150
rect 12914 2148 12970 2150
rect 12994 2148 13050 2150
rect 16687 2202 16743 2204
rect 16767 2202 16823 2204
rect 16847 2202 16903 2204
rect 16927 2202 16983 2204
rect 16687 2150 16733 2202
rect 16733 2150 16743 2202
rect 16767 2150 16797 2202
rect 16797 2150 16809 2202
rect 16809 2150 16823 2202
rect 16847 2150 16861 2202
rect 16861 2150 16873 2202
rect 16873 2150 16903 2202
rect 16927 2150 16937 2202
rect 16937 2150 16983 2202
rect 16687 2148 16743 2150
rect 16767 2148 16823 2150
rect 16847 2148 16903 2150
rect 16927 2148 16983 2150
rect 1398 720 1454 776
<< metal3 >>
rect 0 17234 800 17264
rect 4153 17234 4219 17237
rect 0 17232 4219 17234
rect 0 17176 4158 17232
rect 4214 17176 4219 17232
rect 0 17174 4219 17176
rect 0 17144 800 17174
rect 4153 17171 4219 17174
rect 2912 15808 3228 15809
rect 0 15738 800 15768
rect 2912 15744 2918 15808
rect 2982 15744 2998 15808
rect 3062 15744 3078 15808
rect 3142 15744 3158 15808
rect 3222 15744 3228 15808
rect 2912 15743 3228 15744
rect 6845 15808 7161 15809
rect 6845 15744 6851 15808
rect 6915 15744 6931 15808
rect 6995 15744 7011 15808
rect 7075 15744 7091 15808
rect 7155 15744 7161 15808
rect 6845 15743 7161 15744
rect 10778 15808 11094 15809
rect 10778 15744 10784 15808
rect 10848 15744 10864 15808
rect 10928 15744 10944 15808
rect 11008 15744 11024 15808
rect 11088 15744 11094 15808
rect 10778 15743 11094 15744
rect 14711 15808 15027 15809
rect 14711 15744 14717 15808
rect 14781 15744 14797 15808
rect 14861 15744 14877 15808
rect 14941 15744 14957 15808
rect 15021 15744 15027 15808
rect 14711 15743 15027 15744
rect 2773 15738 2839 15741
rect 0 15736 2839 15738
rect 0 15680 2778 15736
rect 2834 15680 2839 15736
rect 0 15678 2839 15680
rect 0 15648 800 15678
rect 2773 15675 2839 15678
rect 4878 15264 5194 15265
rect 4878 15200 4884 15264
rect 4948 15200 4964 15264
rect 5028 15200 5044 15264
rect 5108 15200 5124 15264
rect 5188 15200 5194 15264
rect 4878 15199 5194 15200
rect 8811 15264 9127 15265
rect 8811 15200 8817 15264
rect 8881 15200 8897 15264
rect 8961 15200 8977 15264
rect 9041 15200 9057 15264
rect 9121 15200 9127 15264
rect 8811 15199 9127 15200
rect 12744 15264 13060 15265
rect 12744 15200 12750 15264
rect 12814 15200 12830 15264
rect 12894 15200 12910 15264
rect 12974 15200 12990 15264
rect 13054 15200 13060 15264
rect 12744 15199 13060 15200
rect 16677 15264 16993 15265
rect 16677 15200 16683 15264
rect 16747 15200 16763 15264
rect 16827 15200 16843 15264
rect 16907 15200 16923 15264
rect 16987 15200 16993 15264
rect 16677 15199 16993 15200
rect 2912 14720 3228 14721
rect 2912 14656 2918 14720
rect 2982 14656 2998 14720
rect 3062 14656 3078 14720
rect 3142 14656 3158 14720
rect 3222 14656 3228 14720
rect 2912 14655 3228 14656
rect 6845 14720 7161 14721
rect 6845 14656 6851 14720
rect 6915 14656 6931 14720
rect 6995 14656 7011 14720
rect 7075 14656 7091 14720
rect 7155 14656 7161 14720
rect 6845 14655 7161 14656
rect 10778 14720 11094 14721
rect 10778 14656 10784 14720
rect 10848 14656 10864 14720
rect 10928 14656 10944 14720
rect 11008 14656 11024 14720
rect 11088 14656 11094 14720
rect 10778 14655 11094 14656
rect 14711 14720 15027 14721
rect 14711 14656 14717 14720
rect 14781 14656 14797 14720
rect 14861 14656 14877 14720
rect 14941 14656 14957 14720
rect 15021 14656 15027 14720
rect 14711 14655 15027 14656
rect 0 14242 800 14272
rect 1669 14242 1735 14245
rect 0 14240 1735 14242
rect 0 14184 1674 14240
rect 1730 14184 1735 14240
rect 0 14182 1735 14184
rect 0 14152 800 14182
rect 1669 14179 1735 14182
rect 4878 14176 5194 14177
rect 4878 14112 4884 14176
rect 4948 14112 4964 14176
rect 5028 14112 5044 14176
rect 5108 14112 5124 14176
rect 5188 14112 5194 14176
rect 4878 14111 5194 14112
rect 8811 14176 9127 14177
rect 8811 14112 8817 14176
rect 8881 14112 8897 14176
rect 8961 14112 8977 14176
rect 9041 14112 9057 14176
rect 9121 14112 9127 14176
rect 8811 14111 9127 14112
rect 12744 14176 13060 14177
rect 12744 14112 12750 14176
rect 12814 14112 12830 14176
rect 12894 14112 12910 14176
rect 12974 14112 12990 14176
rect 13054 14112 13060 14176
rect 12744 14111 13060 14112
rect 16677 14176 16993 14177
rect 16677 14112 16683 14176
rect 16747 14112 16763 14176
rect 16827 14112 16843 14176
rect 16907 14112 16923 14176
rect 16987 14112 16993 14176
rect 16677 14111 16993 14112
rect 10869 14106 10935 14109
rect 11881 14106 11947 14109
rect 10869 14104 11947 14106
rect 10869 14048 10874 14104
rect 10930 14048 11886 14104
rect 11942 14048 11947 14104
rect 10869 14046 11947 14048
rect 10869 14043 10935 14046
rect 11881 14043 11947 14046
rect 4061 13970 4127 13973
rect 14089 13970 14155 13973
rect 4061 13968 14155 13970
rect 4061 13912 4066 13968
rect 4122 13912 14094 13968
rect 14150 13912 14155 13968
rect 4061 13910 14155 13912
rect 4061 13907 4127 13910
rect 14089 13907 14155 13910
rect 2912 13632 3228 13633
rect 2912 13568 2918 13632
rect 2982 13568 2998 13632
rect 3062 13568 3078 13632
rect 3142 13568 3158 13632
rect 3222 13568 3228 13632
rect 2912 13567 3228 13568
rect 6845 13632 7161 13633
rect 6845 13568 6851 13632
rect 6915 13568 6931 13632
rect 6995 13568 7011 13632
rect 7075 13568 7091 13632
rect 7155 13568 7161 13632
rect 6845 13567 7161 13568
rect 10778 13632 11094 13633
rect 10778 13568 10784 13632
rect 10848 13568 10864 13632
rect 10928 13568 10944 13632
rect 11008 13568 11024 13632
rect 11088 13568 11094 13632
rect 10778 13567 11094 13568
rect 14711 13632 15027 13633
rect 14711 13568 14717 13632
rect 14781 13568 14797 13632
rect 14861 13568 14877 13632
rect 14941 13568 14957 13632
rect 15021 13568 15027 13632
rect 14711 13567 15027 13568
rect 4878 13088 5194 13089
rect 4878 13024 4884 13088
rect 4948 13024 4964 13088
rect 5028 13024 5044 13088
rect 5108 13024 5124 13088
rect 5188 13024 5194 13088
rect 4878 13023 5194 13024
rect 8811 13088 9127 13089
rect 8811 13024 8817 13088
rect 8881 13024 8897 13088
rect 8961 13024 8977 13088
rect 9041 13024 9057 13088
rect 9121 13024 9127 13088
rect 8811 13023 9127 13024
rect 12744 13088 13060 13089
rect 12744 13024 12750 13088
rect 12814 13024 12830 13088
rect 12894 13024 12910 13088
rect 12974 13024 12990 13088
rect 13054 13024 13060 13088
rect 12744 13023 13060 13024
rect 16677 13088 16993 13089
rect 16677 13024 16683 13088
rect 16747 13024 16763 13088
rect 16827 13024 16843 13088
rect 16907 13024 16923 13088
rect 16987 13024 16993 13088
rect 16677 13023 16993 13024
rect 0 12746 800 12776
rect 1669 12746 1735 12749
rect 0 12744 1735 12746
rect 0 12688 1674 12744
rect 1730 12688 1735 12744
rect 0 12686 1735 12688
rect 0 12656 800 12686
rect 1669 12683 1735 12686
rect 2912 12544 3228 12545
rect 2912 12480 2918 12544
rect 2982 12480 2998 12544
rect 3062 12480 3078 12544
rect 3142 12480 3158 12544
rect 3222 12480 3228 12544
rect 2912 12479 3228 12480
rect 6845 12544 7161 12545
rect 6845 12480 6851 12544
rect 6915 12480 6931 12544
rect 6995 12480 7011 12544
rect 7075 12480 7091 12544
rect 7155 12480 7161 12544
rect 6845 12479 7161 12480
rect 10778 12544 11094 12545
rect 10778 12480 10784 12544
rect 10848 12480 10864 12544
rect 10928 12480 10944 12544
rect 11008 12480 11024 12544
rect 11088 12480 11094 12544
rect 10778 12479 11094 12480
rect 14711 12544 15027 12545
rect 14711 12480 14717 12544
rect 14781 12480 14797 12544
rect 14861 12480 14877 12544
rect 14941 12480 14957 12544
rect 15021 12480 15027 12544
rect 14711 12479 15027 12480
rect 4878 12000 5194 12001
rect 4878 11936 4884 12000
rect 4948 11936 4964 12000
rect 5028 11936 5044 12000
rect 5108 11936 5124 12000
rect 5188 11936 5194 12000
rect 4878 11935 5194 11936
rect 8811 12000 9127 12001
rect 8811 11936 8817 12000
rect 8881 11936 8897 12000
rect 8961 11936 8977 12000
rect 9041 11936 9057 12000
rect 9121 11936 9127 12000
rect 8811 11935 9127 11936
rect 12744 12000 13060 12001
rect 12744 11936 12750 12000
rect 12814 11936 12830 12000
rect 12894 11936 12910 12000
rect 12974 11936 12990 12000
rect 13054 11936 13060 12000
rect 12744 11935 13060 11936
rect 16677 12000 16993 12001
rect 16677 11936 16683 12000
rect 16747 11936 16763 12000
rect 16827 11936 16843 12000
rect 16907 11936 16923 12000
rect 16987 11936 16993 12000
rect 16677 11935 16993 11936
rect 2912 11456 3228 11457
rect 2912 11392 2918 11456
rect 2982 11392 2998 11456
rect 3062 11392 3078 11456
rect 3142 11392 3158 11456
rect 3222 11392 3228 11456
rect 2912 11391 3228 11392
rect 6845 11456 7161 11457
rect 6845 11392 6851 11456
rect 6915 11392 6931 11456
rect 6995 11392 7011 11456
rect 7075 11392 7091 11456
rect 7155 11392 7161 11456
rect 6845 11391 7161 11392
rect 10778 11456 11094 11457
rect 10778 11392 10784 11456
rect 10848 11392 10864 11456
rect 10928 11392 10944 11456
rect 11008 11392 11024 11456
rect 11088 11392 11094 11456
rect 10778 11391 11094 11392
rect 14711 11456 15027 11457
rect 14711 11392 14717 11456
rect 14781 11392 14797 11456
rect 14861 11392 14877 11456
rect 14941 11392 14957 11456
rect 15021 11392 15027 11456
rect 14711 11391 15027 11392
rect 0 11250 800 11280
rect 1669 11250 1735 11253
rect 0 11248 1735 11250
rect 0 11192 1674 11248
rect 1730 11192 1735 11248
rect 0 11190 1735 11192
rect 0 11160 800 11190
rect 1669 11187 1735 11190
rect 4878 10912 5194 10913
rect 4878 10848 4884 10912
rect 4948 10848 4964 10912
rect 5028 10848 5044 10912
rect 5108 10848 5124 10912
rect 5188 10848 5194 10912
rect 4878 10847 5194 10848
rect 8811 10912 9127 10913
rect 8811 10848 8817 10912
rect 8881 10848 8897 10912
rect 8961 10848 8977 10912
rect 9041 10848 9057 10912
rect 9121 10848 9127 10912
rect 8811 10847 9127 10848
rect 12744 10912 13060 10913
rect 12744 10848 12750 10912
rect 12814 10848 12830 10912
rect 12894 10848 12910 10912
rect 12974 10848 12990 10912
rect 13054 10848 13060 10912
rect 12744 10847 13060 10848
rect 16677 10912 16993 10913
rect 16677 10848 16683 10912
rect 16747 10848 16763 10912
rect 16827 10848 16843 10912
rect 16907 10848 16923 10912
rect 16987 10848 16993 10912
rect 16677 10847 16993 10848
rect 2912 10368 3228 10369
rect 2912 10304 2918 10368
rect 2982 10304 2998 10368
rect 3062 10304 3078 10368
rect 3142 10304 3158 10368
rect 3222 10304 3228 10368
rect 2912 10303 3228 10304
rect 6845 10368 7161 10369
rect 6845 10304 6851 10368
rect 6915 10304 6931 10368
rect 6995 10304 7011 10368
rect 7075 10304 7091 10368
rect 7155 10304 7161 10368
rect 6845 10303 7161 10304
rect 10778 10368 11094 10369
rect 10778 10304 10784 10368
rect 10848 10304 10864 10368
rect 10928 10304 10944 10368
rect 11008 10304 11024 10368
rect 11088 10304 11094 10368
rect 10778 10303 11094 10304
rect 14711 10368 15027 10369
rect 14711 10304 14717 10368
rect 14781 10304 14797 10368
rect 14861 10304 14877 10368
rect 14941 10304 14957 10368
rect 15021 10304 15027 10368
rect 14711 10303 15027 10304
rect 4878 9824 5194 9825
rect 0 9754 800 9784
rect 4878 9760 4884 9824
rect 4948 9760 4964 9824
rect 5028 9760 5044 9824
rect 5108 9760 5124 9824
rect 5188 9760 5194 9824
rect 4878 9759 5194 9760
rect 8811 9824 9127 9825
rect 8811 9760 8817 9824
rect 8881 9760 8897 9824
rect 8961 9760 8977 9824
rect 9041 9760 9057 9824
rect 9121 9760 9127 9824
rect 8811 9759 9127 9760
rect 12744 9824 13060 9825
rect 12744 9760 12750 9824
rect 12814 9760 12830 9824
rect 12894 9760 12910 9824
rect 12974 9760 12990 9824
rect 13054 9760 13060 9824
rect 12744 9759 13060 9760
rect 16677 9824 16993 9825
rect 16677 9760 16683 9824
rect 16747 9760 16763 9824
rect 16827 9760 16843 9824
rect 16907 9760 16923 9824
rect 16987 9760 16993 9824
rect 16677 9759 16993 9760
rect 1761 9754 1827 9757
rect 0 9752 1827 9754
rect 0 9696 1766 9752
rect 1822 9696 1827 9752
rect 0 9694 1827 9696
rect 0 9664 800 9694
rect 1761 9691 1827 9694
rect 3366 9692 3372 9756
rect 3436 9754 3442 9756
rect 3969 9754 4035 9757
rect 3436 9752 4035 9754
rect 3436 9696 3974 9752
rect 4030 9696 4035 9752
rect 3436 9694 4035 9696
rect 3436 9692 3442 9694
rect 3969 9691 4035 9694
rect 2912 9280 3228 9281
rect 2912 9216 2918 9280
rect 2982 9216 2998 9280
rect 3062 9216 3078 9280
rect 3142 9216 3158 9280
rect 3222 9216 3228 9280
rect 2912 9215 3228 9216
rect 6845 9280 7161 9281
rect 6845 9216 6851 9280
rect 6915 9216 6931 9280
rect 6995 9216 7011 9280
rect 7075 9216 7091 9280
rect 7155 9216 7161 9280
rect 6845 9215 7161 9216
rect 10778 9280 11094 9281
rect 10778 9216 10784 9280
rect 10848 9216 10864 9280
rect 10928 9216 10944 9280
rect 11008 9216 11024 9280
rect 11088 9216 11094 9280
rect 10778 9215 11094 9216
rect 14711 9280 15027 9281
rect 14711 9216 14717 9280
rect 14781 9216 14797 9280
rect 14861 9216 14877 9280
rect 14941 9216 14957 9280
rect 15021 9216 15027 9280
rect 14711 9215 15027 9216
rect 4878 8736 5194 8737
rect 4878 8672 4884 8736
rect 4948 8672 4964 8736
rect 5028 8672 5044 8736
rect 5108 8672 5124 8736
rect 5188 8672 5194 8736
rect 4878 8671 5194 8672
rect 8811 8736 9127 8737
rect 8811 8672 8817 8736
rect 8881 8672 8897 8736
rect 8961 8672 8977 8736
rect 9041 8672 9057 8736
rect 9121 8672 9127 8736
rect 8811 8671 9127 8672
rect 12744 8736 13060 8737
rect 12744 8672 12750 8736
rect 12814 8672 12830 8736
rect 12894 8672 12910 8736
rect 12974 8672 12990 8736
rect 13054 8672 13060 8736
rect 12744 8671 13060 8672
rect 16677 8736 16993 8737
rect 16677 8672 16683 8736
rect 16747 8672 16763 8736
rect 16827 8672 16843 8736
rect 16907 8672 16923 8736
rect 16987 8672 16993 8736
rect 16677 8671 16993 8672
rect 0 8258 800 8288
rect 1761 8258 1827 8261
rect 0 8256 1827 8258
rect 0 8200 1766 8256
rect 1822 8200 1827 8256
rect 0 8198 1827 8200
rect 0 8168 800 8198
rect 1761 8195 1827 8198
rect 2912 8192 3228 8193
rect 2912 8128 2918 8192
rect 2982 8128 2998 8192
rect 3062 8128 3078 8192
rect 3142 8128 3158 8192
rect 3222 8128 3228 8192
rect 2912 8127 3228 8128
rect 6845 8192 7161 8193
rect 6845 8128 6851 8192
rect 6915 8128 6931 8192
rect 6995 8128 7011 8192
rect 7075 8128 7091 8192
rect 7155 8128 7161 8192
rect 6845 8127 7161 8128
rect 10778 8192 11094 8193
rect 10778 8128 10784 8192
rect 10848 8128 10864 8192
rect 10928 8128 10944 8192
rect 11008 8128 11024 8192
rect 11088 8128 11094 8192
rect 10778 8127 11094 8128
rect 14711 8192 15027 8193
rect 14711 8128 14717 8192
rect 14781 8128 14797 8192
rect 14861 8128 14877 8192
rect 14941 8128 14957 8192
rect 15021 8128 15027 8192
rect 14711 8127 15027 8128
rect 4878 7648 5194 7649
rect 4878 7584 4884 7648
rect 4948 7584 4964 7648
rect 5028 7584 5044 7648
rect 5108 7584 5124 7648
rect 5188 7584 5194 7648
rect 4878 7583 5194 7584
rect 8811 7648 9127 7649
rect 8811 7584 8817 7648
rect 8881 7584 8897 7648
rect 8961 7584 8977 7648
rect 9041 7584 9057 7648
rect 9121 7584 9127 7648
rect 8811 7583 9127 7584
rect 12744 7648 13060 7649
rect 12744 7584 12750 7648
rect 12814 7584 12830 7648
rect 12894 7584 12910 7648
rect 12974 7584 12990 7648
rect 13054 7584 13060 7648
rect 12744 7583 13060 7584
rect 16677 7648 16993 7649
rect 16677 7584 16683 7648
rect 16747 7584 16763 7648
rect 16827 7584 16843 7648
rect 16907 7584 16923 7648
rect 16987 7584 16993 7648
rect 16677 7583 16993 7584
rect 5165 7306 5231 7309
rect 6729 7306 6795 7309
rect 5165 7304 6795 7306
rect 5165 7248 5170 7304
rect 5226 7248 6734 7304
rect 6790 7248 6795 7304
rect 5165 7246 6795 7248
rect 5165 7243 5231 7246
rect 6729 7243 6795 7246
rect 2912 7104 3228 7105
rect 2912 7040 2918 7104
rect 2982 7040 2998 7104
rect 3062 7040 3078 7104
rect 3142 7040 3158 7104
rect 3222 7040 3228 7104
rect 2912 7039 3228 7040
rect 6845 7104 7161 7105
rect 6845 7040 6851 7104
rect 6915 7040 6931 7104
rect 6995 7040 7011 7104
rect 7075 7040 7091 7104
rect 7155 7040 7161 7104
rect 6845 7039 7161 7040
rect 10778 7104 11094 7105
rect 10778 7040 10784 7104
rect 10848 7040 10864 7104
rect 10928 7040 10944 7104
rect 11008 7040 11024 7104
rect 11088 7040 11094 7104
rect 10778 7039 11094 7040
rect 14711 7104 15027 7105
rect 14711 7040 14717 7104
rect 14781 7040 14797 7104
rect 14861 7040 14877 7104
rect 14941 7040 14957 7104
rect 15021 7040 15027 7104
rect 14711 7039 15027 7040
rect 0 6762 800 6792
rect 1669 6762 1735 6765
rect 0 6760 1735 6762
rect 0 6704 1674 6760
rect 1730 6704 1735 6760
rect 0 6702 1735 6704
rect 0 6672 800 6702
rect 1669 6699 1735 6702
rect 4878 6560 5194 6561
rect 4878 6496 4884 6560
rect 4948 6496 4964 6560
rect 5028 6496 5044 6560
rect 5108 6496 5124 6560
rect 5188 6496 5194 6560
rect 4878 6495 5194 6496
rect 8811 6560 9127 6561
rect 8811 6496 8817 6560
rect 8881 6496 8897 6560
rect 8961 6496 8977 6560
rect 9041 6496 9057 6560
rect 9121 6496 9127 6560
rect 8811 6495 9127 6496
rect 12744 6560 13060 6561
rect 12744 6496 12750 6560
rect 12814 6496 12830 6560
rect 12894 6496 12910 6560
rect 12974 6496 12990 6560
rect 13054 6496 13060 6560
rect 12744 6495 13060 6496
rect 16677 6560 16993 6561
rect 16677 6496 16683 6560
rect 16747 6496 16763 6560
rect 16827 6496 16843 6560
rect 16907 6496 16923 6560
rect 16987 6496 16993 6560
rect 16677 6495 16993 6496
rect 2912 6016 3228 6017
rect 2912 5952 2918 6016
rect 2982 5952 2998 6016
rect 3062 5952 3078 6016
rect 3142 5952 3158 6016
rect 3222 5952 3228 6016
rect 2912 5951 3228 5952
rect 6845 6016 7161 6017
rect 6845 5952 6851 6016
rect 6915 5952 6931 6016
rect 6995 5952 7011 6016
rect 7075 5952 7091 6016
rect 7155 5952 7161 6016
rect 6845 5951 7161 5952
rect 10778 6016 11094 6017
rect 10778 5952 10784 6016
rect 10848 5952 10864 6016
rect 10928 5952 10944 6016
rect 11008 5952 11024 6016
rect 11088 5952 11094 6016
rect 10778 5951 11094 5952
rect 14711 6016 15027 6017
rect 14711 5952 14717 6016
rect 14781 5952 14797 6016
rect 14861 5952 14877 6016
rect 14941 5952 14957 6016
rect 15021 5952 15027 6016
rect 14711 5951 15027 5952
rect 4878 5472 5194 5473
rect 4878 5408 4884 5472
rect 4948 5408 4964 5472
rect 5028 5408 5044 5472
rect 5108 5408 5124 5472
rect 5188 5408 5194 5472
rect 4878 5407 5194 5408
rect 8811 5472 9127 5473
rect 8811 5408 8817 5472
rect 8881 5408 8897 5472
rect 8961 5408 8977 5472
rect 9041 5408 9057 5472
rect 9121 5408 9127 5472
rect 8811 5407 9127 5408
rect 12744 5472 13060 5473
rect 12744 5408 12750 5472
rect 12814 5408 12830 5472
rect 12894 5408 12910 5472
rect 12974 5408 12990 5472
rect 13054 5408 13060 5472
rect 12744 5407 13060 5408
rect 16677 5472 16993 5473
rect 16677 5408 16683 5472
rect 16747 5408 16763 5472
rect 16827 5408 16843 5472
rect 16907 5408 16923 5472
rect 16987 5408 16993 5472
rect 16677 5407 16993 5408
rect 0 5266 800 5296
rect 1485 5266 1551 5269
rect 0 5264 1551 5266
rect 0 5208 1490 5264
rect 1546 5208 1551 5264
rect 0 5206 1551 5208
rect 0 5176 800 5206
rect 1485 5203 1551 5206
rect 2912 4928 3228 4929
rect 2912 4864 2918 4928
rect 2982 4864 2998 4928
rect 3062 4864 3078 4928
rect 3142 4864 3158 4928
rect 3222 4864 3228 4928
rect 2912 4863 3228 4864
rect 6845 4928 7161 4929
rect 6845 4864 6851 4928
rect 6915 4864 6931 4928
rect 6995 4864 7011 4928
rect 7075 4864 7091 4928
rect 7155 4864 7161 4928
rect 6845 4863 7161 4864
rect 10778 4928 11094 4929
rect 10778 4864 10784 4928
rect 10848 4864 10864 4928
rect 10928 4864 10944 4928
rect 11008 4864 11024 4928
rect 11088 4864 11094 4928
rect 10778 4863 11094 4864
rect 14711 4928 15027 4929
rect 14711 4864 14717 4928
rect 14781 4864 14797 4928
rect 14861 4864 14877 4928
rect 14941 4864 14957 4928
rect 15021 4864 15027 4928
rect 14711 4863 15027 4864
rect 4878 4384 5194 4385
rect 4878 4320 4884 4384
rect 4948 4320 4964 4384
rect 5028 4320 5044 4384
rect 5108 4320 5124 4384
rect 5188 4320 5194 4384
rect 4878 4319 5194 4320
rect 8811 4384 9127 4385
rect 8811 4320 8817 4384
rect 8881 4320 8897 4384
rect 8961 4320 8977 4384
rect 9041 4320 9057 4384
rect 9121 4320 9127 4384
rect 8811 4319 9127 4320
rect 12744 4384 13060 4385
rect 12744 4320 12750 4384
rect 12814 4320 12830 4384
rect 12894 4320 12910 4384
rect 12974 4320 12990 4384
rect 13054 4320 13060 4384
rect 12744 4319 13060 4320
rect 16677 4384 16993 4385
rect 16677 4320 16683 4384
rect 16747 4320 16763 4384
rect 16827 4320 16843 4384
rect 16907 4320 16923 4384
rect 16987 4320 16993 4384
rect 16677 4319 16993 4320
rect 2037 4042 2103 4045
rect 3366 4042 3372 4044
rect 2037 4040 3372 4042
rect 2037 3984 2042 4040
rect 2098 3984 3372 4040
rect 2037 3982 3372 3984
rect 2037 3979 2103 3982
rect 3366 3980 3372 3982
rect 3436 3980 3442 4044
rect 2912 3840 3228 3841
rect 0 3770 800 3800
rect 2912 3776 2918 3840
rect 2982 3776 2998 3840
rect 3062 3776 3078 3840
rect 3142 3776 3158 3840
rect 3222 3776 3228 3840
rect 2912 3775 3228 3776
rect 6845 3840 7161 3841
rect 6845 3776 6851 3840
rect 6915 3776 6931 3840
rect 6995 3776 7011 3840
rect 7075 3776 7091 3840
rect 7155 3776 7161 3840
rect 6845 3775 7161 3776
rect 10778 3840 11094 3841
rect 10778 3776 10784 3840
rect 10848 3776 10864 3840
rect 10928 3776 10944 3840
rect 11008 3776 11024 3840
rect 11088 3776 11094 3840
rect 10778 3775 11094 3776
rect 14711 3840 15027 3841
rect 14711 3776 14717 3840
rect 14781 3776 14797 3840
rect 14861 3776 14877 3840
rect 14941 3776 14957 3840
rect 15021 3776 15027 3840
rect 14711 3775 15027 3776
rect 1393 3770 1459 3773
rect 0 3768 1459 3770
rect 0 3712 1398 3768
rect 1454 3712 1459 3768
rect 0 3710 1459 3712
rect 0 3680 800 3710
rect 1393 3707 1459 3710
rect 4878 3296 5194 3297
rect 4878 3232 4884 3296
rect 4948 3232 4964 3296
rect 5028 3232 5044 3296
rect 5108 3232 5124 3296
rect 5188 3232 5194 3296
rect 4878 3231 5194 3232
rect 8811 3296 9127 3297
rect 8811 3232 8817 3296
rect 8881 3232 8897 3296
rect 8961 3232 8977 3296
rect 9041 3232 9057 3296
rect 9121 3232 9127 3296
rect 8811 3231 9127 3232
rect 12744 3296 13060 3297
rect 12744 3232 12750 3296
rect 12814 3232 12830 3296
rect 12894 3232 12910 3296
rect 12974 3232 12990 3296
rect 13054 3232 13060 3296
rect 12744 3231 13060 3232
rect 16677 3296 16993 3297
rect 16677 3232 16683 3296
rect 16747 3232 16763 3296
rect 16827 3232 16843 3296
rect 16907 3232 16923 3296
rect 16987 3232 16993 3296
rect 16677 3231 16993 3232
rect 2912 2752 3228 2753
rect 2912 2688 2918 2752
rect 2982 2688 2998 2752
rect 3062 2688 3078 2752
rect 3142 2688 3158 2752
rect 3222 2688 3228 2752
rect 2912 2687 3228 2688
rect 6845 2752 7161 2753
rect 6845 2688 6851 2752
rect 6915 2688 6931 2752
rect 6995 2688 7011 2752
rect 7075 2688 7091 2752
rect 7155 2688 7161 2752
rect 6845 2687 7161 2688
rect 10778 2752 11094 2753
rect 10778 2688 10784 2752
rect 10848 2688 10864 2752
rect 10928 2688 10944 2752
rect 11008 2688 11024 2752
rect 11088 2688 11094 2752
rect 10778 2687 11094 2688
rect 14711 2752 15027 2753
rect 14711 2688 14717 2752
rect 14781 2688 14797 2752
rect 14861 2688 14877 2752
rect 14941 2688 14957 2752
rect 15021 2688 15027 2752
rect 14711 2687 15027 2688
rect 0 2274 800 2304
rect 1761 2274 1827 2277
rect 0 2272 1827 2274
rect 0 2216 1766 2272
rect 1822 2216 1827 2272
rect 0 2214 1827 2216
rect 0 2184 800 2214
rect 1761 2211 1827 2214
rect 4878 2208 5194 2209
rect 4878 2144 4884 2208
rect 4948 2144 4964 2208
rect 5028 2144 5044 2208
rect 5108 2144 5124 2208
rect 5188 2144 5194 2208
rect 4878 2143 5194 2144
rect 8811 2208 9127 2209
rect 8811 2144 8817 2208
rect 8881 2144 8897 2208
rect 8961 2144 8977 2208
rect 9041 2144 9057 2208
rect 9121 2144 9127 2208
rect 8811 2143 9127 2144
rect 12744 2208 13060 2209
rect 12744 2144 12750 2208
rect 12814 2144 12830 2208
rect 12894 2144 12910 2208
rect 12974 2144 12990 2208
rect 13054 2144 13060 2208
rect 12744 2143 13060 2144
rect 16677 2208 16993 2209
rect 16677 2144 16683 2208
rect 16747 2144 16763 2208
rect 16827 2144 16843 2208
rect 16907 2144 16923 2208
rect 16987 2144 16993 2208
rect 16677 2143 16993 2144
rect 0 778 800 808
rect 1393 778 1459 781
rect 0 776 1459 778
rect 0 720 1398 776
rect 1454 720 1459 776
rect 0 718 1459 720
rect 0 688 800 718
rect 1393 715 1459 718
<< via3 >>
rect 2918 15804 2982 15808
rect 2918 15748 2922 15804
rect 2922 15748 2978 15804
rect 2978 15748 2982 15804
rect 2918 15744 2982 15748
rect 2998 15804 3062 15808
rect 2998 15748 3002 15804
rect 3002 15748 3058 15804
rect 3058 15748 3062 15804
rect 2998 15744 3062 15748
rect 3078 15804 3142 15808
rect 3078 15748 3082 15804
rect 3082 15748 3138 15804
rect 3138 15748 3142 15804
rect 3078 15744 3142 15748
rect 3158 15804 3222 15808
rect 3158 15748 3162 15804
rect 3162 15748 3218 15804
rect 3218 15748 3222 15804
rect 3158 15744 3222 15748
rect 6851 15804 6915 15808
rect 6851 15748 6855 15804
rect 6855 15748 6911 15804
rect 6911 15748 6915 15804
rect 6851 15744 6915 15748
rect 6931 15804 6995 15808
rect 6931 15748 6935 15804
rect 6935 15748 6991 15804
rect 6991 15748 6995 15804
rect 6931 15744 6995 15748
rect 7011 15804 7075 15808
rect 7011 15748 7015 15804
rect 7015 15748 7071 15804
rect 7071 15748 7075 15804
rect 7011 15744 7075 15748
rect 7091 15804 7155 15808
rect 7091 15748 7095 15804
rect 7095 15748 7151 15804
rect 7151 15748 7155 15804
rect 7091 15744 7155 15748
rect 10784 15804 10848 15808
rect 10784 15748 10788 15804
rect 10788 15748 10844 15804
rect 10844 15748 10848 15804
rect 10784 15744 10848 15748
rect 10864 15804 10928 15808
rect 10864 15748 10868 15804
rect 10868 15748 10924 15804
rect 10924 15748 10928 15804
rect 10864 15744 10928 15748
rect 10944 15804 11008 15808
rect 10944 15748 10948 15804
rect 10948 15748 11004 15804
rect 11004 15748 11008 15804
rect 10944 15744 11008 15748
rect 11024 15804 11088 15808
rect 11024 15748 11028 15804
rect 11028 15748 11084 15804
rect 11084 15748 11088 15804
rect 11024 15744 11088 15748
rect 14717 15804 14781 15808
rect 14717 15748 14721 15804
rect 14721 15748 14777 15804
rect 14777 15748 14781 15804
rect 14717 15744 14781 15748
rect 14797 15804 14861 15808
rect 14797 15748 14801 15804
rect 14801 15748 14857 15804
rect 14857 15748 14861 15804
rect 14797 15744 14861 15748
rect 14877 15804 14941 15808
rect 14877 15748 14881 15804
rect 14881 15748 14937 15804
rect 14937 15748 14941 15804
rect 14877 15744 14941 15748
rect 14957 15804 15021 15808
rect 14957 15748 14961 15804
rect 14961 15748 15017 15804
rect 15017 15748 15021 15804
rect 14957 15744 15021 15748
rect 4884 15260 4948 15264
rect 4884 15204 4888 15260
rect 4888 15204 4944 15260
rect 4944 15204 4948 15260
rect 4884 15200 4948 15204
rect 4964 15260 5028 15264
rect 4964 15204 4968 15260
rect 4968 15204 5024 15260
rect 5024 15204 5028 15260
rect 4964 15200 5028 15204
rect 5044 15260 5108 15264
rect 5044 15204 5048 15260
rect 5048 15204 5104 15260
rect 5104 15204 5108 15260
rect 5044 15200 5108 15204
rect 5124 15260 5188 15264
rect 5124 15204 5128 15260
rect 5128 15204 5184 15260
rect 5184 15204 5188 15260
rect 5124 15200 5188 15204
rect 8817 15260 8881 15264
rect 8817 15204 8821 15260
rect 8821 15204 8877 15260
rect 8877 15204 8881 15260
rect 8817 15200 8881 15204
rect 8897 15260 8961 15264
rect 8897 15204 8901 15260
rect 8901 15204 8957 15260
rect 8957 15204 8961 15260
rect 8897 15200 8961 15204
rect 8977 15260 9041 15264
rect 8977 15204 8981 15260
rect 8981 15204 9037 15260
rect 9037 15204 9041 15260
rect 8977 15200 9041 15204
rect 9057 15260 9121 15264
rect 9057 15204 9061 15260
rect 9061 15204 9117 15260
rect 9117 15204 9121 15260
rect 9057 15200 9121 15204
rect 12750 15260 12814 15264
rect 12750 15204 12754 15260
rect 12754 15204 12810 15260
rect 12810 15204 12814 15260
rect 12750 15200 12814 15204
rect 12830 15260 12894 15264
rect 12830 15204 12834 15260
rect 12834 15204 12890 15260
rect 12890 15204 12894 15260
rect 12830 15200 12894 15204
rect 12910 15260 12974 15264
rect 12910 15204 12914 15260
rect 12914 15204 12970 15260
rect 12970 15204 12974 15260
rect 12910 15200 12974 15204
rect 12990 15260 13054 15264
rect 12990 15204 12994 15260
rect 12994 15204 13050 15260
rect 13050 15204 13054 15260
rect 12990 15200 13054 15204
rect 16683 15260 16747 15264
rect 16683 15204 16687 15260
rect 16687 15204 16743 15260
rect 16743 15204 16747 15260
rect 16683 15200 16747 15204
rect 16763 15260 16827 15264
rect 16763 15204 16767 15260
rect 16767 15204 16823 15260
rect 16823 15204 16827 15260
rect 16763 15200 16827 15204
rect 16843 15260 16907 15264
rect 16843 15204 16847 15260
rect 16847 15204 16903 15260
rect 16903 15204 16907 15260
rect 16843 15200 16907 15204
rect 16923 15260 16987 15264
rect 16923 15204 16927 15260
rect 16927 15204 16983 15260
rect 16983 15204 16987 15260
rect 16923 15200 16987 15204
rect 2918 14716 2982 14720
rect 2918 14660 2922 14716
rect 2922 14660 2978 14716
rect 2978 14660 2982 14716
rect 2918 14656 2982 14660
rect 2998 14716 3062 14720
rect 2998 14660 3002 14716
rect 3002 14660 3058 14716
rect 3058 14660 3062 14716
rect 2998 14656 3062 14660
rect 3078 14716 3142 14720
rect 3078 14660 3082 14716
rect 3082 14660 3138 14716
rect 3138 14660 3142 14716
rect 3078 14656 3142 14660
rect 3158 14716 3222 14720
rect 3158 14660 3162 14716
rect 3162 14660 3218 14716
rect 3218 14660 3222 14716
rect 3158 14656 3222 14660
rect 6851 14716 6915 14720
rect 6851 14660 6855 14716
rect 6855 14660 6911 14716
rect 6911 14660 6915 14716
rect 6851 14656 6915 14660
rect 6931 14716 6995 14720
rect 6931 14660 6935 14716
rect 6935 14660 6991 14716
rect 6991 14660 6995 14716
rect 6931 14656 6995 14660
rect 7011 14716 7075 14720
rect 7011 14660 7015 14716
rect 7015 14660 7071 14716
rect 7071 14660 7075 14716
rect 7011 14656 7075 14660
rect 7091 14716 7155 14720
rect 7091 14660 7095 14716
rect 7095 14660 7151 14716
rect 7151 14660 7155 14716
rect 7091 14656 7155 14660
rect 10784 14716 10848 14720
rect 10784 14660 10788 14716
rect 10788 14660 10844 14716
rect 10844 14660 10848 14716
rect 10784 14656 10848 14660
rect 10864 14716 10928 14720
rect 10864 14660 10868 14716
rect 10868 14660 10924 14716
rect 10924 14660 10928 14716
rect 10864 14656 10928 14660
rect 10944 14716 11008 14720
rect 10944 14660 10948 14716
rect 10948 14660 11004 14716
rect 11004 14660 11008 14716
rect 10944 14656 11008 14660
rect 11024 14716 11088 14720
rect 11024 14660 11028 14716
rect 11028 14660 11084 14716
rect 11084 14660 11088 14716
rect 11024 14656 11088 14660
rect 14717 14716 14781 14720
rect 14717 14660 14721 14716
rect 14721 14660 14777 14716
rect 14777 14660 14781 14716
rect 14717 14656 14781 14660
rect 14797 14716 14861 14720
rect 14797 14660 14801 14716
rect 14801 14660 14857 14716
rect 14857 14660 14861 14716
rect 14797 14656 14861 14660
rect 14877 14716 14941 14720
rect 14877 14660 14881 14716
rect 14881 14660 14937 14716
rect 14937 14660 14941 14716
rect 14877 14656 14941 14660
rect 14957 14716 15021 14720
rect 14957 14660 14961 14716
rect 14961 14660 15017 14716
rect 15017 14660 15021 14716
rect 14957 14656 15021 14660
rect 4884 14172 4948 14176
rect 4884 14116 4888 14172
rect 4888 14116 4944 14172
rect 4944 14116 4948 14172
rect 4884 14112 4948 14116
rect 4964 14172 5028 14176
rect 4964 14116 4968 14172
rect 4968 14116 5024 14172
rect 5024 14116 5028 14172
rect 4964 14112 5028 14116
rect 5044 14172 5108 14176
rect 5044 14116 5048 14172
rect 5048 14116 5104 14172
rect 5104 14116 5108 14172
rect 5044 14112 5108 14116
rect 5124 14172 5188 14176
rect 5124 14116 5128 14172
rect 5128 14116 5184 14172
rect 5184 14116 5188 14172
rect 5124 14112 5188 14116
rect 8817 14172 8881 14176
rect 8817 14116 8821 14172
rect 8821 14116 8877 14172
rect 8877 14116 8881 14172
rect 8817 14112 8881 14116
rect 8897 14172 8961 14176
rect 8897 14116 8901 14172
rect 8901 14116 8957 14172
rect 8957 14116 8961 14172
rect 8897 14112 8961 14116
rect 8977 14172 9041 14176
rect 8977 14116 8981 14172
rect 8981 14116 9037 14172
rect 9037 14116 9041 14172
rect 8977 14112 9041 14116
rect 9057 14172 9121 14176
rect 9057 14116 9061 14172
rect 9061 14116 9117 14172
rect 9117 14116 9121 14172
rect 9057 14112 9121 14116
rect 12750 14172 12814 14176
rect 12750 14116 12754 14172
rect 12754 14116 12810 14172
rect 12810 14116 12814 14172
rect 12750 14112 12814 14116
rect 12830 14172 12894 14176
rect 12830 14116 12834 14172
rect 12834 14116 12890 14172
rect 12890 14116 12894 14172
rect 12830 14112 12894 14116
rect 12910 14172 12974 14176
rect 12910 14116 12914 14172
rect 12914 14116 12970 14172
rect 12970 14116 12974 14172
rect 12910 14112 12974 14116
rect 12990 14172 13054 14176
rect 12990 14116 12994 14172
rect 12994 14116 13050 14172
rect 13050 14116 13054 14172
rect 12990 14112 13054 14116
rect 16683 14172 16747 14176
rect 16683 14116 16687 14172
rect 16687 14116 16743 14172
rect 16743 14116 16747 14172
rect 16683 14112 16747 14116
rect 16763 14172 16827 14176
rect 16763 14116 16767 14172
rect 16767 14116 16823 14172
rect 16823 14116 16827 14172
rect 16763 14112 16827 14116
rect 16843 14172 16907 14176
rect 16843 14116 16847 14172
rect 16847 14116 16903 14172
rect 16903 14116 16907 14172
rect 16843 14112 16907 14116
rect 16923 14172 16987 14176
rect 16923 14116 16927 14172
rect 16927 14116 16983 14172
rect 16983 14116 16987 14172
rect 16923 14112 16987 14116
rect 2918 13628 2982 13632
rect 2918 13572 2922 13628
rect 2922 13572 2978 13628
rect 2978 13572 2982 13628
rect 2918 13568 2982 13572
rect 2998 13628 3062 13632
rect 2998 13572 3002 13628
rect 3002 13572 3058 13628
rect 3058 13572 3062 13628
rect 2998 13568 3062 13572
rect 3078 13628 3142 13632
rect 3078 13572 3082 13628
rect 3082 13572 3138 13628
rect 3138 13572 3142 13628
rect 3078 13568 3142 13572
rect 3158 13628 3222 13632
rect 3158 13572 3162 13628
rect 3162 13572 3218 13628
rect 3218 13572 3222 13628
rect 3158 13568 3222 13572
rect 6851 13628 6915 13632
rect 6851 13572 6855 13628
rect 6855 13572 6911 13628
rect 6911 13572 6915 13628
rect 6851 13568 6915 13572
rect 6931 13628 6995 13632
rect 6931 13572 6935 13628
rect 6935 13572 6991 13628
rect 6991 13572 6995 13628
rect 6931 13568 6995 13572
rect 7011 13628 7075 13632
rect 7011 13572 7015 13628
rect 7015 13572 7071 13628
rect 7071 13572 7075 13628
rect 7011 13568 7075 13572
rect 7091 13628 7155 13632
rect 7091 13572 7095 13628
rect 7095 13572 7151 13628
rect 7151 13572 7155 13628
rect 7091 13568 7155 13572
rect 10784 13628 10848 13632
rect 10784 13572 10788 13628
rect 10788 13572 10844 13628
rect 10844 13572 10848 13628
rect 10784 13568 10848 13572
rect 10864 13628 10928 13632
rect 10864 13572 10868 13628
rect 10868 13572 10924 13628
rect 10924 13572 10928 13628
rect 10864 13568 10928 13572
rect 10944 13628 11008 13632
rect 10944 13572 10948 13628
rect 10948 13572 11004 13628
rect 11004 13572 11008 13628
rect 10944 13568 11008 13572
rect 11024 13628 11088 13632
rect 11024 13572 11028 13628
rect 11028 13572 11084 13628
rect 11084 13572 11088 13628
rect 11024 13568 11088 13572
rect 14717 13628 14781 13632
rect 14717 13572 14721 13628
rect 14721 13572 14777 13628
rect 14777 13572 14781 13628
rect 14717 13568 14781 13572
rect 14797 13628 14861 13632
rect 14797 13572 14801 13628
rect 14801 13572 14857 13628
rect 14857 13572 14861 13628
rect 14797 13568 14861 13572
rect 14877 13628 14941 13632
rect 14877 13572 14881 13628
rect 14881 13572 14937 13628
rect 14937 13572 14941 13628
rect 14877 13568 14941 13572
rect 14957 13628 15021 13632
rect 14957 13572 14961 13628
rect 14961 13572 15017 13628
rect 15017 13572 15021 13628
rect 14957 13568 15021 13572
rect 4884 13084 4948 13088
rect 4884 13028 4888 13084
rect 4888 13028 4944 13084
rect 4944 13028 4948 13084
rect 4884 13024 4948 13028
rect 4964 13084 5028 13088
rect 4964 13028 4968 13084
rect 4968 13028 5024 13084
rect 5024 13028 5028 13084
rect 4964 13024 5028 13028
rect 5044 13084 5108 13088
rect 5044 13028 5048 13084
rect 5048 13028 5104 13084
rect 5104 13028 5108 13084
rect 5044 13024 5108 13028
rect 5124 13084 5188 13088
rect 5124 13028 5128 13084
rect 5128 13028 5184 13084
rect 5184 13028 5188 13084
rect 5124 13024 5188 13028
rect 8817 13084 8881 13088
rect 8817 13028 8821 13084
rect 8821 13028 8877 13084
rect 8877 13028 8881 13084
rect 8817 13024 8881 13028
rect 8897 13084 8961 13088
rect 8897 13028 8901 13084
rect 8901 13028 8957 13084
rect 8957 13028 8961 13084
rect 8897 13024 8961 13028
rect 8977 13084 9041 13088
rect 8977 13028 8981 13084
rect 8981 13028 9037 13084
rect 9037 13028 9041 13084
rect 8977 13024 9041 13028
rect 9057 13084 9121 13088
rect 9057 13028 9061 13084
rect 9061 13028 9117 13084
rect 9117 13028 9121 13084
rect 9057 13024 9121 13028
rect 12750 13084 12814 13088
rect 12750 13028 12754 13084
rect 12754 13028 12810 13084
rect 12810 13028 12814 13084
rect 12750 13024 12814 13028
rect 12830 13084 12894 13088
rect 12830 13028 12834 13084
rect 12834 13028 12890 13084
rect 12890 13028 12894 13084
rect 12830 13024 12894 13028
rect 12910 13084 12974 13088
rect 12910 13028 12914 13084
rect 12914 13028 12970 13084
rect 12970 13028 12974 13084
rect 12910 13024 12974 13028
rect 12990 13084 13054 13088
rect 12990 13028 12994 13084
rect 12994 13028 13050 13084
rect 13050 13028 13054 13084
rect 12990 13024 13054 13028
rect 16683 13084 16747 13088
rect 16683 13028 16687 13084
rect 16687 13028 16743 13084
rect 16743 13028 16747 13084
rect 16683 13024 16747 13028
rect 16763 13084 16827 13088
rect 16763 13028 16767 13084
rect 16767 13028 16823 13084
rect 16823 13028 16827 13084
rect 16763 13024 16827 13028
rect 16843 13084 16907 13088
rect 16843 13028 16847 13084
rect 16847 13028 16903 13084
rect 16903 13028 16907 13084
rect 16843 13024 16907 13028
rect 16923 13084 16987 13088
rect 16923 13028 16927 13084
rect 16927 13028 16983 13084
rect 16983 13028 16987 13084
rect 16923 13024 16987 13028
rect 2918 12540 2982 12544
rect 2918 12484 2922 12540
rect 2922 12484 2978 12540
rect 2978 12484 2982 12540
rect 2918 12480 2982 12484
rect 2998 12540 3062 12544
rect 2998 12484 3002 12540
rect 3002 12484 3058 12540
rect 3058 12484 3062 12540
rect 2998 12480 3062 12484
rect 3078 12540 3142 12544
rect 3078 12484 3082 12540
rect 3082 12484 3138 12540
rect 3138 12484 3142 12540
rect 3078 12480 3142 12484
rect 3158 12540 3222 12544
rect 3158 12484 3162 12540
rect 3162 12484 3218 12540
rect 3218 12484 3222 12540
rect 3158 12480 3222 12484
rect 6851 12540 6915 12544
rect 6851 12484 6855 12540
rect 6855 12484 6911 12540
rect 6911 12484 6915 12540
rect 6851 12480 6915 12484
rect 6931 12540 6995 12544
rect 6931 12484 6935 12540
rect 6935 12484 6991 12540
rect 6991 12484 6995 12540
rect 6931 12480 6995 12484
rect 7011 12540 7075 12544
rect 7011 12484 7015 12540
rect 7015 12484 7071 12540
rect 7071 12484 7075 12540
rect 7011 12480 7075 12484
rect 7091 12540 7155 12544
rect 7091 12484 7095 12540
rect 7095 12484 7151 12540
rect 7151 12484 7155 12540
rect 7091 12480 7155 12484
rect 10784 12540 10848 12544
rect 10784 12484 10788 12540
rect 10788 12484 10844 12540
rect 10844 12484 10848 12540
rect 10784 12480 10848 12484
rect 10864 12540 10928 12544
rect 10864 12484 10868 12540
rect 10868 12484 10924 12540
rect 10924 12484 10928 12540
rect 10864 12480 10928 12484
rect 10944 12540 11008 12544
rect 10944 12484 10948 12540
rect 10948 12484 11004 12540
rect 11004 12484 11008 12540
rect 10944 12480 11008 12484
rect 11024 12540 11088 12544
rect 11024 12484 11028 12540
rect 11028 12484 11084 12540
rect 11084 12484 11088 12540
rect 11024 12480 11088 12484
rect 14717 12540 14781 12544
rect 14717 12484 14721 12540
rect 14721 12484 14777 12540
rect 14777 12484 14781 12540
rect 14717 12480 14781 12484
rect 14797 12540 14861 12544
rect 14797 12484 14801 12540
rect 14801 12484 14857 12540
rect 14857 12484 14861 12540
rect 14797 12480 14861 12484
rect 14877 12540 14941 12544
rect 14877 12484 14881 12540
rect 14881 12484 14937 12540
rect 14937 12484 14941 12540
rect 14877 12480 14941 12484
rect 14957 12540 15021 12544
rect 14957 12484 14961 12540
rect 14961 12484 15017 12540
rect 15017 12484 15021 12540
rect 14957 12480 15021 12484
rect 4884 11996 4948 12000
rect 4884 11940 4888 11996
rect 4888 11940 4944 11996
rect 4944 11940 4948 11996
rect 4884 11936 4948 11940
rect 4964 11996 5028 12000
rect 4964 11940 4968 11996
rect 4968 11940 5024 11996
rect 5024 11940 5028 11996
rect 4964 11936 5028 11940
rect 5044 11996 5108 12000
rect 5044 11940 5048 11996
rect 5048 11940 5104 11996
rect 5104 11940 5108 11996
rect 5044 11936 5108 11940
rect 5124 11996 5188 12000
rect 5124 11940 5128 11996
rect 5128 11940 5184 11996
rect 5184 11940 5188 11996
rect 5124 11936 5188 11940
rect 8817 11996 8881 12000
rect 8817 11940 8821 11996
rect 8821 11940 8877 11996
rect 8877 11940 8881 11996
rect 8817 11936 8881 11940
rect 8897 11996 8961 12000
rect 8897 11940 8901 11996
rect 8901 11940 8957 11996
rect 8957 11940 8961 11996
rect 8897 11936 8961 11940
rect 8977 11996 9041 12000
rect 8977 11940 8981 11996
rect 8981 11940 9037 11996
rect 9037 11940 9041 11996
rect 8977 11936 9041 11940
rect 9057 11996 9121 12000
rect 9057 11940 9061 11996
rect 9061 11940 9117 11996
rect 9117 11940 9121 11996
rect 9057 11936 9121 11940
rect 12750 11996 12814 12000
rect 12750 11940 12754 11996
rect 12754 11940 12810 11996
rect 12810 11940 12814 11996
rect 12750 11936 12814 11940
rect 12830 11996 12894 12000
rect 12830 11940 12834 11996
rect 12834 11940 12890 11996
rect 12890 11940 12894 11996
rect 12830 11936 12894 11940
rect 12910 11996 12974 12000
rect 12910 11940 12914 11996
rect 12914 11940 12970 11996
rect 12970 11940 12974 11996
rect 12910 11936 12974 11940
rect 12990 11996 13054 12000
rect 12990 11940 12994 11996
rect 12994 11940 13050 11996
rect 13050 11940 13054 11996
rect 12990 11936 13054 11940
rect 16683 11996 16747 12000
rect 16683 11940 16687 11996
rect 16687 11940 16743 11996
rect 16743 11940 16747 11996
rect 16683 11936 16747 11940
rect 16763 11996 16827 12000
rect 16763 11940 16767 11996
rect 16767 11940 16823 11996
rect 16823 11940 16827 11996
rect 16763 11936 16827 11940
rect 16843 11996 16907 12000
rect 16843 11940 16847 11996
rect 16847 11940 16903 11996
rect 16903 11940 16907 11996
rect 16843 11936 16907 11940
rect 16923 11996 16987 12000
rect 16923 11940 16927 11996
rect 16927 11940 16983 11996
rect 16983 11940 16987 11996
rect 16923 11936 16987 11940
rect 2918 11452 2982 11456
rect 2918 11396 2922 11452
rect 2922 11396 2978 11452
rect 2978 11396 2982 11452
rect 2918 11392 2982 11396
rect 2998 11452 3062 11456
rect 2998 11396 3002 11452
rect 3002 11396 3058 11452
rect 3058 11396 3062 11452
rect 2998 11392 3062 11396
rect 3078 11452 3142 11456
rect 3078 11396 3082 11452
rect 3082 11396 3138 11452
rect 3138 11396 3142 11452
rect 3078 11392 3142 11396
rect 3158 11452 3222 11456
rect 3158 11396 3162 11452
rect 3162 11396 3218 11452
rect 3218 11396 3222 11452
rect 3158 11392 3222 11396
rect 6851 11452 6915 11456
rect 6851 11396 6855 11452
rect 6855 11396 6911 11452
rect 6911 11396 6915 11452
rect 6851 11392 6915 11396
rect 6931 11452 6995 11456
rect 6931 11396 6935 11452
rect 6935 11396 6991 11452
rect 6991 11396 6995 11452
rect 6931 11392 6995 11396
rect 7011 11452 7075 11456
rect 7011 11396 7015 11452
rect 7015 11396 7071 11452
rect 7071 11396 7075 11452
rect 7011 11392 7075 11396
rect 7091 11452 7155 11456
rect 7091 11396 7095 11452
rect 7095 11396 7151 11452
rect 7151 11396 7155 11452
rect 7091 11392 7155 11396
rect 10784 11452 10848 11456
rect 10784 11396 10788 11452
rect 10788 11396 10844 11452
rect 10844 11396 10848 11452
rect 10784 11392 10848 11396
rect 10864 11452 10928 11456
rect 10864 11396 10868 11452
rect 10868 11396 10924 11452
rect 10924 11396 10928 11452
rect 10864 11392 10928 11396
rect 10944 11452 11008 11456
rect 10944 11396 10948 11452
rect 10948 11396 11004 11452
rect 11004 11396 11008 11452
rect 10944 11392 11008 11396
rect 11024 11452 11088 11456
rect 11024 11396 11028 11452
rect 11028 11396 11084 11452
rect 11084 11396 11088 11452
rect 11024 11392 11088 11396
rect 14717 11452 14781 11456
rect 14717 11396 14721 11452
rect 14721 11396 14777 11452
rect 14777 11396 14781 11452
rect 14717 11392 14781 11396
rect 14797 11452 14861 11456
rect 14797 11396 14801 11452
rect 14801 11396 14857 11452
rect 14857 11396 14861 11452
rect 14797 11392 14861 11396
rect 14877 11452 14941 11456
rect 14877 11396 14881 11452
rect 14881 11396 14937 11452
rect 14937 11396 14941 11452
rect 14877 11392 14941 11396
rect 14957 11452 15021 11456
rect 14957 11396 14961 11452
rect 14961 11396 15017 11452
rect 15017 11396 15021 11452
rect 14957 11392 15021 11396
rect 4884 10908 4948 10912
rect 4884 10852 4888 10908
rect 4888 10852 4944 10908
rect 4944 10852 4948 10908
rect 4884 10848 4948 10852
rect 4964 10908 5028 10912
rect 4964 10852 4968 10908
rect 4968 10852 5024 10908
rect 5024 10852 5028 10908
rect 4964 10848 5028 10852
rect 5044 10908 5108 10912
rect 5044 10852 5048 10908
rect 5048 10852 5104 10908
rect 5104 10852 5108 10908
rect 5044 10848 5108 10852
rect 5124 10908 5188 10912
rect 5124 10852 5128 10908
rect 5128 10852 5184 10908
rect 5184 10852 5188 10908
rect 5124 10848 5188 10852
rect 8817 10908 8881 10912
rect 8817 10852 8821 10908
rect 8821 10852 8877 10908
rect 8877 10852 8881 10908
rect 8817 10848 8881 10852
rect 8897 10908 8961 10912
rect 8897 10852 8901 10908
rect 8901 10852 8957 10908
rect 8957 10852 8961 10908
rect 8897 10848 8961 10852
rect 8977 10908 9041 10912
rect 8977 10852 8981 10908
rect 8981 10852 9037 10908
rect 9037 10852 9041 10908
rect 8977 10848 9041 10852
rect 9057 10908 9121 10912
rect 9057 10852 9061 10908
rect 9061 10852 9117 10908
rect 9117 10852 9121 10908
rect 9057 10848 9121 10852
rect 12750 10908 12814 10912
rect 12750 10852 12754 10908
rect 12754 10852 12810 10908
rect 12810 10852 12814 10908
rect 12750 10848 12814 10852
rect 12830 10908 12894 10912
rect 12830 10852 12834 10908
rect 12834 10852 12890 10908
rect 12890 10852 12894 10908
rect 12830 10848 12894 10852
rect 12910 10908 12974 10912
rect 12910 10852 12914 10908
rect 12914 10852 12970 10908
rect 12970 10852 12974 10908
rect 12910 10848 12974 10852
rect 12990 10908 13054 10912
rect 12990 10852 12994 10908
rect 12994 10852 13050 10908
rect 13050 10852 13054 10908
rect 12990 10848 13054 10852
rect 16683 10908 16747 10912
rect 16683 10852 16687 10908
rect 16687 10852 16743 10908
rect 16743 10852 16747 10908
rect 16683 10848 16747 10852
rect 16763 10908 16827 10912
rect 16763 10852 16767 10908
rect 16767 10852 16823 10908
rect 16823 10852 16827 10908
rect 16763 10848 16827 10852
rect 16843 10908 16907 10912
rect 16843 10852 16847 10908
rect 16847 10852 16903 10908
rect 16903 10852 16907 10908
rect 16843 10848 16907 10852
rect 16923 10908 16987 10912
rect 16923 10852 16927 10908
rect 16927 10852 16983 10908
rect 16983 10852 16987 10908
rect 16923 10848 16987 10852
rect 2918 10364 2982 10368
rect 2918 10308 2922 10364
rect 2922 10308 2978 10364
rect 2978 10308 2982 10364
rect 2918 10304 2982 10308
rect 2998 10364 3062 10368
rect 2998 10308 3002 10364
rect 3002 10308 3058 10364
rect 3058 10308 3062 10364
rect 2998 10304 3062 10308
rect 3078 10364 3142 10368
rect 3078 10308 3082 10364
rect 3082 10308 3138 10364
rect 3138 10308 3142 10364
rect 3078 10304 3142 10308
rect 3158 10364 3222 10368
rect 3158 10308 3162 10364
rect 3162 10308 3218 10364
rect 3218 10308 3222 10364
rect 3158 10304 3222 10308
rect 6851 10364 6915 10368
rect 6851 10308 6855 10364
rect 6855 10308 6911 10364
rect 6911 10308 6915 10364
rect 6851 10304 6915 10308
rect 6931 10364 6995 10368
rect 6931 10308 6935 10364
rect 6935 10308 6991 10364
rect 6991 10308 6995 10364
rect 6931 10304 6995 10308
rect 7011 10364 7075 10368
rect 7011 10308 7015 10364
rect 7015 10308 7071 10364
rect 7071 10308 7075 10364
rect 7011 10304 7075 10308
rect 7091 10364 7155 10368
rect 7091 10308 7095 10364
rect 7095 10308 7151 10364
rect 7151 10308 7155 10364
rect 7091 10304 7155 10308
rect 10784 10364 10848 10368
rect 10784 10308 10788 10364
rect 10788 10308 10844 10364
rect 10844 10308 10848 10364
rect 10784 10304 10848 10308
rect 10864 10364 10928 10368
rect 10864 10308 10868 10364
rect 10868 10308 10924 10364
rect 10924 10308 10928 10364
rect 10864 10304 10928 10308
rect 10944 10364 11008 10368
rect 10944 10308 10948 10364
rect 10948 10308 11004 10364
rect 11004 10308 11008 10364
rect 10944 10304 11008 10308
rect 11024 10364 11088 10368
rect 11024 10308 11028 10364
rect 11028 10308 11084 10364
rect 11084 10308 11088 10364
rect 11024 10304 11088 10308
rect 14717 10364 14781 10368
rect 14717 10308 14721 10364
rect 14721 10308 14777 10364
rect 14777 10308 14781 10364
rect 14717 10304 14781 10308
rect 14797 10364 14861 10368
rect 14797 10308 14801 10364
rect 14801 10308 14857 10364
rect 14857 10308 14861 10364
rect 14797 10304 14861 10308
rect 14877 10364 14941 10368
rect 14877 10308 14881 10364
rect 14881 10308 14937 10364
rect 14937 10308 14941 10364
rect 14877 10304 14941 10308
rect 14957 10364 15021 10368
rect 14957 10308 14961 10364
rect 14961 10308 15017 10364
rect 15017 10308 15021 10364
rect 14957 10304 15021 10308
rect 4884 9820 4948 9824
rect 4884 9764 4888 9820
rect 4888 9764 4944 9820
rect 4944 9764 4948 9820
rect 4884 9760 4948 9764
rect 4964 9820 5028 9824
rect 4964 9764 4968 9820
rect 4968 9764 5024 9820
rect 5024 9764 5028 9820
rect 4964 9760 5028 9764
rect 5044 9820 5108 9824
rect 5044 9764 5048 9820
rect 5048 9764 5104 9820
rect 5104 9764 5108 9820
rect 5044 9760 5108 9764
rect 5124 9820 5188 9824
rect 5124 9764 5128 9820
rect 5128 9764 5184 9820
rect 5184 9764 5188 9820
rect 5124 9760 5188 9764
rect 8817 9820 8881 9824
rect 8817 9764 8821 9820
rect 8821 9764 8877 9820
rect 8877 9764 8881 9820
rect 8817 9760 8881 9764
rect 8897 9820 8961 9824
rect 8897 9764 8901 9820
rect 8901 9764 8957 9820
rect 8957 9764 8961 9820
rect 8897 9760 8961 9764
rect 8977 9820 9041 9824
rect 8977 9764 8981 9820
rect 8981 9764 9037 9820
rect 9037 9764 9041 9820
rect 8977 9760 9041 9764
rect 9057 9820 9121 9824
rect 9057 9764 9061 9820
rect 9061 9764 9117 9820
rect 9117 9764 9121 9820
rect 9057 9760 9121 9764
rect 12750 9820 12814 9824
rect 12750 9764 12754 9820
rect 12754 9764 12810 9820
rect 12810 9764 12814 9820
rect 12750 9760 12814 9764
rect 12830 9820 12894 9824
rect 12830 9764 12834 9820
rect 12834 9764 12890 9820
rect 12890 9764 12894 9820
rect 12830 9760 12894 9764
rect 12910 9820 12974 9824
rect 12910 9764 12914 9820
rect 12914 9764 12970 9820
rect 12970 9764 12974 9820
rect 12910 9760 12974 9764
rect 12990 9820 13054 9824
rect 12990 9764 12994 9820
rect 12994 9764 13050 9820
rect 13050 9764 13054 9820
rect 12990 9760 13054 9764
rect 16683 9820 16747 9824
rect 16683 9764 16687 9820
rect 16687 9764 16743 9820
rect 16743 9764 16747 9820
rect 16683 9760 16747 9764
rect 16763 9820 16827 9824
rect 16763 9764 16767 9820
rect 16767 9764 16823 9820
rect 16823 9764 16827 9820
rect 16763 9760 16827 9764
rect 16843 9820 16907 9824
rect 16843 9764 16847 9820
rect 16847 9764 16903 9820
rect 16903 9764 16907 9820
rect 16843 9760 16907 9764
rect 16923 9820 16987 9824
rect 16923 9764 16927 9820
rect 16927 9764 16983 9820
rect 16983 9764 16987 9820
rect 16923 9760 16987 9764
rect 3372 9692 3436 9756
rect 2918 9276 2982 9280
rect 2918 9220 2922 9276
rect 2922 9220 2978 9276
rect 2978 9220 2982 9276
rect 2918 9216 2982 9220
rect 2998 9276 3062 9280
rect 2998 9220 3002 9276
rect 3002 9220 3058 9276
rect 3058 9220 3062 9276
rect 2998 9216 3062 9220
rect 3078 9276 3142 9280
rect 3078 9220 3082 9276
rect 3082 9220 3138 9276
rect 3138 9220 3142 9276
rect 3078 9216 3142 9220
rect 3158 9276 3222 9280
rect 3158 9220 3162 9276
rect 3162 9220 3218 9276
rect 3218 9220 3222 9276
rect 3158 9216 3222 9220
rect 6851 9276 6915 9280
rect 6851 9220 6855 9276
rect 6855 9220 6911 9276
rect 6911 9220 6915 9276
rect 6851 9216 6915 9220
rect 6931 9276 6995 9280
rect 6931 9220 6935 9276
rect 6935 9220 6991 9276
rect 6991 9220 6995 9276
rect 6931 9216 6995 9220
rect 7011 9276 7075 9280
rect 7011 9220 7015 9276
rect 7015 9220 7071 9276
rect 7071 9220 7075 9276
rect 7011 9216 7075 9220
rect 7091 9276 7155 9280
rect 7091 9220 7095 9276
rect 7095 9220 7151 9276
rect 7151 9220 7155 9276
rect 7091 9216 7155 9220
rect 10784 9276 10848 9280
rect 10784 9220 10788 9276
rect 10788 9220 10844 9276
rect 10844 9220 10848 9276
rect 10784 9216 10848 9220
rect 10864 9276 10928 9280
rect 10864 9220 10868 9276
rect 10868 9220 10924 9276
rect 10924 9220 10928 9276
rect 10864 9216 10928 9220
rect 10944 9276 11008 9280
rect 10944 9220 10948 9276
rect 10948 9220 11004 9276
rect 11004 9220 11008 9276
rect 10944 9216 11008 9220
rect 11024 9276 11088 9280
rect 11024 9220 11028 9276
rect 11028 9220 11084 9276
rect 11084 9220 11088 9276
rect 11024 9216 11088 9220
rect 14717 9276 14781 9280
rect 14717 9220 14721 9276
rect 14721 9220 14777 9276
rect 14777 9220 14781 9276
rect 14717 9216 14781 9220
rect 14797 9276 14861 9280
rect 14797 9220 14801 9276
rect 14801 9220 14857 9276
rect 14857 9220 14861 9276
rect 14797 9216 14861 9220
rect 14877 9276 14941 9280
rect 14877 9220 14881 9276
rect 14881 9220 14937 9276
rect 14937 9220 14941 9276
rect 14877 9216 14941 9220
rect 14957 9276 15021 9280
rect 14957 9220 14961 9276
rect 14961 9220 15017 9276
rect 15017 9220 15021 9276
rect 14957 9216 15021 9220
rect 4884 8732 4948 8736
rect 4884 8676 4888 8732
rect 4888 8676 4944 8732
rect 4944 8676 4948 8732
rect 4884 8672 4948 8676
rect 4964 8732 5028 8736
rect 4964 8676 4968 8732
rect 4968 8676 5024 8732
rect 5024 8676 5028 8732
rect 4964 8672 5028 8676
rect 5044 8732 5108 8736
rect 5044 8676 5048 8732
rect 5048 8676 5104 8732
rect 5104 8676 5108 8732
rect 5044 8672 5108 8676
rect 5124 8732 5188 8736
rect 5124 8676 5128 8732
rect 5128 8676 5184 8732
rect 5184 8676 5188 8732
rect 5124 8672 5188 8676
rect 8817 8732 8881 8736
rect 8817 8676 8821 8732
rect 8821 8676 8877 8732
rect 8877 8676 8881 8732
rect 8817 8672 8881 8676
rect 8897 8732 8961 8736
rect 8897 8676 8901 8732
rect 8901 8676 8957 8732
rect 8957 8676 8961 8732
rect 8897 8672 8961 8676
rect 8977 8732 9041 8736
rect 8977 8676 8981 8732
rect 8981 8676 9037 8732
rect 9037 8676 9041 8732
rect 8977 8672 9041 8676
rect 9057 8732 9121 8736
rect 9057 8676 9061 8732
rect 9061 8676 9117 8732
rect 9117 8676 9121 8732
rect 9057 8672 9121 8676
rect 12750 8732 12814 8736
rect 12750 8676 12754 8732
rect 12754 8676 12810 8732
rect 12810 8676 12814 8732
rect 12750 8672 12814 8676
rect 12830 8732 12894 8736
rect 12830 8676 12834 8732
rect 12834 8676 12890 8732
rect 12890 8676 12894 8732
rect 12830 8672 12894 8676
rect 12910 8732 12974 8736
rect 12910 8676 12914 8732
rect 12914 8676 12970 8732
rect 12970 8676 12974 8732
rect 12910 8672 12974 8676
rect 12990 8732 13054 8736
rect 12990 8676 12994 8732
rect 12994 8676 13050 8732
rect 13050 8676 13054 8732
rect 12990 8672 13054 8676
rect 16683 8732 16747 8736
rect 16683 8676 16687 8732
rect 16687 8676 16743 8732
rect 16743 8676 16747 8732
rect 16683 8672 16747 8676
rect 16763 8732 16827 8736
rect 16763 8676 16767 8732
rect 16767 8676 16823 8732
rect 16823 8676 16827 8732
rect 16763 8672 16827 8676
rect 16843 8732 16907 8736
rect 16843 8676 16847 8732
rect 16847 8676 16903 8732
rect 16903 8676 16907 8732
rect 16843 8672 16907 8676
rect 16923 8732 16987 8736
rect 16923 8676 16927 8732
rect 16927 8676 16983 8732
rect 16983 8676 16987 8732
rect 16923 8672 16987 8676
rect 2918 8188 2982 8192
rect 2918 8132 2922 8188
rect 2922 8132 2978 8188
rect 2978 8132 2982 8188
rect 2918 8128 2982 8132
rect 2998 8188 3062 8192
rect 2998 8132 3002 8188
rect 3002 8132 3058 8188
rect 3058 8132 3062 8188
rect 2998 8128 3062 8132
rect 3078 8188 3142 8192
rect 3078 8132 3082 8188
rect 3082 8132 3138 8188
rect 3138 8132 3142 8188
rect 3078 8128 3142 8132
rect 3158 8188 3222 8192
rect 3158 8132 3162 8188
rect 3162 8132 3218 8188
rect 3218 8132 3222 8188
rect 3158 8128 3222 8132
rect 6851 8188 6915 8192
rect 6851 8132 6855 8188
rect 6855 8132 6911 8188
rect 6911 8132 6915 8188
rect 6851 8128 6915 8132
rect 6931 8188 6995 8192
rect 6931 8132 6935 8188
rect 6935 8132 6991 8188
rect 6991 8132 6995 8188
rect 6931 8128 6995 8132
rect 7011 8188 7075 8192
rect 7011 8132 7015 8188
rect 7015 8132 7071 8188
rect 7071 8132 7075 8188
rect 7011 8128 7075 8132
rect 7091 8188 7155 8192
rect 7091 8132 7095 8188
rect 7095 8132 7151 8188
rect 7151 8132 7155 8188
rect 7091 8128 7155 8132
rect 10784 8188 10848 8192
rect 10784 8132 10788 8188
rect 10788 8132 10844 8188
rect 10844 8132 10848 8188
rect 10784 8128 10848 8132
rect 10864 8188 10928 8192
rect 10864 8132 10868 8188
rect 10868 8132 10924 8188
rect 10924 8132 10928 8188
rect 10864 8128 10928 8132
rect 10944 8188 11008 8192
rect 10944 8132 10948 8188
rect 10948 8132 11004 8188
rect 11004 8132 11008 8188
rect 10944 8128 11008 8132
rect 11024 8188 11088 8192
rect 11024 8132 11028 8188
rect 11028 8132 11084 8188
rect 11084 8132 11088 8188
rect 11024 8128 11088 8132
rect 14717 8188 14781 8192
rect 14717 8132 14721 8188
rect 14721 8132 14777 8188
rect 14777 8132 14781 8188
rect 14717 8128 14781 8132
rect 14797 8188 14861 8192
rect 14797 8132 14801 8188
rect 14801 8132 14857 8188
rect 14857 8132 14861 8188
rect 14797 8128 14861 8132
rect 14877 8188 14941 8192
rect 14877 8132 14881 8188
rect 14881 8132 14937 8188
rect 14937 8132 14941 8188
rect 14877 8128 14941 8132
rect 14957 8188 15021 8192
rect 14957 8132 14961 8188
rect 14961 8132 15017 8188
rect 15017 8132 15021 8188
rect 14957 8128 15021 8132
rect 4884 7644 4948 7648
rect 4884 7588 4888 7644
rect 4888 7588 4944 7644
rect 4944 7588 4948 7644
rect 4884 7584 4948 7588
rect 4964 7644 5028 7648
rect 4964 7588 4968 7644
rect 4968 7588 5024 7644
rect 5024 7588 5028 7644
rect 4964 7584 5028 7588
rect 5044 7644 5108 7648
rect 5044 7588 5048 7644
rect 5048 7588 5104 7644
rect 5104 7588 5108 7644
rect 5044 7584 5108 7588
rect 5124 7644 5188 7648
rect 5124 7588 5128 7644
rect 5128 7588 5184 7644
rect 5184 7588 5188 7644
rect 5124 7584 5188 7588
rect 8817 7644 8881 7648
rect 8817 7588 8821 7644
rect 8821 7588 8877 7644
rect 8877 7588 8881 7644
rect 8817 7584 8881 7588
rect 8897 7644 8961 7648
rect 8897 7588 8901 7644
rect 8901 7588 8957 7644
rect 8957 7588 8961 7644
rect 8897 7584 8961 7588
rect 8977 7644 9041 7648
rect 8977 7588 8981 7644
rect 8981 7588 9037 7644
rect 9037 7588 9041 7644
rect 8977 7584 9041 7588
rect 9057 7644 9121 7648
rect 9057 7588 9061 7644
rect 9061 7588 9117 7644
rect 9117 7588 9121 7644
rect 9057 7584 9121 7588
rect 12750 7644 12814 7648
rect 12750 7588 12754 7644
rect 12754 7588 12810 7644
rect 12810 7588 12814 7644
rect 12750 7584 12814 7588
rect 12830 7644 12894 7648
rect 12830 7588 12834 7644
rect 12834 7588 12890 7644
rect 12890 7588 12894 7644
rect 12830 7584 12894 7588
rect 12910 7644 12974 7648
rect 12910 7588 12914 7644
rect 12914 7588 12970 7644
rect 12970 7588 12974 7644
rect 12910 7584 12974 7588
rect 12990 7644 13054 7648
rect 12990 7588 12994 7644
rect 12994 7588 13050 7644
rect 13050 7588 13054 7644
rect 12990 7584 13054 7588
rect 16683 7644 16747 7648
rect 16683 7588 16687 7644
rect 16687 7588 16743 7644
rect 16743 7588 16747 7644
rect 16683 7584 16747 7588
rect 16763 7644 16827 7648
rect 16763 7588 16767 7644
rect 16767 7588 16823 7644
rect 16823 7588 16827 7644
rect 16763 7584 16827 7588
rect 16843 7644 16907 7648
rect 16843 7588 16847 7644
rect 16847 7588 16903 7644
rect 16903 7588 16907 7644
rect 16843 7584 16907 7588
rect 16923 7644 16987 7648
rect 16923 7588 16927 7644
rect 16927 7588 16983 7644
rect 16983 7588 16987 7644
rect 16923 7584 16987 7588
rect 2918 7100 2982 7104
rect 2918 7044 2922 7100
rect 2922 7044 2978 7100
rect 2978 7044 2982 7100
rect 2918 7040 2982 7044
rect 2998 7100 3062 7104
rect 2998 7044 3002 7100
rect 3002 7044 3058 7100
rect 3058 7044 3062 7100
rect 2998 7040 3062 7044
rect 3078 7100 3142 7104
rect 3078 7044 3082 7100
rect 3082 7044 3138 7100
rect 3138 7044 3142 7100
rect 3078 7040 3142 7044
rect 3158 7100 3222 7104
rect 3158 7044 3162 7100
rect 3162 7044 3218 7100
rect 3218 7044 3222 7100
rect 3158 7040 3222 7044
rect 6851 7100 6915 7104
rect 6851 7044 6855 7100
rect 6855 7044 6911 7100
rect 6911 7044 6915 7100
rect 6851 7040 6915 7044
rect 6931 7100 6995 7104
rect 6931 7044 6935 7100
rect 6935 7044 6991 7100
rect 6991 7044 6995 7100
rect 6931 7040 6995 7044
rect 7011 7100 7075 7104
rect 7011 7044 7015 7100
rect 7015 7044 7071 7100
rect 7071 7044 7075 7100
rect 7011 7040 7075 7044
rect 7091 7100 7155 7104
rect 7091 7044 7095 7100
rect 7095 7044 7151 7100
rect 7151 7044 7155 7100
rect 7091 7040 7155 7044
rect 10784 7100 10848 7104
rect 10784 7044 10788 7100
rect 10788 7044 10844 7100
rect 10844 7044 10848 7100
rect 10784 7040 10848 7044
rect 10864 7100 10928 7104
rect 10864 7044 10868 7100
rect 10868 7044 10924 7100
rect 10924 7044 10928 7100
rect 10864 7040 10928 7044
rect 10944 7100 11008 7104
rect 10944 7044 10948 7100
rect 10948 7044 11004 7100
rect 11004 7044 11008 7100
rect 10944 7040 11008 7044
rect 11024 7100 11088 7104
rect 11024 7044 11028 7100
rect 11028 7044 11084 7100
rect 11084 7044 11088 7100
rect 11024 7040 11088 7044
rect 14717 7100 14781 7104
rect 14717 7044 14721 7100
rect 14721 7044 14777 7100
rect 14777 7044 14781 7100
rect 14717 7040 14781 7044
rect 14797 7100 14861 7104
rect 14797 7044 14801 7100
rect 14801 7044 14857 7100
rect 14857 7044 14861 7100
rect 14797 7040 14861 7044
rect 14877 7100 14941 7104
rect 14877 7044 14881 7100
rect 14881 7044 14937 7100
rect 14937 7044 14941 7100
rect 14877 7040 14941 7044
rect 14957 7100 15021 7104
rect 14957 7044 14961 7100
rect 14961 7044 15017 7100
rect 15017 7044 15021 7100
rect 14957 7040 15021 7044
rect 4884 6556 4948 6560
rect 4884 6500 4888 6556
rect 4888 6500 4944 6556
rect 4944 6500 4948 6556
rect 4884 6496 4948 6500
rect 4964 6556 5028 6560
rect 4964 6500 4968 6556
rect 4968 6500 5024 6556
rect 5024 6500 5028 6556
rect 4964 6496 5028 6500
rect 5044 6556 5108 6560
rect 5044 6500 5048 6556
rect 5048 6500 5104 6556
rect 5104 6500 5108 6556
rect 5044 6496 5108 6500
rect 5124 6556 5188 6560
rect 5124 6500 5128 6556
rect 5128 6500 5184 6556
rect 5184 6500 5188 6556
rect 5124 6496 5188 6500
rect 8817 6556 8881 6560
rect 8817 6500 8821 6556
rect 8821 6500 8877 6556
rect 8877 6500 8881 6556
rect 8817 6496 8881 6500
rect 8897 6556 8961 6560
rect 8897 6500 8901 6556
rect 8901 6500 8957 6556
rect 8957 6500 8961 6556
rect 8897 6496 8961 6500
rect 8977 6556 9041 6560
rect 8977 6500 8981 6556
rect 8981 6500 9037 6556
rect 9037 6500 9041 6556
rect 8977 6496 9041 6500
rect 9057 6556 9121 6560
rect 9057 6500 9061 6556
rect 9061 6500 9117 6556
rect 9117 6500 9121 6556
rect 9057 6496 9121 6500
rect 12750 6556 12814 6560
rect 12750 6500 12754 6556
rect 12754 6500 12810 6556
rect 12810 6500 12814 6556
rect 12750 6496 12814 6500
rect 12830 6556 12894 6560
rect 12830 6500 12834 6556
rect 12834 6500 12890 6556
rect 12890 6500 12894 6556
rect 12830 6496 12894 6500
rect 12910 6556 12974 6560
rect 12910 6500 12914 6556
rect 12914 6500 12970 6556
rect 12970 6500 12974 6556
rect 12910 6496 12974 6500
rect 12990 6556 13054 6560
rect 12990 6500 12994 6556
rect 12994 6500 13050 6556
rect 13050 6500 13054 6556
rect 12990 6496 13054 6500
rect 16683 6556 16747 6560
rect 16683 6500 16687 6556
rect 16687 6500 16743 6556
rect 16743 6500 16747 6556
rect 16683 6496 16747 6500
rect 16763 6556 16827 6560
rect 16763 6500 16767 6556
rect 16767 6500 16823 6556
rect 16823 6500 16827 6556
rect 16763 6496 16827 6500
rect 16843 6556 16907 6560
rect 16843 6500 16847 6556
rect 16847 6500 16903 6556
rect 16903 6500 16907 6556
rect 16843 6496 16907 6500
rect 16923 6556 16987 6560
rect 16923 6500 16927 6556
rect 16927 6500 16983 6556
rect 16983 6500 16987 6556
rect 16923 6496 16987 6500
rect 2918 6012 2982 6016
rect 2918 5956 2922 6012
rect 2922 5956 2978 6012
rect 2978 5956 2982 6012
rect 2918 5952 2982 5956
rect 2998 6012 3062 6016
rect 2998 5956 3002 6012
rect 3002 5956 3058 6012
rect 3058 5956 3062 6012
rect 2998 5952 3062 5956
rect 3078 6012 3142 6016
rect 3078 5956 3082 6012
rect 3082 5956 3138 6012
rect 3138 5956 3142 6012
rect 3078 5952 3142 5956
rect 3158 6012 3222 6016
rect 3158 5956 3162 6012
rect 3162 5956 3218 6012
rect 3218 5956 3222 6012
rect 3158 5952 3222 5956
rect 6851 6012 6915 6016
rect 6851 5956 6855 6012
rect 6855 5956 6911 6012
rect 6911 5956 6915 6012
rect 6851 5952 6915 5956
rect 6931 6012 6995 6016
rect 6931 5956 6935 6012
rect 6935 5956 6991 6012
rect 6991 5956 6995 6012
rect 6931 5952 6995 5956
rect 7011 6012 7075 6016
rect 7011 5956 7015 6012
rect 7015 5956 7071 6012
rect 7071 5956 7075 6012
rect 7011 5952 7075 5956
rect 7091 6012 7155 6016
rect 7091 5956 7095 6012
rect 7095 5956 7151 6012
rect 7151 5956 7155 6012
rect 7091 5952 7155 5956
rect 10784 6012 10848 6016
rect 10784 5956 10788 6012
rect 10788 5956 10844 6012
rect 10844 5956 10848 6012
rect 10784 5952 10848 5956
rect 10864 6012 10928 6016
rect 10864 5956 10868 6012
rect 10868 5956 10924 6012
rect 10924 5956 10928 6012
rect 10864 5952 10928 5956
rect 10944 6012 11008 6016
rect 10944 5956 10948 6012
rect 10948 5956 11004 6012
rect 11004 5956 11008 6012
rect 10944 5952 11008 5956
rect 11024 6012 11088 6016
rect 11024 5956 11028 6012
rect 11028 5956 11084 6012
rect 11084 5956 11088 6012
rect 11024 5952 11088 5956
rect 14717 6012 14781 6016
rect 14717 5956 14721 6012
rect 14721 5956 14777 6012
rect 14777 5956 14781 6012
rect 14717 5952 14781 5956
rect 14797 6012 14861 6016
rect 14797 5956 14801 6012
rect 14801 5956 14857 6012
rect 14857 5956 14861 6012
rect 14797 5952 14861 5956
rect 14877 6012 14941 6016
rect 14877 5956 14881 6012
rect 14881 5956 14937 6012
rect 14937 5956 14941 6012
rect 14877 5952 14941 5956
rect 14957 6012 15021 6016
rect 14957 5956 14961 6012
rect 14961 5956 15017 6012
rect 15017 5956 15021 6012
rect 14957 5952 15021 5956
rect 4884 5468 4948 5472
rect 4884 5412 4888 5468
rect 4888 5412 4944 5468
rect 4944 5412 4948 5468
rect 4884 5408 4948 5412
rect 4964 5468 5028 5472
rect 4964 5412 4968 5468
rect 4968 5412 5024 5468
rect 5024 5412 5028 5468
rect 4964 5408 5028 5412
rect 5044 5468 5108 5472
rect 5044 5412 5048 5468
rect 5048 5412 5104 5468
rect 5104 5412 5108 5468
rect 5044 5408 5108 5412
rect 5124 5468 5188 5472
rect 5124 5412 5128 5468
rect 5128 5412 5184 5468
rect 5184 5412 5188 5468
rect 5124 5408 5188 5412
rect 8817 5468 8881 5472
rect 8817 5412 8821 5468
rect 8821 5412 8877 5468
rect 8877 5412 8881 5468
rect 8817 5408 8881 5412
rect 8897 5468 8961 5472
rect 8897 5412 8901 5468
rect 8901 5412 8957 5468
rect 8957 5412 8961 5468
rect 8897 5408 8961 5412
rect 8977 5468 9041 5472
rect 8977 5412 8981 5468
rect 8981 5412 9037 5468
rect 9037 5412 9041 5468
rect 8977 5408 9041 5412
rect 9057 5468 9121 5472
rect 9057 5412 9061 5468
rect 9061 5412 9117 5468
rect 9117 5412 9121 5468
rect 9057 5408 9121 5412
rect 12750 5468 12814 5472
rect 12750 5412 12754 5468
rect 12754 5412 12810 5468
rect 12810 5412 12814 5468
rect 12750 5408 12814 5412
rect 12830 5468 12894 5472
rect 12830 5412 12834 5468
rect 12834 5412 12890 5468
rect 12890 5412 12894 5468
rect 12830 5408 12894 5412
rect 12910 5468 12974 5472
rect 12910 5412 12914 5468
rect 12914 5412 12970 5468
rect 12970 5412 12974 5468
rect 12910 5408 12974 5412
rect 12990 5468 13054 5472
rect 12990 5412 12994 5468
rect 12994 5412 13050 5468
rect 13050 5412 13054 5468
rect 12990 5408 13054 5412
rect 16683 5468 16747 5472
rect 16683 5412 16687 5468
rect 16687 5412 16743 5468
rect 16743 5412 16747 5468
rect 16683 5408 16747 5412
rect 16763 5468 16827 5472
rect 16763 5412 16767 5468
rect 16767 5412 16823 5468
rect 16823 5412 16827 5468
rect 16763 5408 16827 5412
rect 16843 5468 16907 5472
rect 16843 5412 16847 5468
rect 16847 5412 16903 5468
rect 16903 5412 16907 5468
rect 16843 5408 16907 5412
rect 16923 5468 16987 5472
rect 16923 5412 16927 5468
rect 16927 5412 16983 5468
rect 16983 5412 16987 5468
rect 16923 5408 16987 5412
rect 2918 4924 2982 4928
rect 2918 4868 2922 4924
rect 2922 4868 2978 4924
rect 2978 4868 2982 4924
rect 2918 4864 2982 4868
rect 2998 4924 3062 4928
rect 2998 4868 3002 4924
rect 3002 4868 3058 4924
rect 3058 4868 3062 4924
rect 2998 4864 3062 4868
rect 3078 4924 3142 4928
rect 3078 4868 3082 4924
rect 3082 4868 3138 4924
rect 3138 4868 3142 4924
rect 3078 4864 3142 4868
rect 3158 4924 3222 4928
rect 3158 4868 3162 4924
rect 3162 4868 3218 4924
rect 3218 4868 3222 4924
rect 3158 4864 3222 4868
rect 6851 4924 6915 4928
rect 6851 4868 6855 4924
rect 6855 4868 6911 4924
rect 6911 4868 6915 4924
rect 6851 4864 6915 4868
rect 6931 4924 6995 4928
rect 6931 4868 6935 4924
rect 6935 4868 6991 4924
rect 6991 4868 6995 4924
rect 6931 4864 6995 4868
rect 7011 4924 7075 4928
rect 7011 4868 7015 4924
rect 7015 4868 7071 4924
rect 7071 4868 7075 4924
rect 7011 4864 7075 4868
rect 7091 4924 7155 4928
rect 7091 4868 7095 4924
rect 7095 4868 7151 4924
rect 7151 4868 7155 4924
rect 7091 4864 7155 4868
rect 10784 4924 10848 4928
rect 10784 4868 10788 4924
rect 10788 4868 10844 4924
rect 10844 4868 10848 4924
rect 10784 4864 10848 4868
rect 10864 4924 10928 4928
rect 10864 4868 10868 4924
rect 10868 4868 10924 4924
rect 10924 4868 10928 4924
rect 10864 4864 10928 4868
rect 10944 4924 11008 4928
rect 10944 4868 10948 4924
rect 10948 4868 11004 4924
rect 11004 4868 11008 4924
rect 10944 4864 11008 4868
rect 11024 4924 11088 4928
rect 11024 4868 11028 4924
rect 11028 4868 11084 4924
rect 11084 4868 11088 4924
rect 11024 4864 11088 4868
rect 14717 4924 14781 4928
rect 14717 4868 14721 4924
rect 14721 4868 14777 4924
rect 14777 4868 14781 4924
rect 14717 4864 14781 4868
rect 14797 4924 14861 4928
rect 14797 4868 14801 4924
rect 14801 4868 14857 4924
rect 14857 4868 14861 4924
rect 14797 4864 14861 4868
rect 14877 4924 14941 4928
rect 14877 4868 14881 4924
rect 14881 4868 14937 4924
rect 14937 4868 14941 4924
rect 14877 4864 14941 4868
rect 14957 4924 15021 4928
rect 14957 4868 14961 4924
rect 14961 4868 15017 4924
rect 15017 4868 15021 4924
rect 14957 4864 15021 4868
rect 4884 4380 4948 4384
rect 4884 4324 4888 4380
rect 4888 4324 4944 4380
rect 4944 4324 4948 4380
rect 4884 4320 4948 4324
rect 4964 4380 5028 4384
rect 4964 4324 4968 4380
rect 4968 4324 5024 4380
rect 5024 4324 5028 4380
rect 4964 4320 5028 4324
rect 5044 4380 5108 4384
rect 5044 4324 5048 4380
rect 5048 4324 5104 4380
rect 5104 4324 5108 4380
rect 5044 4320 5108 4324
rect 5124 4380 5188 4384
rect 5124 4324 5128 4380
rect 5128 4324 5184 4380
rect 5184 4324 5188 4380
rect 5124 4320 5188 4324
rect 8817 4380 8881 4384
rect 8817 4324 8821 4380
rect 8821 4324 8877 4380
rect 8877 4324 8881 4380
rect 8817 4320 8881 4324
rect 8897 4380 8961 4384
rect 8897 4324 8901 4380
rect 8901 4324 8957 4380
rect 8957 4324 8961 4380
rect 8897 4320 8961 4324
rect 8977 4380 9041 4384
rect 8977 4324 8981 4380
rect 8981 4324 9037 4380
rect 9037 4324 9041 4380
rect 8977 4320 9041 4324
rect 9057 4380 9121 4384
rect 9057 4324 9061 4380
rect 9061 4324 9117 4380
rect 9117 4324 9121 4380
rect 9057 4320 9121 4324
rect 12750 4380 12814 4384
rect 12750 4324 12754 4380
rect 12754 4324 12810 4380
rect 12810 4324 12814 4380
rect 12750 4320 12814 4324
rect 12830 4380 12894 4384
rect 12830 4324 12834 4380
rect 12834 4324 12890 4380
rect 12890 4324 12894 4380
rect 12830 4320 12894 4324
rect 12910 4380 12974 4384
rect 12910 4324 12914 4380
rect 12914 4324 12970 4380
rect 12970 4324 12974 4380
rect 12910 4320 12974 4324
rect 12990 4380 13054 4384
rect 12990 4324 12994 4380
rect 12994 4324 13050 4380
rect 13050 4324 13054 4380
rect 12990 4320 13054 4324
rect 16683 4380 16747 4384
rect 16683 4324 16687 4380
rect 16687 4324 16743 4380
rect 16743 4324 16747 4380
rect 16683 4320 16747 4324
rect 16763 4380 16827 4384
rect 16763 4324 16767 4380
rect 16767 4324 16823 4380
rect 16823 4324 16827 4380
rect 16763 4320 16827 4324
rect 16843 4380 16907 4384
rect 16843 4324 16847 4380
rect 16847 4324 16903 4380
rect 16903 4324 16907 4380
rect 16843 4320 16907 4324
rect 16923 4380 16987 4384
rect 16923 4324 16927 4380
rect 16927 4324 16983 4380
rect 16983 4324 16987 4380
rect 16923 4320 16987 4324
rect 3372 3980 3436 4044
rect 2918 3836 2982 3840
rect 2918 3780 2922 3836
rect 2922 3780 2978 3836
rect 2978 3780 2982 3836
rect 2918 3776 2982 3780
rect 2998 3836 3062 3840
rect 2998 3780 3002 3836
rect 3002 3780 3058 3836
rect 3058 3780 3062 3836
rect 2998 3776 3062 3780
rect 3078 3836 3142 3840
rect 3078 3780 3082 3836
rect 3082 3780 3138 3836
rect 3138 3780 3142 3836
rect 3078 3776 3142 3780
rect 3158 3836 3222 3840
rect 3158 3780 3162 3836
rect 3162 3780 3218 3836
rect 3218 3780 3222 3836
rect 3158 3776 3222 3780
rect 6851 3836 6915 3840
rect 6851 3780 6855 3836
rect 6855 3780 6911 3836
rect 6911 3780 6915 3836
rect 6851 3776 6915 3780
rect 6931 3836 6995 3840
rect 6931 3780 6935 3836
rect 6935 3780 6991 3836
rect 6991 3780 6995 3836
rect 6931 3776 6995 3780
rect 7011 3836 7075 3840
rect 7011 3780 7015 3836
rect 7015 3780 7071 3836
rect 7071 3780 7075 3836
rect 7011 3776 7075 3780
rect 7091 3836 7155 3840
rect 7091 3780 7095 3836
rect 7095 3780 7151 3836
rect 7151 3780 7155 3836
rect 7091 3776 7155 3780
rect 10784 3836 10848 3840
rect 10784 3780 10788 3836
rect 10788 3780 10844 3836
rect 10844 3780 10848 3836
rect 10784 3776 10848 3780
rect 10864 3836 10928 3840
rect 10864 3780 10868 3836
rect 10868 3780 10924 3836
rect 10924 3780 10928 3836
rect 10864 3776 10928 3780
rect 10944 3836 11008 3840
rect 10944 3780 10948 3836
rect 10948 3780 11004 3836
rect 11004 3780 11008 3836
rect 10944 3776 11008 3780
rect 11024 3836 11088 3840
rect 11024 3780 11028 3836
rect 11028 3780 11084 3836
rect 11084 3780 11088 3836
rect 11024 3776 11088 3780
rect 14717 3836 14781 3840
rect 14717 3780 14721 3836
rect 14721 3780 14777 3836
rect 14777 3780 14781 3836
rect 14717 3776 14781 3780
rect 14797 3836 14861 3840
rect 14797 3780 14801 3836
rect 14801 3780 14857 3836
rect 14857 3780 14861 3836
rect 14797 3776 14861 3780
rect 14877 3836 14941 3840
rect 14877 3780 14881 3836
rect 14881 3780 14937 3836
rect 14937 3780 14941 3836
rect 14877 3776 14941 3780
rect 14957 3836 15021 3840
rect 14957 3780 14961 3836
rect 14961 3780 15017 3836
rect 15017 3780 15021 3836
rect 14957 3776 15021 3780
rect 4884 3292 4948 3296
rect 4884 3236 4888 3292
rect 4888 3236 4944 3292
rect 4944 3236 4948 3292
rect 4884 3232 4948 3236
rect 4964 3292 5028 3296
rect 4964 3236 4968 3292
rect 4968 3236 5024 3292
rect 5024 3236 5028 3292
rect 4964 3232 5028 3236
rect 5044 3292 5108 3296
rect 5044 3236 5048 3292
rect 5048 3236 5104 3292
rect 5104 3236 5108 3292
rect 5044 3232 5108 3236
rect 5124 3292 5188 3296
rect 5124 3236 5128 3292
rect 5128 3236 5184 3292
rect 5184 3236 5188 3292
rect 5124 3232 5188 3236
rect 8817 3292 8881 3296
rect 8817 3236 8821 3292
rect 8821 3236 8877 3292
rect 8877 3236 8881 3292
rect 8817 3232 8881 3236
rect 8897 3292 8961 3296
rect 8897 3236 8901 3292
rect 8901 3236 8957 3292
rect 8957 3236 8961 3292
rect 8897 3232 8961 3236
rect 8977 3292 9041 3296
rect 8977 3236 8981 3292
rect 8981 3236 9037 3292
rect 9037 3236 9041 3292
rect 8977 3232 9041 3236
rect 9057 3292 9121 3296
rect 9057 3236 9061 3292
rect 9061 3236 9117 3292
rect 9117 3236 9121 3292
rect 9057 3232 9121 3236
rect 12750 3292 12814 3296
rect 12750 3236 12754 3292
rect 12754 3236 12810 3292
rect 12810 3236 12814 3292
rect 12750 3232 12814 3236
rect 12830 3292 12894 3296
rect 12830 3236 12834 3292
rect 12834 3236 12890 3292
rect 12890 3236 12894 3292
rect 12830 3232 12894 3236
rect 12910 3292 12974 3296
rect 12910 3236 12914 3292
rect 12914 3236 12970 3292
rect 12970 3236 12974 3292
rect 12910 3232 12974 3236
rect 12990 3292 13054 3296
rect 12990 3236 12994 3292
rect 12994 3236 13050 3292
rect 13050 3236 13054 3292
rect 12990 3232 13054 3236
rect 16683 3292 16747 3296
rect 16683 3236 16687 3292
rect 16687 3236 16743 3292
rect 16743 3236 16747 3292
rect 16683 3232 16747 3236
rect 16763 3292 16827 3296
rect 16763 3236 16767 3292
rect 16767 3236 16823 3292
rect 16823 3236 16827 3292
rect 16763 3232 16827 3236
rect 16843 3292 16907 3296
rect 16843 3236 16847 3292
rect 16847 3236 16903 3292
rect 16903 3236 16907 3292
rect 16843 3232 16907 3236
rect 16923 3292 16987 3296
rect 16923 3236 16927 3292
rect 16927 3236 16983 3292
rect 16983 3236 16987 3292
rect 16923 3232 16987 3236
rect 2918 2748 2982 2752
rect 2918 2692 2922 2748
rect 2922 2692 2978 2748
rect 2978 2692 2982 2748
rect 2918 2688 2982 2692
rect 2998 2748 3062 2752
rect 2998 2692 3002 2748
rect 3002 2692 3058 2748
rect 3058 2692 3062 2748
rect 2998 2688 3062 2692
rect 3078 2748 3142 2752
rect 3078 2692 3082 2748
rect 3082 2692 3138 2748
rect 3138 2692 3142 2748
rect 3078 2688 3142 2692
rect 3158 2748 3222 2752
rect 3158 2692 3162 2748
rect 3162 2692 3218 2748
rect 3218 2692 3222 2748
rect 3158 2688 3222 2692
rect 6851 2748 6915 2752
rect 6851 2692 6855 2748
rect 6855 2692 6911 2748
rect 6911 2692 6915 2748
rect 6851 2688 6915 2692
rect 6931 2748 6995 2752
rect 6931 2692 6935 2748
rect 6935 2692 6991 2748
rect 6991 2692 6995 2748
rect 6931 2688 6995 2692
rect 7011 2748 7075 2752
rect 7011 2692 7015 2748
rect 7015 2692 7071 2748
rect 7071 2692 7075 2748
rect 7011 2688 7075 2692
rect 7091 2748 7155 2752
rect 7091 2692 7095 2748
rect 7095 2692 7151 2748
rect 7151 2692 7155 2748
rect 7091 2688 7155 2692
rect 10784 2748 10848 2752
rect 10784 2692 10788 2748
rect 10788 2692 10844 2748
rect 10844 2692 10848 2748
rect 10784 2688 10848 2692
rect 10864 2748 10928 2752
rect 10864 2692 10868 2748
rect 10868 2692 10924 2748
rect 10924 2692 10928 2748
rect 10864 2688 10928 2692
rect 10944 2748 11008 2752
rect 10944 2692 10948 2748
rect 10948 2692 11004 2748
rect 11004 2692 11008 2748
rect 10944 2688 11008 2692
rect 11024 2748 11088 2752
rect 11024 2692 11028 2748
rect 11028 2692 11084 2748
rect 11084 2692 11088 2748
rect 11024 2688 11088 2692
rect 14717 2748 14781 2752
rect 14717 2692 14721 2748
rect 14721 2692 14777 2748
rect 14777 2692 14781 2748
rect 14717 2688 14781 2692
rect 14797 2748 14861 2752
rect 14797 2692 14801 2748
rect 14801 2692 14857 2748
rect 14857 2692 14861 2748
rect 14797 2688 14861 2692
rect 14877 2748 14941 2752
rect 14877 2692 14881 2748
rect 14881 2692 14937 2748
rect 14937 2692 14941 2748
rect 14877 2688 14941 2692
rect 14957 2748 15021 2752
rect 14957 2692 14961 2748
rect 14961 2692 15017 2748
rect 15017 2692 15021 2748
rect 14957 2688 15021 2692
rect 4884 2204 4948 2208
rect 4884 2148 4888 2204
rect 4888 2148 4944 2204
rect 4944 2148 4948 2204
rect 4884 2144 4948 2148
rect 4964 2204 5028 2208
rect 4964 2148 4968 2204
rect 4968 2148 5024 2204
rect 5024 2148 5028 2204
rect 4964 2144 5028 2148
rect 5044 2204 5108 2208
rect 5044 2148 5048 2204
rect 5048 2148 5104 2204
rect 5104 2148 5108 2204
rect 5044 2144 5108 2148
rect 5124 2204 5188 2208
rect 5124 2148 5128 2204
rect 5128 2148 5184 2204
rect 5184 2148 5188 2204
rect 5124 2144 5188 2148
rect 8817 2204 8881 2208
rect 8817 2148 8821 2204
rect 8821 2148 8877 2204
rect 8877 2148 8881 2204
rect 8817 2144 8881 2148
rect 8897 2204 8961 2208
rect 8897 2148 8901 2204
rect 8901 2148 8957 2204
rect 8957 2148 8961 2204
rect 8897 2144 8961 2148
rect 8977 2204 9041 2208
rect 8977 2148 8981 2204
rect 8981 2148 9037 2204
rect 9037 2148 9041 2204
rect 8977 2144 9041 2148
rect 9057 2204 9121 2208
rect 9057 2148 9061 2204
rect 9061 2148 9117 2204
rect 9117 2148 9121 2204
rect 9057 2144 9121 2148
rect 12750 2204 12814 2208
rect 12750 2148 12754 2204
rect 12754 2148 12810 2204
rect 12810 2148 12814 2204
rect 12750 2144 12814 2148
rect 12830 2204 12894 2208
rect 12830 2148 12834 2204
rect 12834 2148 12890 2204
rect 12890 2148 12894 2204
rect 12830 2144 12894 2148
rect 12910 2204 12974 2208
rect 12910 2148 12914 2204
rect 12914 2148 12970 2204
rect 12970 2148 12974 2204
rect 12910 2144 12974 2148
rect 12990 2204 13054 2208
rect 12990 2148 12994 2204
rect 12994 2148 13050 2204
rect 13050 2148 13054 2204
rect 12990 2144 13054 2148
rect 16683 2204 16747 2208
rect 16683 2148 16687 2204
rect 16687 2148 16743 2204
rect 16743 2148 16747 2204
rect 16683 2144 16747 2148
rect 16763 2204 16827 2208
rect 16763 2148 16767 2204
rect 16767 2148 16823 2204
rect 16823 2148 16827 2204
rect 16763 2144 16827 2148
rect 16843 2204 16907 2208
rect 16843 2148 16847 2204
rect 16847 2148 16903 2204
rect 16903 2148 16907 2204
rect 16843 2144 16907 2148
rect 16923 2204 16987 2208
rect 16923 2148 16927 2204
rect 16927 2148 16983 2204
rect 16983 2148 16987 2204
rect 16923 2144 16987 2148
<< metal4 >>
rect 2910 15808 3230 15824
rect 2910 15744 2918 15808
rect 2982 15744 2998 15808
rect 3062 15744 3078 15808
rect 3142 15744 3158 15808
rect 3222 15744 3230 15808
rect 2910 14720 3230 15744
rect 2910 14656 2918 14720
rect 2982 14656 2998 14720
rect 3062 14656 3078 14720
rect 3142 14656 3158 14720
rect 3222 14656 3230 14720
rect 2910 13632 3230 14656
rect 2910 13568 2918 13632
rect 2982 13568 2998 13632
rect 3062 13568 3078 13632
rect 3142 13568 3158 13632
rect 3222 13568 3230 13632
rect 2910 12544 3230 13568
rect 2910 12480 2918 12544
rect 2982 12480 2998 12544
rect 3062 12480 3078 12544
rect 3142 12480 3158 12544
rect 3222 12480 3230 12544
rect 2910 11456 3230 12480
rect 2910 11392 2918 11456
rect 2982 11392 2998 11456
rect 3062 11392 3078 11456
rect 3142 11392 3158 11456
rect 3222 11392 3230 11456
rect 2910 10368 3230 11392
rect 2910 10304 2918 10368
rect 2982 10304 2998 10368
rect 3062 10304 3078 10368
rect 3142 10304 3158 10368
rect 3222 10304 3230 10368
rect 2910 9280 3230 10304
rect 4876 15264 5196 15824
rect 4876 15200 4884 15264
rect 4948 15200 4964 15264
rect 5028 15200 5044 15264
rect 5108 15200 5124 15264
rect 5188 15200 5196 15264
rect 4876 14176 5196 15200
rect 4876 14112 4884 14176
rect 4948 14112 4964 14176
rect 5028 14112 5044 14176
rect 5108 14112 5124 14176
rect 5188 14112 5196 14176
rect 4876 13088 5196 14112
rect 4876 13024 4884 13088
rect 4948 13024 4964 13088
rect 5028 13024 5044 13088
rect 5108 13024 5124 13088
rect 5188 13024 5196 13088
rect 4876 12000 5196 13024
rect 4876 11936 4884 12000
rect 4948 11936 4964 12000
rect 5028 11936 5044 12000
rect 5108 11936 5124 12000
rect 5188 11936 5196 12000
rect 4876 10912 5196 11936
rect 4876 10848 4884 10912
rect 4948 10848 4964 10912
rect 5028 10848 5044 10912
rect 5108 10848 5124 10912
rect 5188 10848 5196 10912
rect 4876 9824 5196 10848
rect 4876 9760 4884 9824
rect 4948 9760 4964 9824
rect 5028 9760 5044 9824
rect 5108 9760 5124 9824
rect 5188 9760 5196 9824
rect 3371 9756 3437 9757
rect 3371 9692 3372 9756
rect 3436 9692 3437 9756
rect 3371 9691 3437 9692
rect 2910 9216 2918 9280
rect 2982 9216 2998 9280
rect 3062 9216 3078 9280
rect 3142 9216 3158 9280
rect 3222 9216 3230 9280
rect 2910 8192 3230 9216
rect 2910 8128 2918 8192
rect 2982 8128 2998 8192
rect 3062 8128 3078 8192
rect 3142 8128 3158 8192
rect 3222 8128 3230 8192
rect 2910 7104 3230 8128
rect 2910 7040 2918 7104
rect 2982 7040 2998 7104
rect 3062 7040 3078 7104
rect 3142 7040 3158 7104
rect 3222 7040 3230 7104
rect 2910 6016 3230 7040
rect 2910 5952 2918 6016
rect 2982 5952 2998 6016
rect 3062 5952 3078 6016
rect 3142 5952 3158 6016
rect 3222 5952 3230 6016
rect 2910 4928 3230 5952
rect 2910 4864 2918 4928
rect 2982 4864 2998 4928
rect 3062 4864 3078 4928
rect 3142 4864 3158 4928
rect 3222 4864 3230 4928
rect 2910 3840 3230 4864
rect 3374 4045 3434 9691
rect 4876 8736 5196 9760
rect 4876 8672 4884 8736
rect 4948 8672 4964 8736
rect 5028 8672 5044 8736
rect 5108 8672 5124 8736
rect 5188 8672 5196 8736
rect 4876 7648 5196 8672
rect 4876 7584 4884 7648
rect 4948 7584 4964 7648
rect 5028 7584 5044 7648
rect 5108 7584 5124 7648
rect 5188 7584 5196 7648
rect 4876 6560 5196 7584
rect 4876 6496 4884 6560
rect 4948 6496 4964 6560
rect 5028 6496 5044 6560
rect 5108 6496 5124 6560
rect 5188 6496 5196 6560
rect 4876 5472 5196 6496
rect 4876 5408 4884 5472
rect 4948 5408 4964 5472
rect 5028 5408 5044 5472
rect 5108 5408 5124 5472
rect 5188 5408 5196 5472
rect 4876 4384 5196 5408
rect 4876 4320 4884 4384
rect 4948 4320 4964 4384
rect 5028 4320 5044 4384
rect 5108 4320 5124 4384
rect 5188 4320 5196 4384
rect 3371 4044 3437 4045
rect 3371 3980 3372 4044
rect 3436 3980 3437 4044
rect 3371 3979 3437 3980
rect 2910 3776 2918 3840
rect 2982 3776 2998 3840
rect 3062 3776 3078 3840
rect 3142 3776 3158 3840
rect 3222 3776 3230 3840
rect 2910 2752 3230 3776
rect 2910 2688 2918 2752
rect 2982 2688 2998 2752
rect 3062 2688 3078 2752
rect 3142 2688 3158 2752
rect 3222 2688 3230 2752
rect 2910 2128 3230 2688
rect 4876 3296 5196 4320
rect 4876 3232 4884 3296
rect 4948 3232 4964 3296
rect 5028 3232 5044 3296
rect 5108 3232 5124 3296
rect 5188 3232 5196 3296
rect 4876 2208 5196 3232
rect 4876 2144 4884 2208
rect 4948 2144 4964 2208
rect 5028 2144 5044 2208
rect 5108 2144 5124 2208
rect 5188 2144 5196 2208
rect 4876 2128 5196 2144
rect 6843 15808 7163 15824
rect 6843 15744 6851 15808
rect 6915 15744 6931 15808
rect 6995 15744 7011 15808
rect 7075 15744 7091 15808
rect 7155 15744 7163 15808
rect 6843 14720 7163 15744
rect 6843 14656 6851 14720
rect 6915 14656 6931 14720
rect 6995 14656 7011 14720
rect 7075 14656 7091 14720
rect 7155 14656 7163 14720
rect 6843 13632 7163 14656
rect 6843 13568 6851 13632
rect 6915 13568 6931 13632
rect 6995 13568 7011 13632
rect 7075 13568 7091 13632
rect 7155 13568 7163 13632
rect 6843 12544 7163 13568
rect 6843 12480 6851 12544
rect 6915 12480 6931 12544
rect 6995 12480 7011 12544
rect 7075 12480 7091 12544
rect 7155 12480 7163 12544
rect 6843 11456 7163 12480
rect 6843 11392 6851 11456
rect 6915 11392 6931 11456
rect 6995 11392 7011 11456
rect 7075 11392 7091 11456
rect 7155 11392 7163 11456
rect 6843 10368 7163 11392
rect 6843 10304 6851 10368
rect 6915 10304 6931 10368
rect 6995 10304 7011 10368
rect 7075 10304 7091 10368
rect 7155 10304 7163 10368
rect 6843 9280 7163 10304
rect 6843 9216 6851 9280
rect 6915 9216 6931 9280
rect 6995 9216 7011 9280
rect 7075 9216 7091 9280
rect 7155 9216 7163 9280
rect 6843 8192 7163 9216
rect 6843 8128 6851 8192
rect 6915 8128 6931 8192
rect 6995 8128 7011 8192
rect 7075 8128 7091 8192
rect 7155 8128 7163 8192
rect 6843 7104 7163 8128
rect 6843 7040 6851 7104
rect 6915 7040 6931 7104
rect 6995 7040 7011 7104
rect 7075 7040 7091 7104
rect 7155 7040 7163 7104
rect 6843 6016 7163 7040
rect 6843 5952 6851 6016
rect 6915 5952 6931 6016
rect 6995 5952 7011 6016
rect 7075 5952 7091 6016
rect 7155 5952 7163 6016
rect 6843 4928 7163 5952
rect 6843 4864 6851 4928
rect 6915 4864 6931 4928
rect 6995 4864 7011 4928
rect 7075 4864 7091 4928
rect 7155 4864 7163 4928
rect 6843 3840 7163 4864
rect 6843 3776 6851 3840
rect 6915 3776 6931 3840
rect 6995 3776 7011 3840
rect 7075 3776 7091 3840
rect 7155 3776 7163 3840
rect 6843 2752 7163 3776
rect 6843 2688 6851 2752
rect 6915 2688 6931 2752
rect 6995 2688 7011 2752
rect 7075 2688 7091 2752
rect 7155 2688 7163 2752
rect 6843 2128 7163 2688
rect 8809 15264 9129 15824
rect 8809 15200 8817 15264
rect 8881 15200 8897 15264
rect 8961 15200 8977 15264
rect 9041 15200 9057 15264
rect 9121 15200 9129 15264
rect 8809 14176 9129 15200
rect 8809 14112 8817 14176
rect 8881 14112 8897 14176
rect 8961 14112 8977 14176
rect 9041 14112 9057 14176
rect 9121 14112 9129 14176
rect 8809 13088 9129 14112
rect 8809 13024 8817 13088
rect 8881 13024 8897 13088
rect 8961 13024 8977 13088
rect 9041 13024 9057 13088
rect 9121 13024 9129 13088
rect 8809 12000 9129 13024
rect 8809 11936 8817 12000
rect 8881 11936 8897 12000
rect 8961 11936 8977 12000
rect 9041 11936 9057 12000
rect 9121 11936 9129 12000
rect 8809 10912 9129 11936
rect 8809 10848 8817 10912
rect 8881 10848 8897 10912
rect 8961 10848 8977 10912
rect 9041 10848 9057 10912
rect 9121 10848 9129 10912
rect 8809 9824 9129 10848
rect 8809 9760 8817 9824
rect 8881 9760 8897 9824
rect 8961 9760 8977 9824
rect 9041 9760 9057 9824
rect 9121 9760 9129 9824
rect 8809 8736 9129 9760
rect 8809 8672 8817 8736
rect 8881 8672 8897 8736
rect 8961 8672 8977 8736
rect 9041 8672 9057 8736
rect 9121 8672 9129 8736
rect 8809 7648 9129 8672
rect 8809 7584 8817 7648
rect 8881 7584 8897 7648
rect 8961 7584 8977 7648
rect 9041 7584 9057 7648
rect 9121 7584 9129 7648
rect 8809 6560 9129 7584
rect 8809 6496 8817 6560
rect 8881 6496 8897 6560
rect 8961 6496 8977 6560
rect 9041 6496 9057 6560
rect 9121 6496 9129 6560
rect 8809 5472 9129 6496
rect 8809 5408 8817 5472
rect 8881 5408 8897 5472
rect 8961 5408 8977 5472
rect 9041 5408 9057 5472
rect 9121 5408 9129 5472
rect 8809 4384 9129 5408
rect 8809 4320 8817 4384
rect 8881 4320 8897 4384
rect 8961 4320 8977 4384
rect 9041 4320 9057 4384
rect 9121 4320 9129 4384
rect 8809 3296 9129 4320
rect 8809 3232 8817 3296
rect 8881 3232 8897 3296
rect 8961 3232 8977 3296
rect 9041 3232 9057 3296
rect 9121 3232 9129 3296
rect 8809 2208 9129 3232
rect 8809 2144 8817 2208
rect 8881 2144 8897 2208
rect 8961 2144 8977 2208
rect 9041 2144 9057 2208
rect 9121 2144 9129 2208
rect 8809 2128 9129 2144
rect 10776 15808 11096 15824
rect 10776 15744 10784 15808
rect 10848 15744 10864 15808
rect 10928 15744 10944 15808
rect 11008 15744 11024 15808
rect 11088 15744 11096 15808
rect 10776 14720 11096 15744
rect 10776 14656 10784 14720
rect 10848 14656 10864 14720
rect 10928 14656 10944 14720
rect 11008 14656 11024 14720
rect 11088 14656 11096 14720
rect 10776 13632 11096 14656
rect 10776 13568 10784 13632
rect 10848 13568 10864 13632
rect 10928 13568 10944 13632
rect 11008 13568 11024 13632
rect 11088 13568 11096 13632
rect 10776 12544 11096 13568
rect 10776 12480 10784 12544
rect 10848 12480 10864 12544
rect 10928 12480 10944 12544
rect 11008 12480 11024 12544
rect 11088 12480 11096 12544
rect 10776 11456 11096 12480
rect 10776 11392 10784 11456
rect 10848 11392 10864 11456
rect 10928 11392 10944 11456
rect 11008 11392 11024 11456
rect 11088 11392 11096 11456
rect 10776 10368 11096 11392
rect 10776 10304 10784 10368
rect 10848 10304 10864 10368
rect 10928 10304 10944 10368
rect 11008 10304 11024 10368
rect 11088 10304 11096 10368
rect 10776 9280 11096 10304
rect 10776 9216 10784 9280
rect 10848 9216 10864 9280
rect 10928 9216 10944 9280
rect 11008 9216 11024 9280
rect 11088 9216 11096 9280
rect 10776 8192 11096 9216
rect 10776 8128 10784 8192
rect 10848 8128 10864 8192
rect 10928 8128 10944 8192
rect 11008 8128 11024 8192
rect 11088 8128 11096 8192
rect 10776 7104 11096 8128
rect 10776 7040 10784 7104
rect 10848 7040 10864 7104
rect 10928 7040 10944 7104
rect 11008 7040 11024 7104
rect 11088 7040 11096 7104
rect 10776 6016 11096 7040
rect 10776 5952 10784 6016
rect 10848 5952 10864 6016
rect 10928 5952 10944 6016
rect 11008 5952 11024 6016
rect 11088 5952 11096 6016
rect 10776 4928 11096 5952
rect 10776 4864 10784 4928
rect 10848 4864 10864 4928
rect 10928 4864 10944 4928
rect 11008 4864 11024 4928
rect 11088 4864 11096 4928
rect 10776 3840 11096 4864
rect 10776 3776 10784 3840
rect 10848 3776 10864 3840
rect 10928 3776 10944 3840
rect 11008 3776 11024 3840
rect 11088 3776 11096 3840
rect 10776 2752 11096 3776
rect 10776 2688 10784 2752
rect 10848 2688 10864 2752
rect 10928 2688 10944 2752
rect 11008 2688 11024 2752
rect 11088 2688 11096 2752
rect 10776 2128 11096 2688
rect 12742 15264 13062 15824
rect 12742 15200 12750 15264
rect 12814 15200 12830 15264
rect 12894 15200 12910 15264
rect 12974 15200 12990 15264
rect 13054 15200 13062 15264
rect 12742 14176 13062 15200
rect 12742 14112 12750 14176
rect 12814 14112 12830 14176
rect 12894 14112 12910 14176
rect 12974 14112 12990 14176
rect 13054 14112 13062 14176
rect 12742 13088 13062 14112
rect 12742 13024 12750 13088
rect 12814 13024 12830 13088
rect 12894 13024 12910 13088
rect 12974 13024 12990 13088
rect 13054 13024 13062 13088
rect 12742 12000 13062 13024
rect 12742 11936 12750 12000
rect 12814 11936 12830 12000
rect 12894 11936 12910 12000
rect 12974 11936 12990 12000
rect 13054 11936 13062 12000
rect 12742 10912 13062 11936
rect 12742 10848 12750 10912
rect 12814 10848 12830 10912
rect 12894 10848 12910 10912
rect 12974 10848 12990 10912
rect 13054 10848 13062 10912
rect 12742 9824 13062 10848
rect 12742 9760 12750 9824
rect 12814 9760 12830 9824
rect 12894 9760 12910 9824
rect 12974 9760 12990 9824
rect 13054 9760 13062 9824
rect 12742 8736 13062 9760
rect 12742 8672 12750 8736
rect 12814 8672 12830 8736
rect 12894 8672 12910 8736
rect 12974 8672 12990 8736
rect 13054 8672 13062 8736
rect 12742 7648 13062 8672
rect 12742 7584 12750 7648
rect 12814 7584 12830 7648
rect 12894 7584 12910 7648
rect 12974 7584 12990 7648
rect 13054 7584 13062 7648
rect 12742 6560 13062 7584
rect 12742 6496 12750 6560
rect 12814 6496 12830 6560
rect 12894 6496 12910 6560
rect 12974 6496 12990 6560
rect 13054 6496 13062 6560
rect 12742 5472 13062 6496
rect 12742 5408 12750 5472
rect 12814 5408 12830 5472
rect 12894 5408 12910 5472
rect 12974 5408 12990 5472
rect 13054 5408 13062 5472
rect 12742 4384 13062 5408
rect 12742 4320 12750 4384
rect 12814 4320 12830 4384
rect 12894 4320 12910 4384
rect 12974 4320 12990 4384
rect 13054 4320 13062 4384
rect 12742 3296 13062 4320
rect 12742 3232 12750 3296
rect 12814 3232 12830 3296
rect 12894 3232 12910 3296
rect 12974 3232 12990 3296
rect 13054 3232 13062 3296
rect 12742 2208 13062 3232
rect 12742 2144 12750 2208
rect 12814 2144 12830 2208
rect 12894 2144 12910 2208
rect 12974 2144 12990 2208
rect 13054 2144 13062 2208
rect 12742 2128 13062 2144
rect 14709 15808 15029 15824
rect 14709 15744 14717 15808
rect 14781 15744 14797 15808
rect 14861 15744 14877 15808
rect 14941 15744 14957 15808
rect 15021 15744 15029 15808
rect 14709 14720 15029 15744
rect 14709 14656 14717 14720
rect 14781 14656 14797 14720
rect 14861 14656 14877 14720
rect 14941 14656 14957 14720
rect 15021 14656 15029 14720
rect 14709 13632 15029 14656
rect 14709 13568 14717 13632
rect 14781 13568 14797 13632
rect 14861 13568 14877 13632
rect 14941 13568 14957 13632
rect 15021 13568 15029 13632
rect 14709 12544 15029 13568
rect 14709 12480 14717 12544
rect 14781 12480 14797 12544
rect 14861 12480 14877 12544
rect 14941 12480 14957 12544
rect 15021 12480 15029 12544
rect 14709 11456 15029 12480
rect 14709 11392 14717 11456
rect 14781 11392 14797 11456
rect 14861 11392 14877 11456
rect 14941 11392 14957 11456
rect 15021 11392 15029 11456
rect 14709 10368 15029 11392
rect 14709 10304 14717 10368
rect 14781 10304 14797 10368
rect 14861 10304 14877 10368
rect 14941 10304 14957 10368
rect 15021 10304 15029 10368
rect 14709 9280 15029 10304
rect 14709 9216 14717 9280
rect 14781 9216 14797 9280
rect 14861 9216 14877 9280
rect 14941 9216 14957 9280
rect 15021 9216 15029 9280
rect 14709 8192 15029 9216
rect 14709 8128 14717 8192
rect 14781 8128 14797 8192
rect 14861 8128 14877 8192
rect 14941 8128 14957 8192
rect 15021 8128 15029 8192
rect 14709 7104 15029 8128
rect 14709 7040 14717 7104
rect 14781 7040 14797 7104
rect 14861 7040 14877 7104
rect 14941 7040 14957 7104
rect 15021 7040 15029 7104
rect 14709 6016 15029 7040
rect 14709 5952 14717 6016
rect 14781 5952 14797 6016
rect 14861 5952 14877 6016
rect 14941 5952 14957 6016
rect 15021 5952 15029 6016
rect 14709 4928 15029 5952
rect 14709 4864 14717 4928
rect 14781 4864 14797 4928
rect 14861 4864 14877 4928
rect 14941 4864 14957 4928
rect 15021 4864 15029 4928
rect 14709 3840 15029 4864
rect 14709 3776 14717 3840
rect 14781 3776 14797 3840
rect 14861 3776 14877 3840
rect 14941 3776 14957 3840
rect 15021 3776 15029 3840
rect 14709 2752 15029 3776
rect 14709 2688 14717 2752
rect 14781 2688 14797 2752
rect 14861 2688 14877 2752
rect 14941 2688 14957 2752
rect 15021 2688 15029 2752
rect 14709 2128 15029 2688
rect 16675 15264 16995 15824
rect 16675 15200 16683 15264
rect 16747 15200 16763 15264
rect 16827 15200 16843 15264
rect 16907 15200 16923 15264
rect 16987 15200 16995 15264
rect 16675 14176 16995 15200
rect 16675 14112 16683 14176
rect 16747 14112 16763 14176
rect 16827 14112 16843 14176
rect 16907 14112 16923 14176
rect 16987 14112 16995 14176
rect 16675 13088 16995 14112
rect 16675 13024 16683 13088
rect 16747 13024 16763 13088
rect 16827 13024 16843 13088
rect 16907 13024 16923 13088
rect 16987 13024 16995 13088
rect 16675 12000 16995 13024
rect 16675 11936 16683 12000
rect 16747 11936 16763 12000
rect 16827 11936 16843 12000
rect 16907 11936 16923 12000
rect 16987 11936 16995 12000
rect 16675 10912 16995 11936
rect 16675 10848 16683 10912
rect 16747 10848 16763 10912
rect 16827 10848 16843 10912
rect 16907 10848 16923 10912
rect 16987 10848 16995 10912
rect 16675 9824 16995 10848
rect 16675 9760 16683 9824
rect 16747 9760 16763 9824
rect 16827 9760 16843 9824
rect 16907 9760 16923 9824
rect 16987 9760 16995 9824
rect 16675 8736 16995 9760
rect 16675 8672 16683 8736
rect 16747 8672 16763 8736
rect 16827 8672 16843 8736
rect 16907 8672 16923 8736
rect 16987 8672 16995 8736
rect 16675 7648 16995 8672
rect 16675 7584 16683 7648
rect 16747 7584 16763 7648
rect 16827 7584 16843 7648
rect 16907 7584 16923 7648
rect 16987 7584 16995 7648
rect 16675 6560 16995 7584
rect 16675 6496 16683 6560
rect 16747 6496 16763 6560
rect 16827 6496 16843 6560
rect 16907 6496 16923 6560
rect 16987 6496 16995 6560
rect 16675 5472 16995 6496
rect 16675 5408 16683 5472
rect 16747 5408 16763 5472
rect 16827 5408 16843 5472
rect 16907 5408 16923 5472
rect 16987 5408 16995 5472
rect 16675 4384 16995 5408
rect 16675 4320 16683 4384
rect 16747 4320 16763 4384
rect 16827 4320 16843 4384
rect 16907 4320 16923 4384
rect 16987 4320 16995 4384
rect 16675 3296 16995 4320
rect 16675 3232 16683 3296
rect 16747 3232 16763 3296
rect 16827 3232 16843 3296
rect 16907 3232 16923 3296
rect 16987 3232 16995 3296
rect 16675 2208 16995 3232
rect 16675 2144 16683 2208
rect 16747 2144 16763 2208
rect 16827 2144 16843 2208
rect 16907 2144 16923 2208
rect 16987 2144 16995 2208
rect 16675 2128 16995 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__216__1_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 15732 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__2_A
timestamp 1666464484
transform -1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__3_A
timestamp 1666464484
transform 1 0 14904 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__4_A
timestamp 1666464484
transform 1 0 14904 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__6_A
timestamp 1666464484
transform 1 0 4048 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__8_A
timestamp 1666464484
transform -1 0 4784 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1666464484
transform -1 0 6716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 15732 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1666464484
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1666464484
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_9
timestamp 1666464484
transform 1 0 1932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_21
timestamp 1666464484
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_34
timestamp 1666464484
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1666464484
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1666464484
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1666464484
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_11
timestamp 1666464484
transform 1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_15
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_19
timestamp 1666464484
transform 1 0 2852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1666464484
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_34
timestamp 1666464484
transform 1 0 4232 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_40
timestamp 1666464484
transform 1 0 4784 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_52
timestamp 1666464484
transform 1 0 5888 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_64
timestamp 1666464484
transform 1 0 6992 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_76
timestamp 1666464484
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1666464484
transform 1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_13
timestamp 1666464484
transform 1 0 2300 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_21
timestamp 1666464484
transform 1 0 3036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_28
timestamp 1666464484
transform 1 0 3680 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_34
timestamp 1666464484
transform 1 0 4232 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_41
timestamp 1666464484
transform 1 0 4876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1666464484
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_90
timestamp 1666464484
transform 1 0 9384 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_102
timestamp 1666464484
transform 1 0 10488 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1666464484
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_9
timestamp 1666464484
transform 1 0 1932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_13
timestamp 1666464484
transform 1 0 2300 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_18
timestamp 1666464484
transform 1 0 2760 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1666464484
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_34
timestamp 1666464484
transform 1 0 4232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_45
timestamp 1666464484
transform 1 0 5244 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_50
timestamp 1666464484
transform 1 0 5704 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_62
timestamp 1666464484
transform 1 0 6808 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_68
timestamp 1666464484
transform 1 0 7360 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_73
timestamp 1666464484
transform 1 0 7820 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1666464484
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1666464484
transform 1 0 9660 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_11
timestamp 1666464484
transform 1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_20
timestamp 1666464484
transform 1 0 2944 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_36
timestamp 1666464484
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_43
timestamp 1666464484
transform 1 0 5060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_47
timestamp 1666464484
transform 1 0 5428 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1666464484
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_64
timestamp 1666464484
transform 1 0 6992 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_72
timestamp 1666464484
transform 1 0 7728 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_100
timestamp 1666464484
transform 1 0 10304 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_13
timestamp 1666464484
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1666464484
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_35
timestamp 1666464484
transform 1 0 4324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_73
timestamp 1666464484
transform 1 0 7820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1666464484
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_111
timestamp 1666464484
transform 1 0 11316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_123
timestamp 1666464484
transform 1 0 12420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1666464484
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_9
timestamp 1666464484
transform 1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_19
timestamp 1666464484
transform 1 0 2852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_23
timestamp 1666464484
transform 1 0 3220 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1666464484
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_77
timestamp 1666464484
transform 1 0 8188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_88
timestamp 1666464484
transform 1 0 9200 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_96
timestamp 1666464484
transform 1 0 9936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_100
timestamp 1666464484
transform 1 0 10304 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1666464484
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_120
timestamp 1666464484
transform 1 0 12144 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_132
timestamp 1666464484
transform 1 0 13248 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_144
timestamp 1666464484
transform 1 0 14352 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_156
timestamp 1666464484
transform 1 0 15456 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_11
timestamp 1666464484
transform 1 0 2116 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1666464484
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_36
timestamp 1666464484
transform 1 0 4416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_60
timestamp 1666464484
transform 1 0 6624 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1666464484
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_90
timestamp 1666464484
transform 1 0 9384 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_118
timestamp 1666464484
transform 1 0 11960 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_129
timestamp 1666464484
transform 1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1666464484
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_11
timestamp 1666464484
transform 1 0 2116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_19
timestamp 1666464484
transform 1 0 2852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1666464484
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_33
timestamp 1666464484
transform 1 0 4140 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1666464484
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_63
timestamp 1666464484
transform 1 0 6900 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1666464484
transform 1 0 7636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_104
timestamp 1666464484
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_119
timestamp 1666464484
transform 1 0 12052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_126
timestamp 1666464484
transform 1 0 12696 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_133
timestamp 1666464484
transform 1 0 13340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_145
timestamp 1666464484
transform 1 0 14444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_157
timestamp 1666464484
transform 1 0 15548 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1666464484
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_9
timestamp 1666464484
transform 1 0 1932 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_13
timestamp 1666464484
transform 1 0 2300 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_18
timestamp 1666464484
transform 1 0 2760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1666464484
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_36
timestamp 1666464484
transform 1 0 4416 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_44
timestamp 1666464484
transform 1 0 5152 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_73
timestamp 1666464484
transform 1 0 7820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1666464484
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_90
timestamp 1666464484
transform 1 0 9384 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_98
timestamp 1666464484
transform 1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_120
timestamp 1666464484
transform 1 0 12144 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_128
timestamp 1666464484
transform 1 0 12880 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 1666464484
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_9
timestamp 1666464484
transform 1 0 1932 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_17
timestamp 1666464484
transform 1 0 2668 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_38
timestamp 1666464484
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_45
timestamp 1666464484
transform 1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1666464484
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_68
timestamp 1666464484
transform 1 0 7360 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_74
timestamp 1666464484
transform 1 0 7912 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_95
timestamp 1666464484
transform 1 0 9844 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_103
timestamp 1666464484
transform 1 0 10580 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1666464484
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_120
timestamp 1666464484
transform 1 0 12144 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_148
timestamp 1666464484
transform 1 0 14720 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_154
timestamp 1666464484
transform 1 0 15272 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_158
timestamp 1666464484
transform 1 0 15640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1666464484
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1666464484
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_37
timestamp 1666464484
transform 1 0 4508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_61
timestamp 1666464484
transform 1 0 6716 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1666464484
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1666464484
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_117
timestamp 1666464484
transform 1 0 11868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_125
timestamp 1666464484
transform 1 0 12604 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_147
timestamp 1666464484
transform 1 0 14628 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_155
timestamp 1666464484
transform 1 0 15364 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_162
timestamp 1666464484
transform 1 0 16008 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1666464484
transform 1 0 1932 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_14
timestamp 1666464484
transform 1 0 2392 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_42
timestamp 1666464484
transform 1 0 4968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_48
timestamp 1666464484
transform 1 0 5520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1666464484
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_64
timestamp 1666464484
transform 1 0 6992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_72
timestamp 1666464484
transform 1 0 7728 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_96
timestamp 1666464484
transform 1 0 9936 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1666464484
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_138
timestamp 1666464484
transform 1 0 13800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_162
timestamp 1666464484
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_22
timestamp 1666464484
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_38
timestamp 1666464484
transform 1 0 4600 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_44
timestamp 1666464484
transform 1 0 5152 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_78
timestamp 1666464484
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_92
timestamp 1666464484
transform 1 0 9568 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_100
timestamp 1666464484
transform 1 0 10304 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_129
timestamp 1666464484
transform 1 0 12972 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1666464484
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_163
timestamp 1666464484
transform 1 0 16100 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_167
timestamp 1666464484
transform 1 0 16468 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1666464484
transform 1 0 1932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_30
timestamp 1666464484
transform 1 0 3864 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1666464484
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_79
timestamp 1666464484
transform 1 0 8372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_101
timestamp 1666464484
transform 1 0 10396 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1666464484
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_135
timestamp 1666464484
transform 1 0 13524 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_159
timestamp 1666464484
transform 1 0 15732 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1666464484
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_9
timestamp 1666464484
transform 1 0 1932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_13
timestamp 1666464484
transform 1 0 2300 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_18
timestamp 1666464484
transform 1 0 2760 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1666464484
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_33
timestamp 1666464484
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_39
timestamp 1666464484
transform 1 0 4692 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_45
timestamp 1666464484
transform 1 0 5244 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_66
timestamp 1666464484
transform 1 0 7176 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_72
timestamp 1666464484
transform 1 0 7728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1666464484
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1666464484
transform 1 0 9660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_100
timestamp 1666464484
transform 1 0 10304 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_127
timestamp 1666464484
transform 1 0 12788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_131
timestamp 1666464484
transform 1 0 13156 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1666464484
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_146
timestamp 1666464484
transform 1 0 14536 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_160
timestamp 1666464484
transform 1 0 15824 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_10
timestamp 1666464484
transform 1 0 2024 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_16
timestamp 1666464484
transform 1 0 2576 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_21
timestamp 1666464484
transform 1 0 3036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_45
timestamp 1666464484
transform 1 0 5244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_49
timestamp 1666464484
transform 1 0 5612 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1666464484
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1666464484
transform 1 0 6808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_71
timestamp 1666464484
transform 1 0 7636 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_79
timestamp 1666464484
transform 1 0 8372 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_87
timestamp 1666464484
transform 1 0 9108 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1666464484
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_119
timestamp 1666464484
transform 1 0 12052 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_140
timestamp 1666464484
transform 1 0 13984 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1666464484
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_22
timestamp 1666464484
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_52
timestamp 1666464484
transform 1 0 5888 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_76
timestamp 1666464484
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_107
timestamp 1666464484
transform 1 0 10948 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_115
timestamp 1666464484
transform 1 0 11684 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_123
timestamp 1666464484
transform 1 0 12420 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_127
timestamp 1666464484
transform 1 0 12788 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_132
timestamp 1666464484
transform 1 0 13248 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_146
timestamp 1666464484
transform 1 0 14536 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_159
timestamp 1666464484
transform 1 0 15732 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_167
timestamp 1666464484
transform 1 0 16468 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_25
timestamp 1666464484
transform 1 0 3404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_29
timestamp 1666464484
transform 1 0 3772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_33
timestamp 1666464484
transform 1 0 4140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1666464484
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_64
timestamp 1666464484
transform 1 0 6992 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_72
timestamp 1666464484
transform 1 0 7728 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_76
timestamp 1666464484
transform 1 0 8096 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_85
timestamp 1666464484
transform 1 0 8924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1666464484
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_117
timestamp 1666464484
transform 1 0 11868 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_122
timestamp 1666464484
transform 1 0 12328 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_148
timestamp 1666464484
transform 1 0 14720 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_155
timestamp 1666464484
transform 1 0 15364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666464484
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_9
timestamp 1666464484
transform 1 0 1932 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_13
timestamp 1666464484
transform 1 0 2300 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1666464484
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1666464484
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_34
timestamp 1666464484
transform 1 0 4232 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_58
timestamp 1666464484
transform 1 0 6440 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1666464484
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_91
timestamp 1666464484
transform 1 0 9476 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_99
timestamp 1666464484
transform 1 0 10212 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_105
timestamp 1666464484
transform 1 0 10764 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_129
timestamp 1666464484
transform 1 0 12972 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1666464484
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_146
timestamp 1666464484
transform 1 0 14536 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666464484
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_165
timestamp 1666464484
transform 1 0 16284 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_9
timestamp 1666464484
transform 1 0 1932 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_13
timestamp 1666464484
transform 1 0 2300 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_30
timestamp 1666464484
transform 1 0 3864 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1666464484
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_61
timestamp 1666464484
transform 1 0 6716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_100
timestamp 1666464484
transform 1 0 10304 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1666464484
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_119
timestamp 1666464484
transform 1 0 12052 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_130
timestamp 1666464484
transform 1 0 13064 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_138
timestamp 1666464484
transform 1 0 13800 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_145
timestamp 1666464484
transform 1 0 14444 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_157
timestamp 1666464484
transform 1 0 15548 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1666464484
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1666464484
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666464484
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_40
timestamp 1666464484
transform 1 0 4784 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_44
timestamp 1666464484
transform 1 0 5152 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_65
timestamp 1666464484
transform 1 0 7084 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_73
timestamp 1666464484
transform 1 0 7820 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1666464484
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_95
timestamp 1666464484
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_119
timestamp 1666464484
transform 1 0 12052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_126
timestamp 1666464484
transform 1 0 12696 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_146
timestamp 1666464484
transform 1 0 14536 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_152
timestamp 1666464484
transform 1 0 15088 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_164
timestamp 1666464484
transform 1 0 16192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_9
timestamp 1666464484
transform 1 0 1932 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_19
timestamp 1666464484
transform 1 0 2852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_43
timestamp 1666464484
transform 1 0 5060 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1666464484
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_79
timestamp 1666464484
transform 1 0 8372 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_103
timestamp 1666464484
transform 1 0 10580 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1666464484
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_118
timestamp 1666464484
transform 1 0 11960 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_132
timestamp 1666464484
transform 1 0 13248 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_139
timestamp 1666464484
transform 1 0 13892 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_146
timestamp 1666464484
transform 1 0 14536 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_152
timestamp 1666464484
transform 1 0 15088 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1666464484
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_13
timestamp 1666464484
transform 1 0 2300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1666464484
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_37
timestamp 1666464484
transform 1 0 4508 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_45
timestamp 1666464484
transform 1 0 5244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_49
timestamp 1666464484
transform 1 0 5612 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_54
timestamp 1666464484
transform 1 0 6072 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_57
timestamp 1666464484
transform 1 0 6348 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1666464484
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666464484
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_91
timestamp 1666464484
transform 1 0 9476 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1666464484
transform 1 0 10488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_113
timestamp 1666464484
transform 1 0 11500 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_118
timestamp 1666464484
transform 1 0 11960 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_125
timestamp 1666464484
transform 1 0 12604 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_132
timestamp 1666464484
transform 1 0 13248 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1666464484
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_153
timestamp 1666464484
transform 1 0 15180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_159
timestamp 1666464484
transform 1 0 15732 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_167
timestamp 1666464484
transform 1 0 16468 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 16836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 16836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 16836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1666464484
transform 1 0 6256 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1666464484
transform 1 0 11408 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 13248 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _108_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9660 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _109_
timestamp 1666464484
transform 1 0 6532 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _110__10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11224 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _111__11
timestamp 1666464484
transform -1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _112__12
timestamp 1666464484
transform 1 0 14904 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _113__13
timestamp 1666464484
transform 1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _114_
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _115_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7176 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _116_
timestamp 1666464484
transform -1 0 9568 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _117_
timestamp 1666464484
transform 1 0 9108 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _118_
timestamp 1666464484
transform 1 0 10672 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _119_
timestamp 1666464484
transform 1 0 5612 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _120_
timestamp 1666464484
transform 1 0 4048 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _121_
timestamp 1666464484
transform 1 0 4232 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _122_
timestamp 1666464484
transform 1 0 11684 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _123_
timestamp 1666464484
transform 1 0 10396 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _124_
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _125_
timestamp 1666464484
transform 1 0 11684 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _126_
timestamp 1666464484
transform 1 0 5612 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _127_
timestamp 1666464484
transform 1 0 6532 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _128__14
timestamp 1666464484
transform -1 0 15640 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _129__15
timestamp 1666464484
transform -1 0 14536 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _130__16
timestamp 1666464484
transform -1 0 15824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _131__17
timestamp 1666464484
transform -1 0 14536 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _132__18
timestamp 1666464484
transform -1 0 16008 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _133__19
timestamp 1666464484
transform -1 0 12696 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _134__20
timestamp 1666464484
transform -1 0 11960 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _135__21
timestamp 1666464484
transform -1 0 11132 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136__22
timestamp 1666464484
transform -1 0 12604 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _137_
timestamp 1666464484
transform 1 0 3956 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _138_
timestamp 1666464484
transform -1 0 6992 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _139_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2024 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1748 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _141_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11684 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _142_
timestamp 1666464484
transform 1 0 3956 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _143_
timestamp 1666464484
transform 1 0 3956 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1666464484
transform 1 0 14904 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _145_
timestamp 1666464484
transform -1 0 3220 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _146_
timestamp 1666464484
transform 1 0 2852 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _147_
timestamp 1666464484
transform 1 0 15088 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _148_
timestamp 1666464484
transform 1 0 1656 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _149_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1564 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1666464484
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _151_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12420 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _152_
timestamp 1666464484
transform 1 0 12972 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _153_
timestamp 1666464484
transform 1 0 11684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _154_
timestamp 1666464484
transform 1 0 7452 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _155_
timestamp 1666464484
transform 1 0 5336 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _156_
timestamp 1666464484
transform -1 0 3496 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _157_
timestamp 1666464484
transform -1 0 11132 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _158_
timestamp 1666464484
transform -1 0 7728 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _159_
timestamp 1666464484
transform -1 0 3036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _160_
timestamp 1666464484
transform 1 0 3128 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1666464484
transform -1 0 5060 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1666464484
transform -1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4600 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1666464484
transform 1 0 1840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1666464484
transform -1 0 4140 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1666464484
transform -1 0 5244 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _167_
timestamp 1666464484
transform 1 0 7820 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1666464484
transform 1 0 14260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1666464484
transform -1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 1666464484
transform 1 0 3956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1666464484
transform 1 0 10028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1666464484
transform -1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _174_
timestamp 1666464484
transform 1 0 10028 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1666464484
transform 1 0 12420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8188 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  _177_
timestamp 1666464484
transform 1 0 6992 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _178_
timestamp 1666464484
transform -1 0 4416 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _179_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9200 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _180_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 7360 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_4  _183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4508 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _184_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _185_
timestamp 1666464484
transform 1 0 13064 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _186_
timestamp 1666464484
transform -1 0 8280 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8648 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _188_
timestamp 1666464484
transform -1 0 2944 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3036 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1666464484
transform -1 0 3496 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2668 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _192_
timestamp 1666464484
transform -1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _194_
timestamp 1666464484
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _195_
timestamp 1666464484
transform -1 0 2760 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _196_
timestamp 1666464484
transform 1 0 4600 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _197_
timestamp 1666464484
transform 1 0 2300 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1656 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _199_
timestamp 1666464484
transform -1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _200_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2576 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _202_
timestamp 1666464484
transform 1 0 1564 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _203_
timestamp 1666464484
transform 1 0 1564 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _204_
timestamp 1666464484
transform -1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _205_
timestamp 1666464484
transform -1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _206_
timestamp 1666464484
transform -1 0 12052 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _207_
timestamp 1666464484
transform -1 0 12328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _208_
timestamp 1666464484
transform 1 0 13064 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _209_
timestamp 1666464484
transform 1 0 13248 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _210_
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _211_
timestamp 1666464484
transform -1 0 13800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _212_
timestamp 1666464484
transform -1 0 15364 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _213_
timestamp 1666464484
transform 1 0 12972 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _214_
timestamp 1666464484
transform -1 0 8556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1666464484
transform 1 0 12328 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216__1
timestamp 1666464484
transform -1 0 15180 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217__2
timestamp 1666464484
transform -1 0 13892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218__3
timestamp 1666464484
transform -1 0 14536 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219__4
timestamp 1666464484
transform -1 0 14536 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220__5
timestamp 1666464484
transform 1 0 14168 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _221__23
timestamp 1666464484
transform 1 0 13064 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _222_
timestamp 1666464484
transform 1 0 5704 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _223_
timestamp 1666464484
transform 1 0 9108 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _224_
timestamp 1666464484
transform -1 0 10488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _225_
timestamp 1666464484
transform -1 0 10764 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _226_
timestamp 1666464484
transform -1 0 14628 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _227_
timestamp 1666464484
transform -1 0 13708 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _228_
timestamp 1666464484
transform -1 0 13248 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _229_
timestamp 1666464484
transform 1 0 12696 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _230_
timestamp 1666464484
transform -1 0 12972 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _231__6
timestamp 1666464484
transform -1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232__7
timestamp 1666464484
transform -1 0 10304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _233_
timestamp 1666464484
transform -1 0 4876 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _234_
timestamp 1666464484
transform -1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _235_
timestamp 1666464484
transform -1 0 2760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1666464484
transform -1 0 12972 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _237_
timestamp 1666464484
transform -1 0 7820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _238_
timestamp 1666464484
transform -1 0 9936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _239_
timestamp 1666464484
transform -1 0 11132 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _240__8
timestamp 1666464484
transform -1 0 3680 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241__9
timestamp 1666464484
transform -1 0 9384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _242_
timestamp 1666464484
transform -1 0 2760 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _243_
timestamp 1666464484
transform -1 0 2392 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _244_
timestamp 1666464484
transform 1 0 7360 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _245_
timestamp 1666464484
transform -1 0 4416 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _246_
timestamp 1666464484
transform 1 0 9292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _247_
timestamp 1666464484
transform 1 0 8004 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _248_
timestamp 1666464484
transform 1 0 5704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _249_
timestamp 1666464484
transform -1 0 6992 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _250_
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _251_
timestamp 1666464484
transform 1 0 11316 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _252_
timestamp 1666464484
transform 1 0 9108 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _253_
timestamp 1666464484
transform -1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _254__24
timestamp 1666464484
transform -1 0 6072 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3128 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _256_
timestamp 1666464484
transform -1 0 3864 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _257_
timestamp 1666464484
transform -1 0 5060 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _258_
timestamp 1666464484
transform -1 0 3036 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _259_
timestamp 1666464484
transform 1 0 4508 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6072 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _261_
timestamp 1666464484
transform 1 0 6532 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _262_
timestamp 1666464484
transform 1 0 8740 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _263_
timestamp 1666464484
transform 1 0 10212 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _264_
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _265_
timestamp 1666464484
transform -1 0 14720 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _266_
timestamp 1666464484
transform 1 0 14352 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _267_
timestamp 1666464484
transform 1 0 13892 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _268_
timestamp 1666464484
transform 1 0 12880 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _269_
timestamp 1666464484
transform 1 0 14168 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_2  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1564 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _271_
timestamp 1666464484
transform -1 0 10396 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _272_
timestamp 1666464484
transform -1 0 5796 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _273_
timestamp 1666464484
transform 1 0 5244 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _274_
timestamp 1666464484
transform 1 0 4784 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _275_
timestamp 1666464484
transform -1 0 11960 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _276_
timestamp 1666464484
transform 1 0 7544 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _277_
timestamp 1666464484
transform 1 0 9476 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _278_
timestamp 1666464484
transform -1 0 12144 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _279_
timestamp 1666464484
transform -1 0 3036 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _280_
timestamp 1666464484
transform -1 0 8648 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_1  _281_
timestamp 1666464484
transform 1 0 3404 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _282_
timestamp 1666464484
transform 1 0 3128 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _283_
timestamp 1666464484
transform -1 0 6716 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _284_
timestamp 1666464484
transform 1 0 2760 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _285_
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _286_
timestamp 1666464484
transform 1 0 8096 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _287_
timestamp 1666464484
transform 1 0 6256 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _288_
timestamp 1666464484
transform 1 0 5336 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _289_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 13800 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _290_
timestamp 1666464484
transform -1 0 12788 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9016 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _292_
timestamp 1666464484
transform 1 0 6808 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _293_
timestamp 1666464484
transform -1 0 6440 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5888 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__069_
timestamp 1666464484
transform 1 0 9200 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__070_
timestamp 1666464484
transform 1 0 12144 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__071_
timestamp 1666464484
transform -1 0 10948 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__072_
timestamp 1666464484
transform -1 0 9844 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1666464484
transform 1 0 5244 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__068_
timestamp 1666464484
transform -1 0 3864 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__069_
timestamp 1666464484
transform -1 0 7084 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__070_
timestamp 1666464484
transform -1 0 12236 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__071_
timestamp 1666464484
transform -1 0 9660 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__072_
timestamp 1666464484
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1666464484
transform 1 0 6532 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__068_
timestamp 1666464484
transform 1 0 4232 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__069_
timestamp 1666464484
transform 1 0 11684 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__070_
timestamp 1666464484
transform 1 0 14260 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__071_
timestamp 1666464484
transform -1 0 9660 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__072_
timestamp 1666464484
transform 1 0 7820 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1666464484
transform 1 0 6532 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14260 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1666464484
transform -1 0 3036 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1666464484
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1666464484
transform -1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1666464484
transform -1 0 1932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1666464484
transform -1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1666464484
transform 1 0 1564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1666464484
transform 1 0 1564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1666464484
transform -1 0 1932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1666464484
transform -1 0 1932 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1666464484
transform -1 0 1932 0 -1 14144
box -38 -48 406 592
<< labels >>
flabel metal2 s 4434 17200 4490 18000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 io_out[0]
port 1 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 io_out[10]
port 2 nsew signal tristate
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 io_out[11]
port 3 nsew signal tristate
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 io_out[1]
port 4 nsew signal tristate
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 io_out[2]
port 5 nsew signal tristate
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 io_out[3]
port 6 nsew signal tristate
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 io_out[4]
port 7 nsew signal tristate
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 io_out[5]
port 8 nsew signal tristate
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 io_out[6]
port 9 nsew signal tristate
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 io_out[7]
port 10 nsew signal tristate
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 io_out[8]
port 11 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 io_out[9]
port 12 nsew signal tristate
flabel metal2 s 13450 17200 13506 18000 0 FreeSans 224 90 0 0 rst
port 13 nsew signal input
flabel metal4 s 2910 2128 3230 15824 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 6843 2128 7163 15824 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 10776 2128 11096 15824 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 14709 2128 15029 15824 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 4876 2128 5196 15824 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
flabel metal4 s 8809 2128 9129 15824 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
flabel metal4 s 12742 2128 13062 15824 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
flabel metal4 s 16675 2128 16995 15824 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
rlabel metal1 8970 15776 8970 15776 0 vccd1
rlabel via1 9049 15232 9049 15232 0 vssd1
rlabel metal2 12374 14246 12374 14246 0 CIRCUIT_1111.MEMORY_2.d
rlabel metal2 7406 14076 7406 14076 0 CIRCUIT_1111.MEMORY_2.s_currentState
rlabel metal1 7682 12886 7682 12886 0 CIRCUIT_1111.MEMORY_3.d
rlabel metal1 8648 13158 8648 13158 0 CIRCUIT_1111.MEMORY_3.s_currentState
rlabel metal1 6854 12818 6854 12818 0 CIRCUIT_1111.MEMORY_4.d
rlabel metal2 12466 11560 12466 11560 0 CIRCUIT_1111.MEMORY_6.d
rlabel metal2 13294 8126 13294 8126 0 CIRCUIT_1111.MEMORY_6.s_currentState
rlabel metal1 13340 9146 13340 9146 0 CIRCUIT_1111.MEMORY_7.d
rlabel metal1 13110 7412 13110 7412 0 CIRCUIT_1111.MEMORY_7.s_currentState
rlabel metal2 13294 14552 13294 14552 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_1.d
rlabel metal1 13018 15538 13018 15538 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_1.s_currentState
rlabel metal1 13892 10234 13892 10234 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_10.clock
rlabel metal2 15134 9316 15134 9316 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_10.d
rlabel metal1 15456 8942 15456 8942 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_10.s_currentState
rlabel metal2 8142 14756 8142 14756 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_2.d
rlabel metal2 8326 15198 8326 15198 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_2.s_currentState
rlabel metal2 9614 14756 9614 14756 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_3.d
rlabel metal1 10166 14926 10166 14926 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_3.s_currentState
rlabel metal1 11730 14042 11730 14042 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_4.d
rlabel metal2 11822 13702 11822 13702 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_4.s_currentState
rlabel metal1 11730 12886 11730 12886 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_5.d
rlabel metal1 12696 13158 12696 13158 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_5.s_currentState
rlabel metal1 13846 8058 13846 8058 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_6.d
rlabel metal1 13018 7854 13018 7854 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_6.s_currentState
rlabel metal2 13202 13294 13202 13294 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_7.clock
rlabel metal2 13294 11424 13294 11424 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_7.d
rlabel metal2 13386 11492 13386 11492 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_7.s_currentState
rlabel metal2 13570 10234 13570 10234 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_8.s_currentState
rlabel metal2 13662 13022 13662 13022 0 CIRCUIT_1111.custom_counter_10_1.MEMORY_9.s_currentState
rlabel metal1 1932 3706 1932 3706 0 CIRCUIT_1111.full_counter_1.ARITH_1.aEqualsB
rlabel metal2 13846 10744 13846 10744 0 CIRCUIT_1111.full_counter_1.ARITH_2.aEqualsB
rlabel metal1 5520 9554 5520 9554 0 CIRCUIT_1111.full_counter_1.MEMORY_3.s_currentState
rlabel metal1 6946 9588 6946 9588 0 CIRCUIT_1111.full_counter_1.MEMORY_6.s_currentState
rlabel metal1 3864 8398 3864 8398 0 CIRCUIT_1111.full_counter_1.custom_counter_4_1.MEMORY_1.d
rlabel metal1 4922 8330 4922 8330 0 CIRCUIT_1111.full_counter_1.custom_counter_4_1.MEMORY_1.s_currentState
rlabel metal1 6348 9010 6348 9010 0 CIRCUIT_1111.full_counter_1.custom_counter_4_1.MEMORY_2.d
rlabel metal1 2254 9452 2254 9452 0 CIRCUIT_1111.full_counter_1.custom_counter_4_1.MEMORY_2.s_currentState
rlabel metal1 3404 9622 3404 9622 0 CIRCUIT_1111.full_counter_1.custom_counter_4_1.MEMORY_3.d
rlabel metal1 2714 11084 2714 11084 0 CIRCUIT_1111.full_counter_1.custom_counter_4_1.MEMORY_3.s_currentState
rlabel metal1 3634 11662 3634 11662 0 CIRCUIT_1111.full_counter_1.custom_counter_4_1.MEMORY_4.d
rlabel metal1 6210 10030 6210 10030 0 CIRCUIT_1111.full_counter_1.custom_counter_4_1.MEMORY_4.s_currentState
rlabel metal1 4830 12614 4830 12614 0 CIRCUIT_1111.full_counter_1.custom_counter_4_2.MEMORY_1.d
rlabel metal1 5750 11730 5750 11730 0 CIRCUIT_1111.full_counter_1.custom_counter_4_2.MEMORY_1.s_currentState
rlabel metal1 7360 12614 7360 12614 0 CIRCUIT_1111.full_counter_1.custom_counter_4_2.MEMORY_2.d
rlabel metal1 7866 12818 7866 12818 0 CIRCUIT_1111.full_counter_1.custom_counter_4_2.MEMORY_2.s_currentState
rlabel metal1 8188 9486 8188 9486 0 CIRCUIT_1111.full_counter_1.custom_counter_4_2.MEMORY_3.d
rlabel metal1 9522 8976 9522 8976 0 CIRCUIT_1111.full_counter_1.custom_counter_4_2.MEMORY_3.s_currentState
rlabel metal2 10350 9724 10350 9724 0 CIRCUIT_1111.full_counter_1.custom_counter_4_2.MEMORY_4.d
rlabel metal1 11408 10642 11408 10642 0 CIRCUIT_1111.full_counter_1.custom_counter_4_2.MEMORY_4.s_currentState
rlabel metal2 10258 8024 10258 8024 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.ARITH_1.aEqualsB
rlabel metal1 3864 4794 3864 4794 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.ARITH_4.aEqualsB
rlabel metal1 10212 6290 10212 6290 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.MEMORY_5.s_currentState
rlabel metal2 2622 8636 2622 8636 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.MEMORY_6.s_currentState
rlabel metal2 10350 6358 10350 6358 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.custom_counter_4_1.MEMORY_1.d
rlabel metal1 9154 6358 9154 6358 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.custom_counter_4_1.MEMORY_1.s_currentState
rlabel metal1 7820 4182 7820 4182 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.custom_counter_4_1.MEMORY_2.d
rlabel metal2 9890 6834 9890 6834 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.custom_counter_4_1.MEMORY_2.s_currentState
rlabel metal2 9798 6630 9798 6630 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.custom_counter_4_1.MEMORY_3.d
rlabel metal2 11270 7174 11270 7174 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.custom_counter_4_1.MEMORY_3.s_currentState
rlabel metal2 11914 7650 11914 7650 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.custom_counter_4_1.MEMORY_4.d
rlabel metal1 10350 7752 10350 7752 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.custom_counter_4_1.MEMORY_4.s_currentState
rlabel metal2 5474 6936 5474 6936 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.custom_counter_4_2.MEMORY_1.d
rlabel metal1 5520 5202 5520 5202 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.custom_counter_4_2.MEMORY_1.s_currentState
rlabel metal2 5566 5202 5566 5202 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.custom_counter_4_2.MEMORY_2.d
rlabel metal1 3450 7446 3450 7446 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.custom_counter_4_2.MEMORY_2.s_currentState
rlabel metal1 5014 6834 5014 6834 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.custom_counter_4_2.MEMORY_3.d
rlabel metal2 3910 7514 3910 7514 0 CIRCUIT_1111.full_counter_1.seconds_counter_1.custom_counter_4_2.MEMORY_3.s_currentState
rlabel metal1 6486 14994 6486 14994 0 _007_
rlabel metal1 8786 15028 8786 15028 0 _009_
rlabel metal2 10258 14858 10258 14858 0 _011_
rlabel metal1 11132 13294 11132 13294 0 _013_
rlabel metal2 14674 8636 14674 8636 0 _015_
rlabel metal1 13846 13158 13846 13158 0 _017_
rlabel metal2 13938 11356 13938 11356 0 _019_
rlabel metal1 12926 12852 12926 12852 0 _021_
rlabel metal2 14214 9724 14214 9724 0 _023_
rlabel metal2 4462 6052 4462 6052 0 _026_
rlabel metal2 6670 5508 6670 5508 0 _027_
rlabel metal1 5290 5610 5290 5610 0 _028_
rlabel metal1 5888 8330 5888 8330 0 _029_
rlabel metal2 3818 7412 3818 7412 0 _030_
rlabel metal2 11178 6562 11178 6562 0 _031_
rlabel metal1 12374 6766 12374 6766 0 _032_
rlabel metal2 8510 4862 8510 4862 0 _033_
rlabel metal2 7590 4828 7590 4828 0 _034_
rlabel metal2 10534 5882 10534 5882 0 _035_
rlabel metal2 9522 5916 9522 5916 0 _036_
rlabel metal2 11362 8058 11362 8058 0 _037_
rlabel metal2 12098 8092 12098 8092 0 _038_
rlabel metal1 4508 11254 4508 11254 0 _041_
rlabel metal2 2714 11492 2714 11492 0 _042_
rlabel metal2 4462 9316 4462 9316 0 _043_
rlabel metal1 2346 9452 2346 9452 0 _044_
rlabel metal2 5934 9146 5934 9146 0 _045_
rlabel metal2 6670 9180 6670 9180 0 _046_
rlabel metal1 4140 7990 4140 7990 0 _047_
rlabel metal1 11224 9418 11224 9418 0 _048_
rlabel metal1 9844 8942 9844 8942 0 _049_
rlabel metal2 9430 9758 9430 9758 0 _050_
rlabel metal2 8142 10710 8142 10710 0 _051_
rlabel metal2 7314 12002 7314 12002 0 _052_
rlabel metal2 5934 12036 5934 12036 0 _053_
rlabel metal1 6486 9622 6486 9622 0 _054_
rlabel metal1 13110 9078 13110 9078 0 _056_
rlabel metal2 12558 12053 12558 12053 0 _058_
rlabel metal1 9062 12852 9062 12852 0 _060_
rlabel metal1 6808 13294 6808 13294 0 _062_
rlabel metal1 3312 5338 3312 5338 0 _064_
rlabel metal1 14628 12954 14628 12954 0 _065_
rlabel metal1 14766 13498 14766 13498 0 _066_
rlabel metal1 2898 14416 2898 14416 0 _067_
rlabel metal1 12834 14790 12834 14790 0 _068_
rlabel metal2 9246 11526 9246 11526 0 _069_
rlabel metal1 9476 11798 9476 11798 0 _070_
rlabel metal2 10258 11730 10258 11730 0 _071_
rlabel metal1 9568 8058 9568 8058 0 _072_
rlabel metal2 2346 13056 2346 13056 0 _073_
rlabel metal2 2070 15368 2070 15368 0 _074_
rlabel metal1 11914 15504 11914 15504 0 _075_
rlabel metal1 4140 14586 4140 14586 0 _076_
rlabel metal2 13938 14620 13938 14620 0 _077_
rlabel metal2 3174 12920 3174 12920 0 _078_
rlabel metal1 14214 12648 14214 12648 0 _079_
rlabel metal1 1656 11798 1656 11798 0 _080_
rlabel metal1 2070 11526 2070 11526 0 _081_
rlabel metal2 2070 3757 2070 3757 0 _082_
rlabel metal1 11454 11288 11454 11288 0 _083_
rlabel metal2 4186 5882 4186 5882 0 _084_
rlabel metal1 12535 7378 12535 7378 0 _085_
rlabel metal2 2714 6052 2714 6052 0 _086_
rlabel metal2 4370 5950 4370 5950 0 _087_
rlabel metal2 4002 4012 4002 4012 0 _088_
rlabel metal2 8602 6936 8602 6936 0 _089_
rlabel metal2 5198 7327 5198 7327 0 _090_
rlabel metal1 4416 6970 4416 6970 0 _091_
rlabel metal1 5934 7378 5934 7378 0 _092_
rlabel metal1 2806 7344 2806 7344 0 _093_
rlabel metal2 2806 4454 2806 4454 0 _094_
rlabel metal2 8234 7548 8234 7548 0 _095_
rlabel metal2 8418 8874 8418 8874 0 _096_
rlabel metal1 2714 4556 2714 4556 0 _097_
rlabel metal2 2070 5984 2070 5984 0 _098_
rlabel metal1 2530 7480 2530 7480 0 _099_
rlabel metal2 2714 4760 2714 4760 0 _100_
rlabel metal2 1794 4148 1794 4148 0 _101_
rlabel metal1 3220 4726 3220 4726 0 _102_
rlabel metal1 2714 5678 2714 5678 0 _103_
rlabel metal1 2208 5814 2208 5814 0 _104_
rlabel metal2 3450 4930 3450 4930 0 _105_
rlabel metal1 2300 7310 2300 7310 0 _106_
rlabel metal1 5014 14314 5014 14314 0 clk
rlabel metal2 4278 11424 4278 11424 0 clknet_0__068_
rlabel metal1 10488 11526 10488 11526 0 clknet_0__069_
rlabel metal1 13984 10030 13984 10030 0 clknet_0__070_
rlabel metal1 9660 13906 9660 13906 0 clknet_0__071_
rlabel metal1 7038 7888 7038 7888 0 clknet_0__072_
rlabel metal2 6578 14824 6578 14824 0 clknet_0_clk
rlabel metal1 15088 14246 15088 14246 0 clknet_1_0__leaf__068_
rlabel metal1 7452 7990 7452 7990 0 clknet_1_0__leaf__069_
rlabel metal1 13386 11220 13386 11220 0 clknet_1_0__leaf__070_
rlabel metal1 9338 10064 9338 10064 0 clknet_1_0__leaf__071_
rlabel metal1 4646 5712 4646 5712 0 clknet_1_0__leaf__072_
rlabel metal2 12466 14178 12466 14178 0 clknet_1_0__leaf_clk
rlabel metal1 14214 13872 14214 13872 0 clknet_1_1__leaf__068_
rlabel metal2 11178 10778 11178 10778 0 clknet_1_1__leaf__069_
rlabel metal1 15594 11118 15594 11118 0 clknet_1_1__leaf__070_
rlabel metal2 12558 15198 12558 15198 0 clknet_1_1__leaf__071_
rlabel metal1 10626 6324 10626 6324 0 clknet_1_1__leaf__072_
rlabel metal1 6946 13838 6946 13838 0 clknet_1_1__leaf_clk
rlabel metal3 1050 748 1050 748 0 io_out[0]
rlabel via2 2806 15691 2806 15691 0 io_out[10]
rlabel metal1 4646 15674 4646 15674 0 io_out[11]
rlabel metal3 1234 2244 1234 2244 0 io_out[1]
rlabel metal3 1050 3740 1050 3740 0 io_out[2]
rlabel metal1 1610 4726 1610 4726 0 io_out[3]
rlabel metal2 1702 6579 1702 6579 0 io_out[4]
rlabel metal2 1794 8143 1794 8143 0 io_out[5]
rlabel metal2 1794 9163 1794 9163 0 io_out[6]
rlabel metal3 1188 11220 1188 11220 0 io_out[7]
rlabel metal3 1188 12716 1188 12716 0 io_out[8]
rlabel metal2 1702 14127 1702 14127 0 io_out[9]
rlabel metal1 2208 11730 2208 11730 0 net1
rlabel metal1 1564 7514 1564 7514 0 net10
rlabel metal1 10718 12750 10718 12750 0 net11
rlabel metal2 2070 12614 2070 12614 0 net12
rlabel metal1 2162 13906 2162 13906 0 net13
rlabel metal1 3082 12342 3082 12342 0 net14
rlabel metal1 10074 14824 10074 14824 0 net15
rlabel metal1 5014 15062 5014 15062 0 net16
rlabel metal1 7866 14416 7866 14416 0 net17
rlabel metal2 13846 13328 13846 13328 0 net18
rlabel metal2 1610 7412 1610 7412 0 net19
rlabel metal2 1886 3468 1886 3468 0 net2
rlabel metal1 10258 13838 10258 13838 0 net20
rlabel metal2 3542 6528 3542 6528 0 net21
rlabel metal2 9246 7888 9246 7888 0 net22
rlabel metal1 8234 13369 8234 13369 0 net23
rlabel metal1 10764 13838 10764 13838 0 net24
rlabel metal1 12650 11016 12650 11016 0 net25
rlabel metal2 16238 10064 16238 10064 0 net26
rlabel metal2 15502 9112 15502 9112 0 net27
rlabel metal1 14352 13158 14352 13158 0 net28
rlabel metal2 15686 10880 15686 10880 0 net29
rlabel metal1 2530 14892 2530 14892 0 net3
rlabel metal1 14759 11798 14759 11798 0 net30
rlabel metal1 14911 8534 14911 8534 0 net31
rlabel metal2 12558 13770 12558 13770 0 net32
rlabel metal1 11783 14314 11783 14314 0 net33
rlabel metal2 10994 15198 10994 15198 0 net34
rlabel metal2 8694 15232 8694 15232 0 net35
rlabel metal2 13202 14110 13202 14110 0 net36
rlabel metal2 5658 14008 5658 14008 0 net37
rlabel metal2 2438 15266 2438 15266 0 net4
rlabel metal1 1656 2414 1656 2414 0 net5
rlabel metal2 1886 4284 1886 4284 0 net6
rlabel metal2 1886 5066 1886 5066 0 net7
rlabel metal2 1886 6460 1886 6460 0 net8
rlabel metal1 1656 6970 1656 6970 0 net9
rlabel metal1 6302 12818 6302 12818 0 prev_sel
rlabel metal2 13623 17340 13623 17340 0 rst
<< properties >>
string FIXED_BBOX 0 0 18000 18000
<< end >>
