magic
tech sky130B
magscale 1 2
timestamp 1682098768
<< viali >>
rect 1593 18717 1627 18751
rect 1869 18649 1903 18683
rect 4353 17153 4387 17187
rect 4445 17153 4479 17187
rect 6561 17153 6595 17187
rect 6745 17153 6779 17187
rect 7757 17153 7791 17187
rect 7941 17153 7975 17187
rect 4629 17085 4663 17119
rect 4537 16949 4571 16983
rect 6561 16949 6595 16983
rect 7849 16949 7883 16983
rect 7021 16677 7055 16711
rect 4629 16609 4663 16643
rect 6101 16609 6135 16643
rect 6193 16609 6227 16643
rect 6285 16609 6319 16643
rect 6377 16609 6411 16643
rect 7757 16609 7791 16643
rect 3341 16541 3375 16575
rect 3433 16541 3467 16575
rect 4813 16541 4847 16575
rect 7573 16541 7607 16575
rect 8401 16541 8435 16575
rect 10977 16541 11011 16575
rect 14749 16541 14783 16575
rect 14933 16541 14967 16575
rect 3157 16473 3191 16507
rect 7021 16473 7055 16507
rect 8217 16473 8251 16507
rect 8585 16473 8619 16507
rect 11253 16473 11287 16507
rect 3249 16405 3283 16439
rect 4997 16405 5031 16439
rect 5917 16405 5951 16439
rect 7481 16405 7515 16439
rect 14841 16405 14875 16439
rect 9689 16133 9723 16167
rect 12909 16133 12943 16167
rect 3709 16065 3743 16099
rect 4629 16065 4663 16099
rect 4721 16065 4755 16099
rect 4905 16065 4939 16099
rect 4997 16065 5031 16099
rect 5457 16065 5491 16099
rect 5641 16065 5675 16099
rect 6561 16065 6595 16099
rect 7481 16065 7515 16099
rect 7757 16065 7791 16099
rect 9413 16065 9447 16099
rect 10333 16065 10367 16099
rect 12081 16065 12115 16099
rect 13093 16065 13127 16099
rect 13185 16065 13219 16099
rect 13369 16065 13403 16099
rect 13461 16065 13495 16099
rect 14565 16065 14599 16099
rect 14658 16065 14692 16099
rect 14841 16065 14875 16099
rect 14933 16065 14967 16099
rect 15071 16065 15105 16099
rect 16037 16065 16071 16099
rect 3985 15997 4019 16031
rect 4445 15997 4479 16031
rect 6653 15997 6687 16031
rect 6837 15997 6871 16031
rect 7849 15997 7883 16031
rect 9321 15997 9355 16031
rect 9781 15997 9815 16031
rect 12173 15997 12207 16031
rect 12265 15997 12299 16031
rect 15853 15997 15887 16031
rect 15945 15997 15979 16031
rect 16129 15997 16163 16031
rect 5549 15929 5583 15963
rect 7573 15929 7607 15963
rect 15209 15929 15243 15963
rect 3801 15861 3835 15895
rect 3893 15861 3927 15895
rect 6745 15861 6779 15895
rect 7665 15861 7699 15895
rect 9137 15861 9171 15895
rect 10517 15861 10551 15895
rect 11713 15861 11747 15895
rect 15669 15861 15703 15895
rect 9229 15657 9263 15691
rect 10425 15657 10459 15691
rect 10885 15657 10919 15691
rect 14565 15657 14599 15691
rect 16037 15657 16071 15691
rect 17049 15657 17083 15691
rect 7757 15589 7791 15623
rect 12633 15589 12667 15623
rect 13369 15589 13403 15623
rect 2605 15521 2639 15555
rect 12817 15521 12851 15555
rect 2421 15453 2455 15487
rect 7573 15453 7607 15487
rect 7757 15453 7791 15487
rect 9505 15453 9539 15487
rect 10609 15453 10643 15487
rect 10701 15453 10735 15487
rect 10977 15453 11011 15487
rect 11437 15453 11471 15487
rect 11529 15453 11563 15487
rect 12542 15453 12576 15487
rect 13277 15453 13311 15487
rect 13461 15453 13495 15487
rect 14473 15453 14507 15487
rect 14657 15453 14691 15487
rect 16221 15453 16255 15487
rect 16313 15453 16347 15487
rect 16497 15453 16531 15487
rect 16589 15453 16623 15487
rect 17325 15453 17359 15487
rect 17417 15453 17451 15487
rect 17509 15453 17543 15487
rect 17693 15453 17727 15487
rect 9229 15385 9263 15419
rect 12817 15385 12851 15419
rect 1961 15317 1995 15351
rect 2329 15317 2363 15351
rect 9413 15317 9447 15351
rect 8217 15113 8251 15147
rect 14657 15113 14691 15147
rect 16221 15113 16255 15147
rect 17509 15113 17543 15147
rect 18153 15113 18187 15147
rect 7113 15045 7147 15079
rect 7297 15045 7331 15079
rect 13277 15045 13311 15079
rect 15853 15045 15887 15079
rect 16069 15045 16103 15079
rect 18889 15045 18923 15079
rect 2329 14977 2363 15011
rect 2513 14977 2547 15011
rect 7941 14977 7975 15011
rect 11897 14977 11931 15011
rect 11989 14977 12023 15011
rect 12173 14977 12207 15011
rect 12265 14977 12299 15011
rect 13185 14977 13219 15011
rect 14565 14977 14599 15011
rect 14749 14977 14783 15011
rect 18245 14977 18279 15011
rect 18705 14977 18739 15011
rect 18981 14977 19015 15011
rect 8217 14909 8251 14943
rect 13369 14909 13403 14943
rect 17785 14909 17819 14943
rect 12817 14841 12851 14875
rect 18705 14841 18739 14875
rect 2421 14773 2455 14807
rect 7481 14773 7515 14807
rect 8033 14773 8067 14807
rect 11713 14773 11747 14807
rect 16037 14773 16071 14807
rect 17877 14773 17911 14807
rect 17969 14773 18003 14807
rect 7573 14569 7607 14603
rect 8217 14569 8251 14603
rect 12449 14569 12483 14603
rect 15577 14569 15611 14603
rect 9137 14501 9171 14535
rect 16497 14501 16531 14535
rect 4537 14433 4571 14467
rect 6101 14433 6135 14467
rect 7297 14433 7331 14467
rect 9781 14433 9815 14467
rect 10241 14433 10275 14467
rect 11989 14433 12023 14467
rect 18521 14433 18555 14467
rect 2973 14365 3007 14399
rect 3065 14365 3099 14399
rect 3341 14365 3375 14399
rect 3433 14365 3467 14399
rect 4169 14365 4203 14399
rect 4261 14365 4295 14399
rect 4353 14365 4387 14399
rect 4997 14365 5031 14399
rect 5365 14365 5399 14399
rect 6009 14365 6043 14399
rect 6193 14365 6227 14399
rect 7389 14365 7423 14399
rect 9262 14365 9296 14399
rect 9689 14365 9723 14399
rect 10517 14365 10551 14399
rect 10609 14365 10643 14399
rect 10701 14365 10735 14399
rect 10885 14365 10919 14399
rect 11713 14365 11747 14399
rect 11897 14365 11931 14399
rect 12081 14365 12115 14399
rect 12265 14365 12299 14399
rect 13369 14365 13403 14399
rect 13645 14365 13679 14399
rect 15485 14365 15519 14399
rect 15853 14365 15887 14399
rect 16497 14365 16531 14399
rect 16681 14365 16715 14399
rect 18245 14365 18279 14399
rect 18337 14365 18371 14399
rect 1961 14297 1995 14331
rect 2145 14297 2179 14331
rect 3157 14297 3191 14331
rect 5181 14297 5215 14331
rect 5273 14297 5307 14331
rect 8125 14297 8159 14331
rect 2329 14229 2363 14263
rect 2789 14229 2823 14263
rect 5549 14229 5583 14263
rect 6929 14229 6963 14263
rect 9321 14229 9355 14263
rect 13185 14229 13219 14263
rect 13553 14229 13587 14263
rect 16037 14229 16071 14263
rect 18521 14229 18555 14263
rect 2053 14025 2087 14059
rect 2979 14025 3013 14059
rect 5365 14025 5399 14059
rect 9321 14025 9355 14059
rect 11897 14025 11931 14059
rect 15761 14025 15795 14059
rect 17325 14025 17359 14059
rect 19441 14025 19475 14059
rect 19625 14025 19659 14059
rect 3065 13957 3099 13991
rect 6930 13957 6964 13991
rect 9873 13957 9907 13991
rect 10425 13957 10459 13991
rect 14013 13957 14047 13991
rect 15393 13957 15427 13991
rect 16865 13957 16899 13991
rect 1961 13889 1995 13923
rect 2881 13889 2915 13923
rect 3157 13889 3191 13923
rect 4997 13889 5031 13923
rect 5181 13889 5215 13923
rect 6838 13911 6872 13945
rect 7021 13889 7055 13923
rect 7159 13889 7193 13923
rect 7849 13889 7883 13923
rect 8033 13889 8067 13923
rect 8953 13889 8987 13923
rect 10057 13889 10091 13923
rect 12909 13889 12943 13923
rect 14289 13889 14323 13923
rect 14749 13889 14783 13923
rect 15209 13889 15243 13923
rect 15485 13889 15519 13923
rect 15577 13889 15611 13923
rect 18337 13889 18371 13923
rect 18429 13889 18463 13923
rect 18649 13889 18683 13923
rect 19566 13889 19600 13923
rect 2237 13821 2271 13855
rect 6653 13821 6687 13855
rect 7297 13821 7331 13855
rect 8861 13821 8895 13855
rect 11713 13821 11747 13855
rect 12173 13821 12207 13855
rect 12265 13821 12299 13855
rect 14381 13821 14415 13855
rect 18521 13821 18555 13855
rect 20085 13821 20119 13855
rect 7849 13753 7883 13787
rect 14473 13753 14507 13787
rect 17141 13753 17175 13787
rect 19993 13753 20027 13787
rect 1593 13685 1627 13719
rect 13093 13685 13127 13719
rect 14565 13685 14599 13719
rect 18153 13685 18187 13719
rect 7573 13481 7607 13515
rect 9229 13481 9263 13515
rect 13553 13481 13587 13515
rect 14289 13481 14323 13515
rect 17509 13481 17543 13515
rect 11621 13413 11655 13447
rect 4721 13345 4755 13379
rect 4905 13345 4939 13379
rect 18153 13345 18187 13379
rect 2237 13277 2271 13311
rect 7481 13277 7515 13311
rect 9137 13277 9171 13311
rect 9321 13277 9355 13311
rect 11253 13277 11287 13311
rect 11407 13277 11441 13311
rect 13461 13277 13495 13311
rect 14289 13277 14323 13311
rect 14473 13277 14507 13311
rect 17693 13277 17727 13311
rect 17785 13277 17819 13311
rect 18061 13277 18095 13311
rect 19901 13277 19935 13311
rect 2697 13209 2731 13243
rect 19993 13209 20027 13243
rect 4261 13141 4295 13175
rect 4629 13141 4663 13175
rect 4169 12937 4203 12971
rect 5365 12937 5399 12971
rect 6837 12937 6871 12971
rect 15853 12937 15887 12971
rect 16865 12937 16899 12971
rect 18613 12937 18647 12971
rect 20085 12937 20119 12971
rect 2513 12801 2547 12835
rect 4077 12801 4111 12835
rect 5273 12801 5307 12835
rect 6653 12801 6687 12835
rect 7021 12801 7055 12835
rect 7205 12801 7239 12835
rect 9045 12801 9079 12835
rect 11713 12801 11747 12835
rect 13369 12801 13403 12835
rect 15761 12801 15795 12835
rect 16037 12801 16071 12835
rect 17141 12801 17175 12835
rect 17233 12801 17267 12835
rect 18429 12801 18463 12835
rect 18705 12801 18739 12835
rect 19717 12801 19751 12835
rect 19901 12801 19935 12835
rect 3065 12733 3099 12767
rect 4261 12733 4295 12767
rect 5457 12733 5491 12767
rect 8953 12733 8987 12767
rect 9137 12733 9171 12767
rect 9229 12733 9263 12767
rect 11989 12733 12023 12767
rect 13553 12733 13587 12767
rect 17049 12733 17083 12767
rect 17325 12733 17359 12767
rect 11805 12665 11839 12699
rect 18429 12665 18463 12699
rect 3709 12597 3743 12631
rect 4905 12597 4939 12631
rect 7021 12597 7055 12631
rect 8769 12597 8803 12631
rect 11713 12597 11747 12631
rect 19717 12597 19751 12631
rect 9137 12393 9171 12427
rect 11253 12393 11287 12427
rect 11805 12393 11839 12427
rect 14841 12393 14875 12427
rect 15393 12393 15427 12427
rect 17601 12393 17635 12427
rect 19717 12393 19751 12427
rect 20085 12325 20119 12359
rect 2329 12257 2363 12291
rect 2513 12257 2547 12291
rect 3157 12257 3191 12291
rect 3341 12257 3375 12291
rect 5273 12257 5307 12291
rect 5457 12257 5491 12291
rect 7297 12257 7331 12291
rect 12173 12257 12207 12291
rect 14381 12257 14415 12291
rect 16589 12257 16623 12291
rect 19809 12257 19843 12291
rect 3065 12189 3099 12223
rect 6377 12189 6411 12223
rect 6745 12189 6779 12223
rect 7113 12189 7147 12223
rect 7849 12189 7883 12223
rect 8309 12189 8343 12223
rect 8585 12189 8619 12223
rect 9321 12189 9355 12223
rect 9413 12189 9447 12223
rect 10891 12189 10925 12223
rect 11345 12189 11379 12223
rect 11989 12189 12023 12223
rect 12081 12189 12115 12223
rect 12265 12189 12299 12223
rect 13093 12189 13127 12223
rect 13277 12189 13311 12223
rect 14565 12189 14599 12223
rect 14657 12189 14691 12223
rect 14933 12189 14967 12223
rect 15393 12189 15427 12223
rect 15577 12189 15611 12223
rect 16313 12189 16347 12223
rect 17857 12189 17891 12223
rect 17966 12189 18000 12223
rect 18061 12189 18095 12223
rect 18245 12189 18279 12223
rect 19717 12189 19751 12223
rect 8493 12121 8527 12155
rect 9689 12121 9723 12155
rect 9781 12121 9815 12155
rect 10977 12121 11011 12155
rect 11069 12121 11103 12155
rect 16129 12121 16163 12155
rect 1869 12053 1903 12087
rect 2237 12053 2271 12087
rect 3341 12053 3375 12087
rect 4813 12053 4847 12087
rect 5181 12053 5215 12087
rect 8407 12053 8441 12087
rect 10609 12053 10643 12087
rect 13461 12053 13495 12087
rect 2421 11849 2455 11883
rect 2881 11849 2915 11883
rect 7573 11849 7607 11883
rect 12173 11849 12207 11883
rect 12357 11849 12391 11883
rect 13553 11849 13587 11883
rect 19257 11849 19291 11883
rect 20085 11849 20119 11883
rect 4537 11781 4571 11815
rect 8861 11781 8895 11815
rect 9413 11781 9447 11815
rect 14197 11781 14231 11815
rect 15945 11781 15979 11815
rect 19809 11781 19843 11815
rect 2237 11713 2271 11747
rect 3249 11713 3283 11747
rect 4261 11713 4295 11747
rect 4445 11713 4479 11747
rect 4629 11713 4663 11747
rect 5457 11713 5491 11747
rect 7481 11713 7515 11747
rect 9045 11713 9079 11747
rect 10517 11713 10551 11747
rect 10701 11713 10735 11747
rect 10793 11713 10827 11747
rect 11989 11713 12023 11747
rect 12081 11713 12115 11747
rect 13369 11713 13403 11747
rect 13645 11713 13679 11747
rect 14105 11713 14139 11747
rect 14289 11713 14323 11747
rect 15025 11713 15059 11747
rect 15209 11713 15243 11747
rect 15669 11713 15703 11747
rect 15762 11713 15796 11747
rect 16037 11713 16071 11747
rect 16134 11713 16168 11747
rect 17509 11713 17543 11747
rect 18613 11713 18647 11747
rect 19993 11713 20027 11747
rect 2053 11645 2087 11679
rect 3341 11645 3375 11679
rect 5273 11645 5307 11679
rect 5733 11645 5767 11679
rect 7665 11645 7699 11679
rect 10609 11645 10643 11679
rect 17325 11645 17359 11679
rect 18981 11645 19015 11679
rect 5641 11577 5675 11611
rect 11805 11577 11839 11611
rect 18778 11577 18812 11611
rect 3525 11509 3559 11543
rect 4813 11509 4847 11543
rect 7113 11509 7147 11543
rect 10333 11509 10367 11543
rect 13369 11509 13403 11543
rect 15025 11509 15059 11543
rect 16313 11509 16347 11543
rect 17693 11509 17727 11543
rect 18889 11509 18923 11543
rect 12449 11305 12483 11339
rect 14657 11305 14691 11339
rect 16129 11305 16163 11339
rect 1869 11237 1903 11271
rect 6745 11237 6779 11271
rect 14289 11237 14323 11271
rect 16037 11237 16071 11271
rect 4169 11169 4203 11203
rect 7205 11169 7239 11203
rect 7389 11169 7423 11203
rect 16221 11169 16255 11203
rect 19533 11169 19567 11203
rect 20177 11169 20211 11203
rect 1869 11101 1903 11135
rect 2145 11101 2179 11135
rect 3985 11101 4019 11135
rect 12357 11101 12391 11135
rect 13553 11101 13587 11135
rect 15945 11101 15979 11135
rect 17601 11101 17635 11135
rect 19441 11101 19475 11135
rect 19717 11101 19751 11135
rect 2053 11033 2087 11067
rect 7113 11033 7147 11067
rect 13645 11033 13679 11067
rect 14657 11033 14691 11067
rect 14841 10965 14875 10999
rect 17693 10965 17727 10999
rect 19625 10761 19659 10795
rect 1685 10693 1719 10727
rect 1869 10693 1903 10727
rect 10048 10693 10082 10727
rect 18429 10693 18463 10727
rect 8024 10625 8058 10659
rect 13829 10625 13863 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 18613 10625 18647 10659
rect 19625 10625 19659 10659
rect 19993 10625 20027 10659
rect 7757 10557 7791 10591
rect 9781 10557 9815 10591
rect 13921 10557 13955 10591
rect 19441 10557 19475 10591
rect 9137 10489 9171 10523
rect 11161 10421 11195 10455
rect 14013 10421 14047 10455
rect 14197 10421 14231 10455
rect 16957 10421 16991 10455
rect 18705 10421 18739 10455
rect 2973 10217 3007 10251
rect 8401 10217 8435 10251
rect 11621 10217 11655 10251
rect 16681 10217 16715 10251
rect 19625 10217 19659 10251
rect 12955 10149 12989 10183
rect 15669 10149 15703 10183
rect 15761 10149 15795 10183
rect 16865 10149 16899 10183
rect 19809 10149 19843 10183
rect 10333 10081 10367 10115
rect 14565 10081 14599 10115
rect 14657 10081 14691 10115
rect 1593 10013 1627 10047
rect 1860 10013 1894 10047
rect 5089 10013 5123 10047
rect 5356 10013 5390 10047
rect 7021 10013 7055 10047
rect 7277 10013 7311 10047
rect 10057 10013 10091 10047
rect 12817 10013 12851 10047
rect 13093 10013 13127 10047
rect 13277 10013 13311 10047
rect 14473 10013 14507 10047
rect 14749 10013 14783 10047
rect 15393 10013 15427 10047
rect 15577 10013 15611 10047
rect 15853 10013 15887 10047
rect 16037 10013 16071 10047
rect 17417 10013 17451 10047
rect 17877 10013 17911 10047
rect 18061 10013 18095 10047
rect 13185 9945 13219 9979
rect 16497 9945 16531 9979
rect 16697 9945 16731 9979
rect 19441 9945 19475 9979
rect 19641 9945 19675 9979
rect 6469 9877 6503 9911
rect 14289 9877 14323 9911
rect 17601 9877 17635 9911
rect 13093 9673 13127 9707
rect 3056 9605 3090 9639
rect 15485 9605 15519 9639
rect 16865 9605 16899 9639
rect 8033 9537 8067 9571
rect 13001 9537 13035 9571
rect 13185 9537 13219 9571
rect 14289 9537 14323 9571
rect 14473 9537 14507 9571
rect 15117 9537 15151 9571
rect 15301 9537 15335 9571
rect 16129 9537 16163 9571
rect 17049 9537 17083 9571
rect 17141 9537 17175 9571
rect 18521 9537 18555 9571
rect 18889 9537 18923 9571
rect 2789 9469 2823 9503
rect 7757 9469 7791 9503
rect 4169 9401 4203 9435
rect 16865 9401 16899 9435
rect 19717 9401 19751 9435
rect 9137 9333 9171 9367
rect 14381 9333 14415 9367
rect 16221 9333 16255 9367
rect 2973 9129 3007 9163
rect 6009 9129 6043 9163
rect 8493 9129 8527 9163
rect 11713 9129 11747 9163
rect 17877 9129 17911 9163
rect 19901 9129 19935 9163
rect 19717 9061 19751 9095
rect 1593 8993 1627 9027
rect 7113 8993 7147 9027
rect 10425 8993 10459 9027
rect 19441 8993 19475 9027
rect 1860 8925 1894 8959
rect 4629 8925 4663 8959
rect 4896 8925 4930 8959
rect 7380 8925 7414 8959
rect 10149 8925 10183 8959
rect 14381 8925 14415 8959
rect 16589 8925 16623 8959
rect 16957 8925 16991 8959
rect 17049 8925 17083 8959
rect 17417 8925 17451 8959
rect 17509 8925 17543 8959
rect 14565 8857 14599 8891
rect 14749 8789 14783 8823
rect 4353 8585 4387 8619
rect 11161 8585 11195 8619
rect 18245 8585 18279 8619
rect 3240 8517 3274 8551
rect 10048 8517 10082 8551
rect 14197 8517 14231 8551
rect 17233 8517 17267 8551
rect 18521 8517 18555 8551
rect 13185 8449 13219 8483
rect 13369 8449 13403 8483
rect 14013 8449 14047 8483
rect 14105 8449 14139 8483
rect 14335 8449 14369 8483
rect 16865 8449 16899 8483
rect 17049 8449 17083 8483
rect 18429 8449 18463 8483
rect 18613 8449 18647 8483
rect 18797 8449 18831 8483
rect 18889 8449 18923 8483
rect 2973 8381 3007 8415
rect 9781 8381 9815 8415
rect 14473 8381 14507 8415
rect 13277 8313 13311 8347
rect 13829 8245 13863 8279
rect 6193 8041 6227 8075
rect 8401 8041 8435 8075
rect 11345 8041 11379 8075
rect 15577 8041 15611 8075
rect 16957 8041 16991 8075
rect 7021 7905 7055 7939
rect 9965 7905 9999 7939
rect 13277 7905 13311 7939
rect 17601 7905 17635 7939
rect 18613 7905 18647 7939
rect 4813 7837 4847 7871
rect 7288 7837 7322 7871
rect 13093 7837 13127 7871
rect 15209 7837 15243 7871
rect 15577 7837 15611 7871
rect 16865 7837 16899 7871
rect 17049 7837 17083 7871
rect 17509 7837 17543 7871
rect 18521 7837 18555 7871
rect 18705 7837 18739 7871
rect 18797 7837 18831 7871
rect 19441 7837 19475 7871
rect 19625 7837 19659 7871
rect 5080 7769 5114 7803
rect 10232 7769 10266 7803
rect 12633 7701 12667 7735
rect 13001 7701 13035 7735
rect 15393 7701 15427 7735
rect 18337 7701 18371 7735
rect 19533 7701 19567 7735
rect 9137 7497 9171 7531
rect 17785 7497 17819 7531
rect 2605 7361 2639 7395
rect 7849 7361 7883 7395
rect 13001 7361 13035 7395
rect 13093 7361 13127 7395
rect 15209 7361 15243 7395
rect 17693 7361 17727 7395
rect 13185 7293 13219 7327
rect 15301 7293 15335 7327
rect 15485 7293 15519 7327
rect 3893 7157 3927 7191
rect 12633 7157 12667 7191
rect 14841 7157 14875 7191
rect 14289 6953 14323 6987
rect 15485 6953 15519 6987
rect 17417 6953 17451 6987
rect 7297 6885 7331 6919
rect 15945 6885 15979 6919
rect 9781 6817 9815 6851
rect 17325 6817 17359 6851
rect 1593 6749 1627 6783
rect 1849 6749 1883 6783
rect 10048 6749 10082 6783
rect 13461 6749 13495 6783
rect 13645 6749 13679 6783
rect 13737 6749 13771 6783
rect 14473 6749 14507 6783
rect 14565 6749 14599 6783
rect 15669 6749 15703 6783
rect 15761 6749 15795 6783
rect 16037 6749 16071 6783
rect 17141 6749 17175 6783
rect 17417 6749 17451 6783
rect 18245 6749 18279 6783
rect 18613 6749 18647 6783
rect 18705 6749 18739 6783
rect 6009 6681 6043 6715
rect 14841 6681 14875 6715
rect 14933 6681 14967 6715
rect 2973 6613 3007 6647
rect 11161 6613 11195 6647
rect 13277 6613 13311 6647
rect 17601 6613 17635 6647
rect 18337 6613 18371 6647
rect 4169 6409 4203 6443
rect 8493 6409 8527 6443
rect 13001 6409 13035 6443
rect 14841 6409 14875 6443
rect 17049 6409 17083 6443
rect 18337 6409 18371 6443
rect 3056 6341 3090 6375
rect 12909 6341 12943 6375
rect 14473 6341 14507 6375
rect 2789 6273 2823 6307
rect 7380 6273 7414 6307
rect 8953 6273 8987 6307
rect 9220 6273 9254 6307
rect 14657 6273 14691 6307
rect 16037 6273 16071 6307
rect 17233 6273 17267 6307
rect 17509 6273 17543 6307
rect 18521 6273 18555 6307
rect 18797 6273 18831 6307
rect 18981 6273 19015 6307
rect 7113 6205 7147 6239
rect 13185 6205 13219 6239
rect 15853 6205 15887 6239
rect 12541 6137 12575 6171
rect 10333 6069 10367 6103
rect 16221 6069 16255 6103
rect 6745 5865 6779 5899
rect 11161 5865 11195 5899
rect 14381 5865 14415 5899
rect 19717 5797 19751 5831
rect 1593 5729 1627 5763
rect 16681 5729 16715 5763
rect 1869 5661 1903 5695
rect 5365 5661 5399 5695
rect 9781 5661 9815 5695
rect 14657 5661 14691 5695
rect 17325 5661 17359 5695
rect 17509 5661 17543 5695
rect 19441 5661 19475 5695
rect 19625 5661 19659 5695
rect 5632 5593 5666 5627
rect 10048 5593 10082 5627
rect 14381 5593 14415 5627
rect 3157 5525 3191 5559
rect 14565 5525 14599 5559
rect 16129 5525 16163 5559
rect 16497 5525 16531 5559
rect 16589 5525 16623 5559
rect 17417 5525 17451 5559
rect 17049 5321 17083 5355
rect 10048 5253 10082 5287
rect 2513 5185 2547 5219
rect 3913 5185 3947 5219
rect 4169 5185 4203 5219
rect 4629 5185 4663 5219
rect 4896 5185 4930 5219
rect 12909 5185 12943 5219
rect 13829 5185 13863 5219
rect 14381 5185 14415 5219
rect 15209 5185 15243 5219
rect 15301 5185 15335 5219
rect 15393 5185 15427 5219
rect 15577 5185 15611 5219
rect 16957 5185 16991 5219
rect 9781 5117 9815 5151
rect 13001 5117 13035 5151
rect 13185 5117 13219 5151
rect 2789 5049 2823 5083
rect 11161 5049 11195 5083
rect 14933 5049 14967 5083
rect 6009 4981 6043 5015
rect 12541 4981 12575 5015
rect 16957 4709 16991 4743
rect 2053 4641 2087 4675
rect 5273 4641 5307 4675
rect 7113 4641 7147 4675
rect 15669 4641 15703 4675
rect 17141 4641 17175 4675
rect 5540 4573 5574 4607
rect 9781 4573 9815 4607
rect 10048 4573 10082 4607
rect 13553 4573 13587 4607
rect 13645 4573 13679 4607
rect 14473 4573 14507 4607
rect 14657 4573 14691 4607
rect 14750 4551 14784 4585
rect 14875 4573 14909 4607
rect 15577 4573 15611 4607
rect 17233 4573 17267 4607
rect 18061 4573 18095 4607
rect 2320 4505 2354 4539
rect 7380 4505 7414 4539
rect 15117 4505 15151 4539
rect 17509 4505 17543 4539
rect 17601 4505 17635 4539
rect 18153 4505 18187 4539
rect 3433 4437 3467 4471
rect 6653 4437 6687 4471
rect 8493 4437 8527 4471
rect 11161 4437 11195 4471
rect 17049 4233 17083 4267
rect 1593 4097 1627 4131
rect 1860 4097 1894 4131
rect 4537 4097 4571 4131
rect 4804 4097 4838 4131
rect 7113 4097 7147 4131
rect 7380 4097 7414 4131
rect 9864 4097 9898 4131
rect 14197 4097 14231 4131
rect 14381 4097 14415 4131
rect 14657 4097 14691 4131
rect 14841 4097 14875 4131
rect 15025 4097 15059 4131
rect 16865 4097 16899 4131
rect 17233 4097 17267 4131
rect 17417 4097 17451 4131
rect 9597 4029 9631 4063
rect 2973 3893 3007 3927
rect 5917 3893 5951 3927
rect 8493 3893 8527 3927
rect 10977 3893 11011 3927
rect 17233 3893 17267 3927
rect 13001 3689 13035 3723
rect 14289 3689 14323 3723
rect 17233 3689 17267 3723
rect 18245 3689 18279 3723
rect 11069 3621 11103 3655
rect 11805 3621 11839 3655
rect 16773 3621 16807 3655
rect 2053 3553 2087 3587
rect 13461 3553 13495 3587
rect 14565 3553 14599 3587
rect 7021 3485 7055 3519
rect 9689 3485 9723 3519
rect 9956 3485 9990 3519
rect 11805 3485 11839 3519
rect 11989 3485 12023 3519
rect 12081 3485 12115 3519
rect 13185 3485 13219 3519
rect 13369 3485 13403 3519
rect 14473 3485 14507 3519
rect 14933 3485 14967 3519
rect 16957 3485 16991 3519
rect 17049 3485 17083 3519
rect 17325 3485 17359 3519
rect 17969 3485 18003 3519
rect 18061 3485 18095 3519
rect 18337 3485 18371 3519
rect 2320 3417 2354 3451
rect 7288 3417 7322 3451
rect 14841 3417 14875 3451
rect 3433 3349 3467 3383
rect 8401 3349 8435 3383
rect 14657 3349 14691 3383
rect 17785 3349 17819 3383
rect 1869 3145 1903 3179
rect 5549 3145 5583 3179
rect 10057 3145 10091 3179
rect 13645 3145 13679 3179
rect 14197 3145 14231 3179
rect 16221 3145 16255 3179
rect 2605 3077 2639 3111
rect 4353 3077 4387 3111
rect 4813 3077 4847 3111
rect 6837 3077 6871 3111
rect 6929 3077 6963 3111
rect 7849 3077 7883 3111
rect 9597 3077 9631 3111
rect 15853 3077 15887 3111
rect 16069 3077 16103 3111
rect 1777 3009 1811 3043
rect 1961 3009 1995 3043
rect 4997 3009 5031 3043
rect 5089 3009 5123 3043
rect 5733 3009 5767 3043
rect 6009 3009 6043 3043
rect 6745 3009 6779 3043
rect 10241 3009 10275 3043
rect 12541 3009 12575 3043
rect 12725 3009 12759 3043
rect 13461 3009 13495 3043
rect 14105 3009 14139 3043
rect 14289 3009 14323 3043
rect 14933 3009 14967 3043
rect 15209 3009 15243 3043
rect 15393 3009 15427 3043
rect 17049 3009 17083 3043
rect 6561 2941 6595 2975
rect 7297 2941 7331 2975
rect 10517 2941 10551 2975
rect 12357 2941 12391 2975
rect 13277 2941 13311 2975
rect 17141 2941 17175 2975
rect 17417 2941 17451 2975
rect 14749 2873 14783 2907
rect 4813 2805 4847 2839
rect 5917 2805 5951 2839
rect 10425 2805 10459 2839
rect 16037 2805 16071 2839
rect 2973 2601 3007 2635
rect 3341 2601 3375 2635
rect 3985 2601 4019 2635
rect 5641 2601 5675 2635
rect 7665 2601 7699 2635
rect 8309 2601 8343 2635
rect 14841 2601 14875 2635
rect 2237 2533 2271 2567
rect 4077 2533 4111 2567
rect 5825 2533 5859 2567
rect 10977 2533 11011 2567
rect 11897 2533 11931 2567
rect 11989 2533 12023 2567
rect 9597 2465 9631 2499
rect 2237 2397 2271 2431
rect 2513 2397 2547 2431
rect 3157 2397 3191 2431
rect 3433 2397 3467 2431
rect 3985 2397 4019 2431
rect 4261 2397 4295 2431
rect 7665 2397 7699 2431
rect 7849 2397 7883 2431
rect 8309 2397 8343 2431
rect 8585 2397 8619 2431
rect 9864 2397 9898 2431
rect 11897 2397 11931 2431
rect 15025 2397 15059 2431
rect 15301 2397 15335 2431
rect 5457 2329 5491 2363
rect 5673 2329 5707 2363
rect 8493 2329 8527 2363
rect 12173 2329 12207 2363
rect 2421 2261 2455 2295
rect 15209 2261 15243 2295
<< metal1 >>
rect 1104 19610 21043 19632
rect 1104 19558 5894 19610
rect 5946 19558 5958 19610
rect 6010 19558 6022 19610
rect 6074 19558 6086 19610
rect 6138 19558 6150 19610
rect 6202 19558 10839 19610
rect 10891 19558 10903 19610
rect 10955 19558 10967 19610
rect 11019 19558 11031 19610
rect 11083 19558 11095 19610
rect 11147 19558 15784 19610
rect 15836 19558 15848 19610
rect 15900 19558 15912 19610
rect 15964 19558 15976 19610
rect 16028 19558 16040 19610
rect 16092 19558 20729 19610
rect 20781 19558 20793 19610
rect 20845 19558 20857 19610
rect 20909 19558 20921 19610
rect 20973 19558 20985 19610
rect 21037 19558 21043 19610
rect 1104 19536 21043 19558
rect 1104 19066 20884 19088
rect 1104 19014 3422 19066
rect 3474 19014 3486 19066
rect 3538 19014 3550 19066
rect 3602 19014 3614 19066
rect 3666 19014 3678 19066
rect 3730 19014 8367 19066
rect 8419 19014 8431 19066
rect 8483 19014 8495 19066
rect 8547 19014 8559 19066
rect 8611 19014 8623 19066
rect 8675 19014 13312 19066
rect 13364 19014 13376 19066
rect 13428 19014 13440 19066
rect 13492 19014 13504 19066
rect 13556 19014 13568 19066
rect 13620 19014 18257 19066
rect 18309 19014 18321 19066
rect 18373 19014 18385 19066
rect 18437 19014 18449 19066
rect 18501 19014 18513 19066
rect 18565 19014 20884 19066
rect 1104 18992 20884 19014
rect 1581 18751 1639 18757
rect 1581 18717 1593 18751
rect 1627 18748 1639 18751
rect 2314 18748 2320 18760
rect 1627 18720 2320 18748
rect 1627 18717 1639 18720
rect 1581 18711 1639 18717
rect 2314 18708 2320 18720
rect 2372 18708 2378 18760
rect 1854 18680 1860 18692
rect 1815 18652 1860 18680
rect 1854 18640 1860 18652
rect 1912 18640 1918 18692
rect 1104 18522 21043 18544
rect 1104 18470 5894 18522
rect 5946 18470 5958 18522
rect 6010 18470 6022 18522
rect 6074 18470 6086 18522
rect 6138 18470 6150 18522
rect 6202 18470 10839 18522
rect 10891 18470 10903 18522
rect 10955 18470 10967 18522
rect 11019 18470 11031 18522
rect 11083 18470 11095 18522
rect 11147 18470 15784 18522
rect 15836 18470 15848 18522
rect 15900 18470 15912 18522
rect 15964 18470 15976 18522
rect 16028 18470 16040 18522
rect 16092 18470 20729 18522
rect 20781 18470 20793 18522
rect 20845 18470 20857 18522
rect 20909 18470 20921 18522
rect 20973 18470 20985 18522
rect 21037 18470 21043 18522
rect 1104 18448 21043 18470
rect 1104 17978 20884 18000
rect 1104 17926 3422 17978
rect 3474 17926 3486 17978
rect 3538 17926 3550 17978
rect 3602 17926 3614 17978
rect 3666 17926 3678 17978
rect 3730 17926 8367 17978
rect 8419 17926 8431 17978
rect 8483 17926 8495 17978
rect 8547 17926 8559 17978
rect 8611 17926 8623 17978
rect 8675 17926 13312 17978
rect 13364 17926 13376 17978
rect 13428 17926 13440 17978
rect 13492 17926 13504 17978
rect 13556 17926 13568 17978
rect 13620 17926 18257 17978
rect 18309 17926 18321 17978
rect 18373 17926 18385 17978
rect 18437 17926 18449 17978
rect 18501 17926 18513 17978
rect 18565 17926 20884 17978
rect 1104 17904 20884 17926
rect 1104 17434 21043 17456
rect 1104 17382 5894 17434
rect 5946 17382 5958 17434
rect 6010 17382 6022 17434
rect 6074 17382 6086 17434
rect 6138 17382 6150 17434
rect 6202 17382 10839 17434
rect 10891 17382 10903 17434
rect 10955 17382 10967 17434
rect 11019 17382 11031 17434
rect 11083 17382 11095 17434
rect 11147 17382 15784 17434
rect 15836 17382 15848 17434
rect 15900 17382 15912 17434
rect 15964 17382 15976 17434
rect 16028 17382 16040 17434
rect 16092 17382 20729 17434
rect 20781 17382 20793 17434
rect 20845 17382 20857 17434
rect 20909 17382 20921 17434
rect 20973 17382 20985 17434
rect 21037 17382 21043 17434
rect 1104 17360 21043 17382
rect 5626 17212 5632 17264
rect 5684 17252 5690 17264
rect 5684 17224 7972 17252
rect 5684 17212 5690 17224
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17153 4399 17187
rect 4341 17147 4399 17153
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17184 4491 17187
rect 5534 17184 5540 17196
rect 4479 17156 5540 17184
rect 4479 17153 4491 17156
rect 4433 17147 4491 17153
rect 4356 17048 4384 17147
rect 5534 17144 5540 17156
rect 5592 17184 5598 17196
rect 6748 17193 6776 17224
rect 7944 17196 7972 17224
rect 6549 17187 6607 17193
rect 6549 17184 6561 17187
rect 5592 17156 6561 17184
rect 5592 17144 5598 17156
rect 6549 17153 6561 17156
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 6733 17187 6791 17193
rect 6733 17153 6745 17187
rect 6779 17153 6791 17187
rect 7742 17184 7748 17196
rect 7703 17156 7748 17184
rect 6733 17147 6791 17153
rect 4617 17119 4675 17125
rect 4617 17085 4629 17119
rect 4663 17116 4675 17119
rect 5626 17116 5632 17128
rect 4663 17088 5632 17116
rect 4663 17085 4675 17088
rect 4617 17079 4675 17085
rect 5626 17076 5632 17088
rect 5684 17076 5690 17128
rect 6564 17116 6592 17147
rect 7742 17144 7748 17156
rect 7800 17144 7806 17196
rect 7926 17144 7932 17196
rect 7984 17184 7990 17196
rect 7984 17156 8077 17184
rect 7984 17144 7990 17156
rect 6822 17116 6828 17128
rect 6564 17088 6828 17116
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 4982 17048 4988 17060
rect 4356 17020 4988 17048
rect 4982 17008 4988 17020
rect 5040 17008 5046 17060
rect 4522 16940 4528 16992
rect 4580 16980 4586 16992
rect 4580 16952 4625 16980
rect 4580 16940 4586 16952
rect 6086 16940 6092 16992
rect 6144 16980 6150 16992
rect 6546 16980 6552 16992
rect 6144 16952 6552 16980
rect 6144 16940 6150 16952
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 7558 16940 7564 16992
rect 7616 16980 7622 16992
rect 7837 16983 7895 16989
rect 7837 16980 7849 16983
rect 7616 16952 7849 16980
rect 7616 16940 7622 16952
rect 7837 16949 7849 16952
rect 7883 16949 7895 16983
rect 7837 16943 7895 16949
rect 1104 16890 20884 16912
rect 1104 16838 3422 16890
rect 3474 16838 3486 16890
rect 3538 16838 3550 16890
rect 3602 16838 3614 16890
rect 3666 16838 3678 16890
rect 3730 16838 8367 16890
rect 8419 16838 8431 16890
rect 8483 16838 8495 16890
rect 8547 16838 8559 16890
rect 8611 16838 8623 16890
rect 8675 16838 13312 16890
rect 13364 16838 13376 16890
rect 13428 16838 13440 16890
rect 13492 16838 13504 16890
rect 13556 16838 13568 16890
rect 13620 16838 18257 16890
rect 18309 16838 18321 16890
rect 18373 16838 18385 16890
rect 18437 16838 18449 16890
rect 18501 16838 18513 16890
rect 18565 16838 20884 16890
rect 1104 16816 20884 16838
rect 5626 16776 5632 16788
rect 4816 16748 5632 16776
rect 4816 16708 4844 16748
rect 5626 16736 5632 16748
rect 5684 16736 5690 16788
rect 4632 16680 4844 16708
rect 4632 16649 4660 16680
rect 4982 16668 4988 16720
rect 5040 16708 5046 16720
rect 6914 16708 6920 16720
rect 5040 16680 6920 16708
rect 5040 16668 5046 16680
rect 4617 16643 4675 16649
rect 4617 16609 4629 16643
rect 4663 16609 4675 16643
rect 5534 16640 5540 16652
rect 4617 16603 4675 16609
rect 4816 16612 5540 16640
rect 3326 16572 3332 16584
rect 3287 16544 3332 16572
rect 3326 16532 3332 16544
rect 3384 16532 3390 16584
rect 3421 16575 3479 16581
rect 3421 16541 3433 16575
rect 3467 16572 3479 16575
rect 4522 16572 4528 16584
rect 3467 16544 4528 16572
rect 3467 16541 3479 16544
rect 3421 16535 3479 16541
rect 4522 16532 4528 16544
rect 4580 16532 4586 16584
rect 4816 16581 4844 16612
rect 5534 16600 5540 16612
rect 5592 16600 5598 16652
rect 6086 16640 6092 16652
rect 6047 16612 6092 16640
rect 6086 16600 6092 16612
rect 6144 16600 6150 16652
rect 6288 16649 6316 16680
rect 6914 16668 6920 16680
rect 6972 16708 6978 16720
rect 7009 16711 7067 16717
rect 7009 16708 7021 16711
rect 6972 16680 7021 16708
rect 6972 16668 6978 16680
rect 7009 16677 7021 16680
rect 7055 16677 7067 16711
rect 7009 16671 7067 16677
rect 6181 16643 6239 16649
rect 6181 16609 6193 16643
rect 6227 16609 6239 16643
rect 6181 16603 6239 16609
rect 6273 16643 6331 16649
rect 6273 16609 6285 16643
rect 6319 16609 6331 16643
rect 6273 16603 6331 16609
rect 6365 16643 6423 16649
rect 6365 16609 6377 16643
rect 6411 16640 6423 16643
rect 7745 16643 7803 16649
rect 7745 16640 7757 16643
rect 6411 16612 7757 16640
rect 6411 16609 6423 16612
rect 6365 16603 6423 16609
rect 7745 16609 7757 16612
rect 7791 16609 7803 16643
rect 15562 16640 15568 16652
rect 7745 16603 7803 16609
rect 14752 16612 15568 16640
rect 4801 16575 4859 16581
rect 4801 16541 4813 16575
rect 4847 16541 4859 16575
rect 4801 16535 4859 16541
rect 5718 16532 5724 16584
rect 5776 16572 5782 16584
rect 6196 16572 6224 16603
rect 7558 16572 7564 16584
rect 5776 16544 6224 16572
rect 7519 16544 7564 16572
rect 5776 16532 5782 16544
rect 7558 16532 7564 16544
rect 7616 16532 7622 16584
rect 7926 16532 7932 16584
rect 7984 16572 7990 16584
rect 8389 16575 8447 16581
rect 8389 16572 8401 16575
rect 7984 16544 8401 16572
rect 7984 16532 7990 16544
rect 8389 16541 8401 16544
rect 8435 16541 8447 16575
rect 8389 16535 8447 16541
rect 10965 16575 11023 16581
rect 10965 16541 10977 16575
rect 11011 16572 11023 16575
rect 11514 16572 11520 16584
rect 11011 16544 11520 16572
rect 11011 16541 11023 16544
rect 10965 16535 11023 16541
rect 11514 16532 11520 16544
rect 11572 16532 11578 16584
rect 14752 16581 14780 16612
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 14737 16575 14795 16581
rect 14737 16541 14749 16575
rect 14783 16541 14795 16575
rect 14737 16535 14795 16541
rect 14921 16575 14979 16581
rect 14921 16541 14933 16575
rect 14967 16541 14979 16575
rect 14921 16535 14979 16541
rect 3145 16507 3203 16513
rect 3145 16473 3157 16507
rect 3191 16504 3203 16507
rect 4706 16504 4712 16516
rect 3191 16476 4712 16504
rect 3191 16473 3203 16476
rect 3145 16467 3203 16473
rect 4706 16464 4712 16476
rect 4764 16504 4770 16516
rect 4764 16476 6316 16504
rect 4764 16464 4770 16476
rect 3234 16436 3240 16448
rect 3195 16408 3240 16436
rect 3234 16396 3240 16408
rect 3292 16396 3298 16448
rect 4985 16439 5043 16445
rect 4985 16405 4997 16439
rect 5031 16436 5043 16439
rect 5166 16436 5172 16448
rect 5031 16408 5172 16436
rect 5031 16405 5043 16408
rect 4985 16399 5043 16405
rect 5166 16396 5172 16408
rect 5224 16396 5230 16448
rect 5810 16396 5816 16448
rect 5868 16436 5874 16448
rect 5905 16439 5963 16445
rect 5905 16436 5917 16439
rect 5868 16408 5917 16436
rect 5868 16396 5874 16408
rect 5905 16405 5917 16408
rect 5951 16405 5963 16439
rect 6288 16436 6316 16476
rect 6822 16464 6828 16516
rect 6880 16504 6886 16516
rect 7009 16507 7067 16513
rect 7009 16504 7021 16507
rect 6880 16476 7021 16504
rect 6880 16464 6886 16476
rect 7009 16473 7021 16476
rect 7055 16473 7067 16507
rect 7009 16467 7067 16473
rect 7742 16464 7748 16516
rect 7800 16504 7806 16516
rect 8205 16507 8263 16513
rect 8205 16504 8217 16507
rect 7800 16476 8217 16504
rect 7800 16464 7806 16476
rect 8205 16473 8217 16476
rect 8251 16473 8263 16507
rect 8205 16467 8263 16473
rect 8573 16507 8631 16513
rect 8573 16473 8585 16507
rect 8619 16473 8631 16507
rect 8573 16467 8631 16473
rect 11241 16507 11299 16513
rect 11241 16473 11253 16507
rect 11287 16504 11299 16507
rect 11698 16504 11704 16516
rect 11287 16476 11704 16504
rect 11287 16473 11299 16476
rect 11241 16467 11299 16473
rect 7466 16436 7472 16448
rect 6288 16408 7472 16436
rect 5905 16399 5963 16405
rect 7466 16396 7472 16408
rect 7524 16436 7530 16448
rect 8588 16436 8616 16467
rect 11698 16464 11704 16476
rect 11756 16464 11762 16516
rect 14642 16464 14648 16516
rect 14700 16504 14706 16516
rect 14936 16504 14964 16535
rect 14700 16476 14964 16504
rect 14700 16464 14706 16476
rect 7524 16408 8616 16436
rect 14829 16439 14887 16445
rect 7524 16396 7530 16408
rect 14829 16405 14841 16439
rect 14875 16436 14887 16439
rect 15102 16436 15108 16448
rect 14875 16408 15108 16436
rect 14875 16405 14887 16408
rect 14829 16399 14887 16405
rect 15102 16396 15108 16408
rect 15160 16396 15166 16448
rect 1104 16346 21043 16368
rect 1104 16294 5894 16346
rect 5946 16294 5958 16346
rect 6010 16294 6022 16346
rect 6074 16294 6086 16346
rect 6138 16294 6150 16346
rect 6202 16294 10839 16346
rect 10891 16294 10903 16346
rect 10955 16294 10967 16346
rect 11019 16294 11031 16346
rect 11083 16294 11095 16346
rect 11147 16294 15784 16346
rect 15836 16294 15848 16346
rect 15900 16294 15912 16346
rect 15964 16294 15976 16346
rect 16028 16294 16040 16346
rect 16092 16294 20729 16346
rect 20781 16294 20793 16346
rect 20845 16294 20857 16346
rect 20909 16294 20921 16346
rect 20973 16294 20985 16346
rect 21037 16294 21043 16346
rect 1104 16272 21043 16294
rect 3326 16192 3332 16244
rect 3384 16232 3390 16244
rect 5718 16232 5724 16244
rect 3384 16204 5724 16232
rect 3384 16192 3390 16204
rect 3712 16136 4936 16164
rect 3712 16105 3740 16136
rect 3697 16099 3755 16105
rect 3697 16065 3709 16099
rect 3743 16065 3755 16099
rect 3697 16059 3755 16065
rect 4617 16099 4675 16105
rect 4617 16065 4629 16099
rect 4663 16065 4675 16099
rect 4617 16059 4675 16065
rect 3973 16031 4031 16037
rect 3973 15997 3985 16031
rect 4019 16028 4031 16031
rect 4433 16031 4491 16037
rect 4433 16028 4445 16031
rect 4019 16000 4445 16028
rect 4019 15997 4031 16000
rect 3973 15991 4031 15997
rect 4433 15997 4445 16000
rect 4479 15997 4491 16031
rect 4433 15991 4491 15997
rect 4632 15960 4660 16059
rect 4706 16056 4712 16108
rect 4764 16096 4770 16108
rect 4908 16105 4936 16136
rect 4893 16099 4951 16105
rect 4764 16068 4809 16096
rect 4764 16056 4770 16068
rect 4893 16065 4905 16099
rect 4939 16065 4951 16099
rect 4893 16059 4951 16065
rect 4908 16028 4936 16059
rect 4982 16056 4988 16108
rect 5040 16096 5046 16108
rect 5460 16105 5488 16204
rect 5718 16192 5724 16204
rect 5776 16192 5782 16244
rect 11698 16192 11704 16244
rect 11756 16232 11762 16244
rect 11756 16204 15700 16232
rect 11756 16192 11762 16204
rect 9677 16167 9735 16173
rect 9677 16133 9689 16167
rect 9723 16164 9735 16167
rect 12897 16167 12955 16173
rect 12897 16164 12909 16167
rect 9723 16136 12909 16164
rect 9723 16133 9735 16136
rect 9677 16127 9735 16133
rect 12897 16133 12909 16136
rect 12943 16133 12955 16167
rect 12897 16127 12955 16133
rect 5445 16099 5503 16105
rect 5040 16068 5085 16096
rect 5040 16056 5046 16068
rect 5445 16065 5457 16099
rect 5491 16065 5503 16099
rect 5626 16096 5632 16108
rect 5587 16068 5632 16096
rect 5445 16059 5503 16065
rect 5626 16056 5632 16068
rect 5684 16056 5690 16108
rect 6546 16096 6552 16108
rect 6507 16068 6552 16096
rect 6546 16056 6552 16068
rect 6604 16056 6610 16108
rect 7469 16099 7527 16105
rect 7469 16065 7481 16099
rect 7515 16065 7527 16099
rect 7469 16059 7527 16065
rect 5166 16028 5172 16040
rect 4908 16000 5172 16028
rect 5166 15988 5172 16000
rect 5224 16028 5230 16040
rect 6641 16031 6699 16037
rect 6641 16028 6653 16031
rect 5224 16000 6653 16028
rect 5224 15988 5230 16000
rect 6641 15997 6653 16000
rect 6687 15997 6699 16031
rect 6641 15991 6699 15997
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 6914 16028 6920 16040
rect 6871 16000 6920 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 6914 15988 6920 16000
rect 6972 16028 6978 16040
rect 7282 16028 7288 16040
rect 6972 16000 7288 16028
rect 6972 15988 6978 16000
rect 7282 15988 7288 16000
rect 7340 16028 7346 16040
rect 7484 16028 7512 16059
rect 7558 16056 7564 16108
rect 7616 16096 7622 16108
rect 7745 16099 7803 16105
rect 7745 16096 7757 16099
rect 7616 16068 7757 16096
rect 7616 16056 7622 16068
rect 7745 16065 7757 16068
rect 7791 16065 7803 16099
rect 9398 16096 9404 16108
rect 9359 16068 9404 16096
rect 7745 16059 7803 16065
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 9692 16068 10333 16096
rect 9692 16040 9720 16068
rect 10321 16065 10333 16068
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 11238 16056 11244 16108
rect 11296 16096 11302 16108
rect 12069 16099 12127 16105
rect 12069 16096 12081 16099
rect 11296 16068 12081 16096
rect 11296 16056 11302 16068
rect 12069 16065 12081 16068
rect 12115 16065 12127 16099
rect 13078 16096 13084 16108
rect 13039 16068 13084 16096
rect 12069 16059 12127 16065
rect 13078 16056 13084 16068
rect 13136 16056 13142 16108
rect 13173 16099 13231 16105
rect 13173 16065 13185 16099
rect 13219 16096 13231 16099
rect 13280 16096 13308 16204
rect 15194 16164 15200 16176
rect 13372 16136 15200 16164
rect 13372 16105 13400 16136
rect 15194 16124 15200 16136
rect 15252 16124 15258 16176
rect 15672 16108 15700 16204
rect 13219 16068 13308 16096
rect 13357 16099 13415 16105
rect 13219 16065 13231 16068
rect 13173 16059 13231 16065
rect 13357 16065 13369 16099
rect 13403 16065 13415 16099
rect 13357 16059 13415 16065
rect 13449 16099 13507 16105
rect 13449 16065 13461 16099
rect 13495 16096 13507 16099
rect 14366 16096 14372 16108
rect 13495 16068 14372 16096
rect 13495 16065 13507 16068
rect 13449 16059 13507 16065
rect 14366 16056 14372 16068
rect 14424 16056 14430 16108
rect 14550 16096 14556 16108
rect 14511 16068 14556 16096
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 14642 16056 14648 16108
rect 14700 16096 14706 16108
rect 14829 16099 14887 16105
rect 14700 16068 14793 16096
rect 14700 16056 14706 16068
rect 14829 16065 14841 16099
rect 14875 16065 14887 16099
rect 14829 16059 14887 16065
rect 7340 16000 7512 16028
rect 7340 15988 7346 16000
rect 7834 15988 7840 16040
rect 7892 16028 7898 16040
rect 9309 16031 9367 16037
rect 7892 16000 7937 16028
rect 7892 15988 7898 16000
rect 9309 15997 9321 16031
rect 9355 16028 9367 16031
rect 9674 16028 9680 16040
rect 9355 16000 9680 16028
rect 9355 15997 9367 16000
rect 9309 15991 9367 15997
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 9769 16031 9827 16037
rect 9769 15997 9781 16031
rect 9815 15997 9827 16031
rect 9769 15991 9827 15997
rect 5074 15960 5080 15972
rect 4632 15932 5080 15960
rect 5074 15920 5080 15932
rect 5132 15960 5138 15972
rect 5537 15963 5595 15969
rect 5537 15960 5549 15963
rect 5132 15932 5549 15960
rect 5132 15920 5138 15932
rect 5537 15929 5549 15932
rect 5583 15929 5595 15963
rect 5537 15923 5595 15929
rect 7466 15920 7472 15972
rect 7524 15960 7530 15972
rect 7561 15963 7619 15969
rect 7561 15960 7573 15963
rect 7524 15932 7573 15960
rect 7524 15920 7530 15932
rect 7561 15929 7573 15932
rect 7607 15929 7619 15963
rect 7561 15923 7619 15929
rect 9214 15920 9220 15972
rect 9272 15960 9278 15972
rect 9784 15960 9812 15991
rect 11790 15988 11796 16040
rect 11848 16028 11854 16040
rect 12161 16031 12219 16037
rect 12161 16028 12173 16031
rect 11848 16000 12173 16028
rect 11848 15988 11854 16000
rect 12161 15997 12173 16000
rect 12207 15997 12219 16031
rect 12161 15991 12219 15997
rect 12253 16031 12311 16037
rect 12253 15997 12265 16031
rect 12299 15997 12311 16031
rect 14660 16028 14688 16056
rect 12253 15991 12311 15997
rect 13188 16000 14688 16028
rect 9272 15932 9812 15960
rect 9272 15920 9278 15932
rect 11330 15920 11336 15972
rect 11388 15960 11394 15972
rect 12268 15960 12296 15991
rect 13188 15972 13216 16000
rect 14734 15988 14740 16040
rect 14792 16028 14798 16040
rect 14844 16028 14872 16059
rect 14918 16056 14924 16108
rect 14976 16096 14982 16108
rect 15102 16105 15108 16108
rect 15059 16099 15108 16105
rect 14976 16068 15021 16096
rect 14976 16056 14982 16068
rect 15059 16065 15071 16099
rect 15105 16065 15108 16099
rect 15059 16059 15108 16065
rect 15102 16056 15108 16059
rect 15160 16056 15166 16108
rect 15654 16056 15660 16108
rect 15712 16096 15718 16108
rect 16025 16099 16083 16105
rect 16025 16096 16037 16099
rect 15712 16068 16037 16096
rect 15712 16056 15718 16068
rect 16025 16065 16037 16068
rect 16071 16065 16083 16099
rect 16025 16059 16083 16065
rect 14792 16000 14872 16028
rect 15841 16031 15899 16037
rect 14792 15988 14798 16000
rect 15841 15997 15853 16031
rect 15887 15997 15899 16031
rect 15841 15991 15899 15997
rect 11388 15932 12296 15960
rect 11388 15920 11394 15932
rect 3786 15892 3792 15904
rect 3747 15864 3792 15892
rect 3786 15852 3792 15864
rect 3844 15852 3850 15904
rect 3881 15895 3939 15901
rect 3881 15861 3893 15895
rect 3927 15892 3939 15895
rect 4706 15892 4712 15904
rect 3927 15864 4712 15892
rect 3927 15861 3939 15864
rect 3881 15855 3939 15861
rect 4706 15852 4712 15864
rect 4764 15852 4770 15904
rect 6733 15895 6791 15901
rect 6733 15861 6745 15895
rect 6779 15892 6791 15895
rect 6914 15892 6920 15904
rect 6779 15864 6920 15892
rect 6779 15861 6791 15864
rect 6733 15855 6791 15861
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 7650 15852 7656 15904
rect 7708 15892 7714 15904
rect 7708 15864 7753 15892
rect 7708 15852 7714 15864
rect 8846 15852 8852 15904
rect 8904 15892 8910 15904
rect 9125 15895 9183 15901
rect 9125 15892 9137 15895
rect 8904 15864 9137 15892
rect 8904 15852 8910 15864
rect 9125 15861 9137 15864
rect 9171 15861 9183 15895
rect 9125 15855 9183 15861
rect 10410 15852 10416 15904
rect 10468 15892 10474 15904
rect 10505 15895 10563 15901
rect 10505 15892 10517 15895
rect 10468 15864 10517 15892
rect 10468 15852 10474 15864
rect 10505 15861 10517 15864
rect 10551 15861 10563 15895
rect 10505 15855 10563 15861
rect 10870 15852 10876 15904
rect 10928 15892 10934 15904
rect 11701 15895 11759 15901
rect 11701 15892 11713 15895
rect 10928 15864 11713 15892
rect 10928 15852 10934 15864
rect 11701 15861 11713 15864
rect 11747 15861 11759 15895
rect 12268 15892 12296 15932
rect 13170 15920 13176 15972
rect 13228 15920 13234 15972
rect 14182 15920 14188 15972
rect 14240 15960 14246 15972
rect 14550 15960 14556 15972
rect 14240 15932 14556 15960
rect 14240 15920 14246 15932
rect 14550 15920 14556 15932
rect 14608 15920 14614 15972
rect 15197 15963 15255 15969
rect 15197 15929 15209 15963
rect 15243 15960 15255 15963
rect 15856 15960 15884 15991
rect 15930 15988 15936 16040
rect 15988 16028 15994 16040
rect 16117 16031 16175 16037
rect 15988 16000 16033 16028
rect 15988 15988 15994 16000
rect 16117 15997 16129 16031
rect 16163 16028 16175 16031
rect 17034 16028 17040 16040
rect 16163 16000 17040 16028
rect 16163 15997 16175 16000
rect 16117 15991 16175 15997
rect 17034 15988 17040 16000
rect 17092 15988 17098 16040
rect 15243 15932 15884 15960
rect 15243 15929 15255 15932
rect 15197 15923 15255 15929
rect 14642 15892 14648 15904
rect 12268 15864 14648 15892
rect 11701 15855 11759 15861
rect 14642 15852 14648 15864
rect 14700 15852 14706 15904
rect 15657 15895 15715 15901
rect 15657 15861 15669 15895
rect 15703 15892 15715 15895
rect 16114 15892 16120 15904
rect 15703 15864 16120 15892
rect 15703 15861 15715 15864
rect 15657 15855 15715 15861
rect 16114 15852 16120 15864
rect 16172 15852 16178 15904
rect 1104 15802 20884 15824
rect 1104 15750 3422 15802
rect 3474 15750 3486 15802
rect 3538 15750 3550 15802
rect 3602 15750 3614 15802
rect 3666 15750 3678 15802
rect 3730 15750 8367 15802
rect 8419 15750 8431 15802
rect 8483 15750 8495 15802
rect 8547 15750 8559 15802
rect 8611 15750 8623 15802
rect 8675 15750 13312 15802
rect 13364 15750 13376 15802
rect 13428 15750 13440 15802
rect 13492 15750 13504 15802
rect 13556 15750 13568 15802
rect 13620 15750 18257 15802
rect 18309 15750 18321 15802
rect 18373 15750 18385 15802
rect 18437 15750 18449 15802
rect 18501 15750 18513 15802
rect 18565 15750 20884 15802
rect 1104 15728 20884 15750
rect 9214 15688 9220 15700
rect 9175 15660 9220 15688
rect 9214 15648 9220 15660
rect 9272 15648 9278 15700
rect 9398 15648 9404 15700
rect 9456 15688 9462 15700
rect 10413 15691 10471 15697
rect 10413 15688 10425 15691
rect 9456 15660 10425 15688
rect 9456 15648 9462 15660
rect 10413 15657 10425 15660
rect 10459 15657 10471 15691
rect 10870 15688 10876 15700
rect 10831 15660 10876 15688
rect 10413 15651 10471 15657
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 12526 15648 12532 15700
rect 12584 15688 12590 15700
rect 14553 15691 14611 15697
rect 12584 15660 14504 15688
rect 12584 15648 12590 15660
rect 6822 15580 6828 15632
rect 6880 15620 6886 15632
rect 7745 15623 7803 15629
rect 7745 15620 7757 15623
rect 6880 15592 7757 15620
rect 6880 15580 6886 15592
rect 7745 15589 7757 15592
rect 7791 15589 7803 15623
rect 9858 15620 9864 15632
rect 7745 15583 7803 15589
rect 9508 15592 9864 15620
rect 2593 15555 2651 15561
rect 2593 15521 2605 15555
rect 2639 15552 2651 15555
rect 3142 15552 3148 15564
rect 2639 15524 3148 15552
rect 2639 15521 2651 15524
rect 2593 15515 2651 15521
rect 3142 15512 3148 15524
rect 3200 15512 3206 15564
rect 2409 15487 2467 15493
rect 2409 15453 2421 15487
rect 2455 15484 2467 15487
rect 3234 15484 3240 15496
rect 2455 15456 3240 15484
rect 2455 15453 2467 15456
rect 2409 15447 2467 15453
rect 3234 15444 3240 15456
rect 3292 15444 3298 15496
rect 7561 15487 7619 15493
rect 7561 15453 7573 15487
rect 7607 15453 7619 15487
rect 7742 15484 7748 15496
rect 7703 15456 7748 15484
rect 7561 15447 7619 15453
rect 7576 15416 7604 15447
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 9508 15493 9536 15592
rect 9858 15580 9864 15592
rect 9916 15580 9922 15632
rect 12621 15623 12679 15629
rect 12621 15589 12633 15623
rect 12667 15620 12679 15623
rect 13078 15620 13084 15632
rect 12667 15592 13084 15620
rect 12667 15589 12679 15592
rect 12621 15583 12679 15589
rect 13078 15580 13084 15592
rect 13136 15620 13142 15632
rect 13354 15620 13360 15632
rect 13136 15592 13360 15620
rect 13136 15580 13142 15592
rect 13354 15580 13360 15592
rect 13412 15580 13418 15632
rect 14476 15620 14504 15660
rect 14553 15657 14565 15691
rect 14599 15688 14611 15691
rect 14734 15688 14740 15700
rect 14599 15660 14740 15688
rect 14599 15657 14611 15660
rect 14553 15651 14611 15657
rect 14734 15648 14740 15660
rect 14792 15648 14798 15700
rect 15930 15648 15936 15700
rect 15988 15688 15994 15700
rect 16025 15691 16083 15697
rect 16025 15688 16037 15691
rect 15988 15660 16037 15688
rect 15988 15648 15994 15660
rect 16025 15657 16037 15660
rect 16071 15657 16083 15691
rect 17034 15688 17040 15700
rect 16995 15660 17040 15688
rect 16025 15651 16083 15657
rect 17034 15648 17040 15660
rect 17092 15648 17098 15700
rect 14918 15620 14924 15632
rect 14476 15592 14924 15620
rect 14918 15580 14924 15592
rect 14976 15580 14982 15632
rect 15286 15580 15292 15632
rect 15344 15620 15350 15632
rect 15344 15592 17724 15620
rect 15344 15580 15350 15592
rect 12805 15555 12863 15561
rect 12805 15552 12817 15555
rect 12268 15524 12817 15552
rect 9493 15487 9551 15493
rect 9493 15453 9505 15487
rect 9539 15453 9551 15487
rect 9493 15447 9551 15453
rect 10597 15487 10655 15493
rect 10597 15453 10609 15487
rect 10643 15453 10655 15487
rect 10597 15447 10655 15453
rect 8018 15416 8024 15428
rect 7576 15388 8024 15416
rect 8018 15376 8024 15388
rect 8076 15376 8082 15428
rect 9217 15419 9275 15425
rect 9217 15385 9229 15419
rect 9263 15416 9275 15419
rect 10410 15416 10416 15428
rect 9263 15388 10416 15416
rect 9263 15385 9275 15388
rect 9217 15379 9275 15385
rect 10410 15376 10416 15388
rect 10468 15376 10474 15428
rect 10612 15416 10640 15447
rect 10686 15444 10692 15496
rect 10744 15484 10750 15496
rect 10965 15487 11023 15493
rect 10744 15456 10789 15484
rect 10744 15444 10750 15456
rect 10965 15453 10977 15487
rect 11011 15484 11023 15487
rect 11054 15484 11060 15496
rect 11011 15456 11060 15484
rect 11011 15453 11023 15456
rect 10965 15447 11023 15453
rect 11054 15444 11060 15456
rect 11112 15444 11118 15496
rect 11422 15484 11428 15496
rect 11383 15456 11428 15484
rect 11422 15444 11428 15456
rect 11480 15444 11486 15496
rect 11514 15444 11520 15496
rect 11572 15484 11578 15496
rect 12268 15484 12296 15524
rect 12805 15521 12817 15524
rect 12851 15552 12863 15555
rect 13814 15552 13820 15564
rect 12851 15524 13820 15552
rect 12851 15521 12863 15524
rect 12805 15515 12863 15521
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 16666 15552 16672 15564
rect 14660 15524 16672 15552
rect 14660 15496 14688 15524
rect 11572 15456 12296 15484
rect 11572 15444 11578 15456
rect 12526 15444 12532 15496
rect 12584 15484 12590 15496
rect 12584 15456 12629 15484
rect 12584 15444 12590 15456
rect 13170 15444 13176 15496
rect 13228 15484 13234 15496
rect 13265 15487 13323 15493
rect 13265 15484 13277 15487
rect 13228 15456 13277 15484
rect 13228 15444 13234 15456
rect 13265 15453 13277 15456
rect 13311 15453 13323 15487
rect 13265 15447 13323 15453
rect 13449 15487 13507 15493
rect 13449 15453 13461 15487
rect 13495 15484 13507 15487
rect 13630 15484 13636 15496
rect 13495 15456 13636 15484
rect 13495 15453 13507 15456
rect 13449 15447 13507 15453
rect 13630 15444 13636 15456
rect 13688 15444 13694 15496
rect 14458 15484 14464 15496
rect 14419 15456 14464 15484
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 14642 15484 14648 15496
rect 14603 15456 14648 15484
rect 14642 15444 14648 15456
rect 14700 15444 14706 15496
rect 16316 15493 16344 15524
rect 16666 15512 16672 15524
rect 16724 15512 16730 15564
rect 16209 15487 16267 15493
rect 16209 15453 16221 15487
rect 16255 15453 16267 15487
rect 16209 15447 16267 15453
rect 16301 15487 16359 15493
rect 16301 15453 16313 15487
rect 16347 15453 16359 15487
rect 16482 15484 16488 15496
rect 16443 15456 16488 15484
rect 16301 15447 16359 15453
rect 12805 15419 12863 15425
rect 12805 15416 12817 15419
rect 10612 15388 12817 15416
rect 12805 15385 12817 15388
rect 12851 15385 12863 15419
rect 16224 15416 16252 15447
rect 16482 15444 16488 15456
rect 16540 15444 16546 15496
rect 16577 15487 16635 15493
rect 16577 15453 16589 15487
rect 16623 15484 16635 15487
rect 17313 15487 17371 15493
rect 17313 15484 17325 15487
rect 16623 15456 17325 15484
rect 16623 15453 16635 15456
rect 16577 15447 16635 15453
rect 16942 15416 16948 15428
rect 16224 15388 16948 15416
rect 12805 15379 12863 15385
rect 16942 15376 16948 15388
rect 17000 15376 17006 15428
rect 1946 15348 1952 15360
rect 1907 15320 1952 15348
rect 1946 15308 1952 15320
rect 2004 15308 2010 15360
rect 2222 15308 2228 15360
rect 2280 15348 2286 15360
rect 2317 15351 2375 15357
rect 2317 15348 2329 15351
rect 2280 15320 2329 15348
rect 2280 15308 2286 15320
rect 2317 15317 2329 15320
rect 2363 15317 2375 15351
rect 2317 15311 2375 15317
rect 9401 15351 9459 15357
rect 9401 15317 9413 15351
rect 9447 15348 9459 15351
rect 9766 15348 9772 15360
rect 9447 15320 9772 15348
rect 9447 15317 9459 15320
rect 9401 15311 9459 15317
rect 9766 15308 9772 15320
rect 9824 15348 9830 15360
rect 11054 15348 11060 15360
rect 9824 15320 11060 15348
rect 9824 15308 9830 15320
rect 11054 15308 11060 15320
rect 11112 15348 11118 15360
rect 11698 15348 11704 15360
rect 11112 15320 11704 15348
rect 11112 15308 11118 15320
rect 11698 15308 11704 15320
rect 11756 15308 11762 15360
rect 15470 15308 15476 15360
rect 15528 15348 15534 15360
rect 17052 15348 17080 15456
rect 17313 15453 17325 15456
rect 17359 15453 17371 15487
rect 17313 15447 17371 15453
rect 17405 15487 17463 15493
rect 17405 15453 17417 15487
rect 17451 15453 17463 15487
rect 17405 15447 17463 15453
rect 17420 15416 17448 15447
rect 17494 15444 17500 15496
rect 17552 15484 17558 15496
rect 17696 15493 17724 15592
rect 17681 15487 17739 15493
rect 17552 15456 17597 15484
rect 17552 15444 17558 15456
rect 17681 15453 17693 15487
rect 17727 15453 17739 15487
rect 17681 15447 17739 15453
rect 18414 15416 18420 15428
rect 17420 15388 18420 15416
rect 18414 15376 18420 15388
rect 18472 15376 18478 15428
rect 15528 15320 17080 15348
rect 15528 15308 15534 15320
rect 1104 15258 21043 15280
rect 1104 15206 5894 15258
rect 5946 15206 5958 15258
rect 6010 15206 6022 15258
rect 6074 15206 6086 15258
rect 6138 15206 6150 15258
rect 6202 15206 10839 15258
rect 10891 15206 10903 15258
rect 10955 15206 10967 15258
rect 11019 15206 11031 15258
rect 11083 15206 11095 15258
rect 11147 15206 15784 15258
rect 15836 15206 15848 15258
rect 15900 15206 15912 15258
rect 15964 15206 15976 15258
rect 16028 15206 16040 15258
rect 16092 15206 20729 15258
rect 20781 15206 20793 15258
rect 20845 15206 20857 15258
rect 20909 15206 20921 15258
rect 20973 15206 20985 15258
rect 21037 15206 21043 15258
rect 1104 15184 21043 15206
rect 7834 15104 7840 15156
rect 7892 15144 7898 15156
rect 8205 15147 8263 15153
rect 8205 15144 8217 15147
rect 7892 15116 8217 15144
rect 7892 15104 7898 15116
rect 8205 15113 8217 15116
rect 8251 15113 8263 15147
rect 8205 15107 8263 15113
rect 9674 15104 9680 15156
rect 9732 15144 9738 15156
rect 14274 15144 14280 15156
rect 9732 15116 14280 15144
rect 9732 15104 9738 15116
rect 5718 15036 5724 15088
rect 5776 15076 5782 15088
rect 7101 15079 7159 15085
rect 7101 15076 7113 15079
rect 5776 15048 7113 15076
rect 5776 15036 5782 15048
rect 7101 15045 7113 15048
rect 7147 15045 7159 15079
rect 7282 15076 7288 15088
rect 7243 15048 7288 15076
rect 7101 15039 7159 15045
rect 7282 15036 7288 15048
rect 7340 15036 7346 15088
rect 11422 15036 11428 15088
rect 11480 15076 11486 15088
rect 11480 15048 12020 15076
rect 11480 15036 11486 15048
rect 11992 15020 12020 15048
rect 2038 14968 2044 15020
rect 2096 15008 2102 15020
rect 2317 15011 2375 15017
rect 2317 15008 2329 15011
rect 2096 14980 2329 15008
rect 2096 14968 2102 14980
rect 2317 14977 2329 14980
rect 2363 14977 2375 15011
rect 2317 14971 2375 14977
rect 2501 15011 2559 15017
rect 2501 14977 2513 15011
rect 2547 14977 2559 15011
rect 7926 15008 7932 15020
rect 7887 14980 7932 15008
rect 2501 14971 2559 14977
rect 2222 14900 2228 14952
rect 2280 14940 2286 14952
rect 2516 14940 2544 14971
rect 7926 14968 7932 14980
rect 7984 14968 7990 15020
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 14977 11943 15011
rect 11885 14971 11943 14977
rect 2280 14912 2544 14940
rect 2280 14900 2286 14912
rect 8018 14900 8024 14952
rect 8076 14940 8082 14952
rect 8205 14943 8263 14949
rect 8205 14940 8217 14943
rect 8076 14912 8217 14940
rect 8076 14900 8082 14912
rect 8205 14909 8217 14912
rect 8251 14909 8263 14943
rect 8205 14903 8263 14909
rect 3878 14832 3884 14884
rect 3936 14872 3942 14884
rect 7098 14872 7104 14884
rect 3936 14844 7104 14872
rect 3936 14832 3942 14844
rect 7098 14832 7104 14844
rect 7156 14832 7162 14884
rect 7282 14832 7288 14884
rect 7340 14872 7346 14884
rect 11900 14872 11928 14971
rect 11974 14968 11980 15020
rect 12032 15008 12038 15020
rect 12158 15008 12164 15020
rect 12032 14980 12077 15008
rect 12119 14980 12164 15008
rect 12032 14968 12038 14980
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 12268 15017 12296 15116
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 14458 15104 14464 15156
rect 14516 15144 14522 15156
rect 14645 15147 14703 15153
rect 14645 15144 14657 15147
rect 14516 15116 14657 15144
rect 14516 15104 14522 15116
rect 14645 15113 14657 15116
rect 14691 15113 14703 15147
rect 16206 15144 16212 15156
rect 16119 15116 16212 15144
rect 14645 15107 14703 15113
rect 16206 15104 16212 15116
rect 16264 15144 16270 15156
rect 16482 15144 16488 15156
rect 16264 15116 16488 15144
rect 16264 15104 16270 15116
rect 16482 15104 16488 15116
rect 16540 15104 16546 15156
rect 17494 15144 17500 15156
rect 17455 15116 17500 15144
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 18141 15147 18199 15153
rect 18141 15113 18153 15147
rect 18187 15144 18199 15147
rect 19978 15144 19984 15156
rect 18187 15116 19984 15144
rect 18187 15113 18199 15116
rect 18141 15107 18199 15113
rect 19978 15104 19984 15116
rect 20036 15104 20042 15156
rect 13265 15079 13323 15085
rect 13265 15045 13277 15079
rect 13311 15076 13323 15079
rect 15841 15079 15899 15085
rect 15841 15076 15853 15079
rect 13311 15048 15853 15076
rect 13311 15045 13323 15048
rect 13265 15039 13323 15045
rect 15841 15045 15853 15048
rect 15887 15045 15899 15079
rect 15841 15039 15899 15045
rect 16057 15079 16115 15085
rect 16057 15045 16069 15079
rect 16103 15076 16115 15079
rect 16666 15076 16672 15088
rect 16103 15048 16672 15076
rect 16103 15045 16115 15048
rect 16057 15039 16115 15045
rect 12253 15011 12311 15017
rect 12253 14977 12265 15011
rect 12299 14977 12311 15011
rect 12253 14971 12311 14977
rect 13173 15011 13231 15017
rect 13173 14977 13185 15011
rect 13219 15008 13231 15011
rect 13722 15008 13728 15020
rect 13219 14980 13728 15008
rect 13219 14977 13231 14980
rect 13173 14971 13231 14977
rect 13722 14968 13728 14980
rect 13780 15008 13786 15020
rect 13780 14980 14504 15008
rect 13780 14968 13786 14980
rect 13354 14940 13360 14952
rect 13315 14912 13360 14940
rect 13354 14900 13360 14912
rect 13412 14900 13418 14952
rect 14476 14940 14504 14980
rect 14550 14968 14556 15020
rect 14608 15008 14614 15020
rect 14737 15011 14795 15017
rect 14608 14980 14653 15008
rect 14608 14968 14614 14980
rect 14737 14977 14749 15011
rect 14783 15008 14795 15011
rect 15010 15008 15016 15020
rect 14783 14980 15016 15008
rect 14783 14977 14795 14980
rect 14737 14971 14795 14977
rect 15010 14968 15016 14980
rect 15068 14968 15074 15020
rect 15856 15008 15884 15039
rect 16666 15036 16672 15048
rect 16724 15036 16730 15088
rect 17862 15036 17868 15088
rect 17920 15076 17926 15088
rect 18877 15079 18935 15085
rect 18877 15076 18889 15079
rect 17920 15048 18889 15076
rect 17920 15036 17926 15048
rect 18877 15045 18889 15048
rect 18923 15045 18935 15079
rect 18877 15039 18935 15045
rect 16390 15008 16396 15020
rect 15856 14980 16396 15008
rect 16390 14968 16396 14980
rect 16448 14968 16454 15020
rect 18233 15011 18291 15017
rect 18233 14977 18245 15011
rect 18279 14977 18291 15011
rect 18690 15008 18696 15020
rect 18651 14980 18696 15008
rect 18233 14971 18291 14977
rect 17773 14943 17831 14949
rect 17773 14940 17785 14943
rect 14476 14912 17785 14940
rect 17773 14909 17785 14912
rect 17819 14909 17831 14943
rect 17773 14903 17831 14909
rect 12805 14875 12863 14881
rect 12805 14872 12817 14875
rect 7340 14844 8064 14872
rect 11900 14844 12817 14872
rect 7340 14832 7346 14844
rect 2409 14807 2467 14813
rect 2409 14773 2421 14807
rect 2455 14804 2467 14807
rect 3142 14804 3148 14816
rect 2455 14776 3148 14804
rect 2455 14773 2467 14776
rect 2409 14767 2467 14773
rect 3142 14764 3148 14776
rect 3200 14764 3206 14816
rect 6822 14764 6828 14816
rect 6880 14804 6886 14816
rect 8036 14813 8064 14844
rect 12805 14841 12817 14844
rect 12851 14841 12863 14875
rect 12805 14835 12863 14841
rect 17126 14832 17132 14884
rect 17184 14872 17190 14884
rect 18248 14872 18276 14971
rect 18690 14968 18696 14980
rect 18748 14968 18754 15020
rect 18966 15008 18972 15020
rect 18927 14980 18972 15008
rect 18966 14968 18972 14980
rect 19024 14968 19030 15020
rect 17184 14844 18276 14872
rect 17184 14832 17190 14844
rect 18414 14832 18420 14884
rect 18472 14872 18478 14884
rect 18693 14875 18751 14881
rect 18693 14872 18705 14875
rect 18472 14844 18705 14872
rect 18472 14832 18478 14844
rect 18693 14841 18705 14844
rect 18739 14841 18751 14875
rect 18693 14835 18751 14841
rect 7469 14807 7527 14813
rect 7469 14804 7481 14807
rect 6880 14776 7481 14804
rect 6880 14764 6886 14776
rect 7469 14773 7481 14776
rect 7515 14773 7527 14807
rect 7469 14767 7527 14773
rect 8021 14807 8079 14813
rect 8021 14773 8033 14807
rect 8067 14804 8079 14807
rect 8202 14804 8208 14816
rect 8067 14776 8208 14804
rect 8067 14773 8079 14776
rect 8021 14767 8079 14773
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 11701 14807 11759 14813
rect 11701 14804 11713 14807
rect 10652 14776 11713 14804
rect 10652 14764 10658 14776
rect 11701 14773 11713 14776
rect 11747 14773 11759 14807
rect 11701 14767 11759 14773
rect 11790 14764 11796 14816
rect 11848 14804 11854 14816
rect 13078 14804 13084 14816
rect 11848 14776 13084 14804
rect 11848 14764 11854 14776
rect 13078 14764 13084 14776
rect 13136 14764 13142 14816
rect 14090 14764 14096 14816
rect 14148 14804 14154 14816
rect 16025 14807 16083 14813
rect 16025 14804 16037 14807
rect 14148 14776 16037 14804
rect 14148 14764 14154 14776
rect 16025 14773 16037 14776
rect 16071 14773 16083 14807
rect 17862 14804 17868 14816
rect 17823 14776 17868 14804
rect 16025 14767 16083 14773
rect 17862 14764 17868 14776
rect 17920 14764 17926 14816
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 18012 14776 18057 14804
rect 18012 14764 18018 14776
rect 1104 14714 20884 14736
rect 1104 14662 3422 14714
rect 3474 14662 3486 14714
rect 3538 14662 3550 14714
rect 3602 14662 3614 14714
rect 3666 14662 3678 14714
rect 3730 14662 8367 14714
rect 8419 14662 8431 14714
rect 8483 14662 8495 14714
rect 8547 14662 8559 14714
rect 8611 14662 8623 14714
rect 8675 14662 13312 14714
rect 13364 14662 13376 14714
rect 13428 14662 13440 14714
rect 13492 14662 13504 14714
rect 13556 14662 13568 14714
rect 13620 14662 18257 14714
rect 18309 14662 18321 14714
rect 18373 14662 18385 14714
rect 18437 14662 18449 14714
rect 18501 14662 18513 14714
rect 18565 14662 20884 14714
rect 1104 14640 20884 14662
rect 3050 14560 3056 14612
rect 3108 14600 3114 14612
rect 3786 14600 3792 14612
rect 3108 14572 3792 14600
rect 3108 14560 3114 14572
rect 3786 14560 3792 14572
rect 3844 14600 3850 14612
rect 7561 14603 7619 14609
rect 7561 14600 7573 14603
rect 3844 14572 7573 14600
rect 3844 14560 3850 14572
rect 7561 14569 7573 14572
rect 7607 14569 7619 14603
rect 8202 14600 8208 14612
rect 8163 14572 8208 14600
rect 7561 14563 7619 14569
rect 8202 14560 8208 14572
rect 8260 14560 8266 14612
rect 10686 14560 10692 14612
rect 10744 14600 10750 14612
rect 10744 14572 12112 14600
rect 10744 14560 10750 14572
rect 4154 14492 4160 14544
rect 4212 14532 4218 14544
rect 4982 14532 4988 14544
rect 4212 14504 4988 14532
rect 4212 14492 4218 14504
rect 4982 14492 4988 14504
rect 5040 14492 5046 14544
rect 9125 14535 9183 14541
rect 9125 14501 9137 14535
rect 9171 14532 9183 14535
rect 9490 14532 9496 14544
rect 9171 14504 9496 14532
rect 9171 14501 9183 14504
rect 9125 14495 9183 14501
rect 9490 14492 9496 14504
rect 9548 14492 9554 14544
rect 11238 14532 11244 14544
rect 10612 14504 11244 14532
rect 4525 14467 4583 14473
rect 4525 14464 4537 14467
rect 2976 14436 4537 14464
rect 2976 14405 3004 14436
rect 4525 14433 4537 14436
rect 4571 14433 4583 14467
rect 5000 14464 5028 14492
rect 5000 14436 5212 14464
rect 4525 14427 4583 14433
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14365 3019 14399
rect 2961 14359 3019 14365
rect 3050 14356 3056 14408
rect 3108 14396 3114 14408
rect 3326 14396 3332 14408
rect 3108 14368 3153 14396
rect 3287 14368 3332 14396
rect 3108 14356 3114 14368
rect 3326 14356 3332 14368
rect 3384 14356 3390 14408
rect 3418 14356 3424 14408
rect 3476 14396 3482 14408
rect 3878 14396 3884 14408
rect 3476 14368 3884 14396
rect 3476 14356 3482 14368
rect 3878 14356 3884 14368
rect 3936 14356 3942 14408
rect 4154 14396 4160 14408
rect 4115 14368 4160 14396
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 4249 14399 4307 14405
rect 4249 14365 4261 14399
rect 4295 14365 4307 14399
rect 4249 14359 4307 14365
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14365 4399 14399
rect 4341 14359 4399 14365
rect 4985 14399 5043 14405
rect 4985 14365 4997 14399
rect 5031 14396 5043 14399
rect 5074 14396 5080 14408
rect 5031 14368 5080 14396
rect 5031 14365 5043 14368
rect 4985 14359 5043 14365
rect 1949 14331 2007 14337
rect 1949 14297 1961 14331
rect 1995 14328 2007 14331
rect 2038 14328 2044 14340
rect 1995 14300 2044 14328
rect 1995 14297 2007 14300
rect 1949 14291 2007 14297
rect 2038 14288 2044 14300
rect 2096 14288 2102 14340
rect 2133 14331 2191 14337
rect 2133 14297 2145 14331
rect 2179 14328 2191 14331
rect 2222 14328 2228 14340
rect 2179 14300 2228 14328
rect 2179 14297 2191 14300
rect 2133 14291 2191 14297
rect 2222 14288 2228 14300
rect 2280 14288 2286 14340
rect 3145 14331 3203 14337
rect 3145 14297 3157 14331
rect 3191 14328 3203 14331
rect 3234 14328 3240 14340
rect 3191 14300 3240 14328
rect 3191 14297 3203 14300
rect 3145 14291 3203 14297
rect 3234 14288 3240 14300
rect 3292 14288 3298 14340
rect 2317 14263 2375 14269
rect 2317 14229 2329 14263
rect 2363 14260 2375 14263
rect 2406 14260 2412 14272
rect 2363 14232 2412 14260
rect 2363 14229 2375 14232
rect 2317 14223 2375 14229
rect 2406 14220 2412 14232
rect 2464 14220 2470 14272
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 4264 14260 4292 14359
rect 4356 14328 4384 14359
rect 5074 14356 5080 14368
rect 5132 14356 5138 14408
rect 5184 14396 5212 14436
rect 5258 14424 5264 14476
rect 5316 14464 5322 14476
rect 6089 14467 6147 14473
rect 6089 14464 6101 14467
rect 5316 14436 6101 14464
rect 5316 14424 5322 14436
rect 6089 14433 6101 14436
rect 6135 14433 6147 14467
rect 6089 14427 6147 14433
rect 7285 14467 7343 14473
rect 7285 14433 7297 14467
rect 7331 14464 7343 14467
rect 7558 14464 7564 14476
rect 7331 14436 7564 14464
rect 7331 14433 7343 14436
rect 7285 14427 7343 14433
rect 7558 14424 7564 14436
rect 7616 14464 7622 14476
rect 7926 14464 7932 14476
rect 7616 14436 7932 14464
rect 7616 14424 7622 14436
rect 7926 14424 7932 14436
rect 7984 14424 7990 14476
rect 9769 14467 9827 14473
rect 9769 14433 9781 14467
rect 9815 14464 9827 14467
rect 10229 14467 10287 14473
rect 10229 14464 10241 14467
rect 9815 14436 10241 14464
rect 9815 14433 9827 14436
rect 9769 14427 9827 14433
rect 10229 14433 10241 14436
rect 10275 14433 10287 14467
rect 10612 14464 10640 14504
rect 11238 14492 11244 14504
rect 11296 14532 11302 14544
rect 11514 14532 11520 14544
rect 11296 14504 11520 14532
rect 11296 14492 11302 14504
rect 11514 14492 11520 14504
rect 11572 14492 11578 14544
rect 11606 14492 11612 14544
rect 11664 14532 11670 14544
rect 11664 14504 12020 14532
rect 11664 14492 11670 14504
rect 11790 14464 11796 14476
rect 10229 14427 10287 14433
rect 10520 14436 10640 14464
rect 10704 14436 11796 14464
rect 5353 14399 5411 14405
rect 5184 14368 5304 14396
rect 5166 14328 5172 14340
rect 4356 14300 5172 14328
rect 5166 14288 5172 14300
rect 5224 14288 5230 14340
rect 5276 14337 5304 14368
rect 5353 14365 5365 14399
rect 5399 14396 5411 14399
rect 5718 14396 5724 14408
rect 5399 14368 5724 14396
rect 5399 14365 5411 14368
rect 5353 14359 5411 14365
rect 5718 14356 5724 14368
rect 5776 14356 5782 14408
rect 5810 14356 5816 14408
rect 5868 14396 5874 14408
rect 5997 14399 6055 14405
rect 5997 14396 6009 14399
rect 5868 14368 6009 14396
rect 5868 14356 5874 14368
rect 5997 14365 6009 14368
rect 6043 14365 6055 14399
rect 5997 14359 6055 14365
rect 6181 14399 6239 14405
rect 6181 14365 6193 14399
rect 6227 14365 6239 14399
rect 6181 14359 6239 14365
rect 7377 14399 7435 14405
rect 7377 14365 7389 14399
rect 7423 14396 7435 14399
rect 8018 14396 8024 14408
rect 7423 14368 8024 14396
rect 7423 14365 7435 14368
rect 7377 14359 7435 14365
rect 5261 14331 5319 14337
rect 5261 14297 5273 14331
rect 5307 14297 5319 14331
rect 6196 14328 6224 14359
rect 8018 14356 8024 14368
rect 8076 14356 8082 14408
rect 9214 14356 9220 14408
rect 9272 14405 9278 14408
rect 9272 14399 9308 14405
rect 9296 14365 9308 14399
rect 9674 14396 9680 14408
rect 9587 14368 9680 14396
rect 9272 14359 9308 14365
rect 9272 14356 9278 14359
rect 9674 14356 9680 14368
rect 9732 14396 9738 14408
rect 9950 14396 9956 14408
rect 9732 14368 9956 14396
rect 9732 14356 9738 14368
rect 9950 14356 9956 14368
rect 10008 14356 10014 14408
rect 10520 14405 10548 14436
rect 10704 14405 10732 14436
rect 11790 14424 11796 14436
rect 11848 14424 11854 14476
rect 11992 14473 12020 14504
rect 11977 14467 12035 14473
rect 11977 14433 11989 14467
rect 12023 14433 12035 14467
rect 11977 14427 12035 14433
rect 12084 14464 12112 14572
rect 12158 14560 12164 14612
rect 12216 14600 12222 14612
rect 12437 14603 12495 14609
rect 12437 14600 12449 14603
rect 12216 14572 12449 14600
rect 12216 14560 12222 14572
rect 12437 14569 12449 14572
rect 12483 14569 12495 14603
rect 12437 14563 12495 14569
rect 14274 14560 14280 14612
rect 14332 14600 14338 14612
rect 14826 14600 14832 14612
rect 14332 14572 14832 14600
rect 14332 14560 14338 14572
rect 14826 14560 14832 14572
rect 14884 14600 14890 14612
rect 15470 14600 15476 14612
rect 14884 14572 15476 14600
rect 14884 14560 14890 14572
rect 15470 14560 15476 14572
rect 15528 14600 15534 14612
rect 15565 14603 15623 14609
rect 15565 14600 15577 14603
rect 15528 14572 15577 14600
rect 15528 14560 15534 14572
rect 15565 14569 15577 14572
rect 15611 14569 15623 14603
rect 19610 14600 19616 14612
rect 15565 14563 15623 14569
rect 15856 14572 19616 14600
rect 15562 14464 15568 14476
rect 12084 14436 15568 14464
rect 10505 14399 10563 14405
rect 10505 14365 10517 14399
rect 10551 14365 10563 14399
rect 10505 14359 10563 14365
rect 10597 14399 10655 14405
rect 10597 14365 10609 14399
rect 10643 14365 10655 14399
rect 10597 14359 10655 14365
rect 10689 14399 10747 14405
rect 10689 14365 10701 14399
rect 10735 14365 10747 14399
rect 10689 14359 10747 14365
rect 7282 14328 7288 14340
rect 6196 14300 7288 14328
rect 5261 14291 5319 14297
rect 7282 14288 7288 14300
rect 7340 14288 7346 14340
rect 8113 14331 8171 14337
rect 8113 14328 8125 14331
rect 7484 14300 8125 14328
rect 7484 14272 7512 14300
rect 8113 14297 8125 14300
rect 8159 14297 8171 14331
rect 10612 14328 10640 14359
rect 10778 14356 10784 14408
rect 10836 14396 10842 14408
rect 10873 14399 10931 14405
rect 10873 14396 10885 14399
rect 10836 14368 10885 14396
rect 10836 14356 10842 14368
rect 10873 14365 10885 14368
rect 10919 14365 10931 14399
rect 11698 14396 11704 14408
rect 11659 14368 11704 14396
rect 10873 14359 10931 14365
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 12084 14405 12112 14436
rect 15562 14424 15568 14436
rect 15620 14424 15626 14476
rect 15856 14464 15884 14572
rect 19610 14560 19616 14572
rect 19668 14560 19674 14612
rect 16298 14492 16304 14544
rect 16356 14532 16362 14544
rect 16485 14535 16543 14541
rect 16485 14532 16497 14535
rect 16356 14504 16497 14532
rect 16356 14492 16362 14504
rect 16485 14501 16497 14504
rect 16531 14501 16543 14535
rect 16485 14495 16543 14501
rect 18509 14467 18567 14473
rect 18509 14464 18521 14467
rect 15764 14436 15884 14464
rect 16500 14436 18521 14464
rect 11885 14399 11943 14405
rect 11885 14365 11897 14399
rect 11931 14365 11943 14399
rect 11885 14359 11943 14365
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14365 12127 14399
rect 12069 14359 12127 14365
rect 12253 14399 12311 14405
rect 12253 14365 12265 14399
rect 12299 14396 12311 14399
rect 13170 14396 13176 14408
rect 12299 14368 13176 14396
rect 12299 14365 12311 14368
rect 12253 14359 12311 14365
rect 11330 14328 11336 14340
rect 10612 14300 11336 14328
rect 8113 14291 8171 14297
rect 11330 14288 11336 14300
rect 11388 14288 11394 14340
rect 11900 14328 11928 14359
rect 13170 14356 13176 14368
rect 13228 14356 13234 14408
rect 13354 14396 13360 14408
rect 13315 14368 13360 14396
rect 13354 14356 13360 14368
rect 13412 14356 13418 14408
rect 13630 14396 13636 14408
rect 13543 14368 13636 14396
rect 13630 14356 13636 14368
rect 13688 14396 13694 14408
rect 14090 14396 14096 14408
rect 13688 14368 14096 14396
rect 13688 14356 13694 14368
rect 14090 14356 14096 14368
rect 14148 14356 14154 14408
rect 14550 14356 14556 14408
rect 14608 14396 14614 14408
rect 15473 14399 15531 14405
rect 15473 14396 15485 14399
rect 14608 14368 15485 14396
rect 14608 14356 14614 14368
rect 15473 14365 15485 14368
rect 15519 14396 15531 14399
rect 15764 14396 15792 14436
rect 16500 14408 16528 14436
rect 18509 14433 18521 14436
rect 18555 14433 18567 14467
rect 18509 14427 18567 14433
rect 15519 14368 15792 14396
rect 15841 14399 15899 14405
rect 15519 14365 15531 14368
rect 15473 14359 15531 14365
rect 15841 14365 15853 14399
rect 15887 14396 15899 14399
rect 16206 14396 16212 14408
rect 15887 14368 16212 14396
rect 15887 14365 15899 14368
rect 15841 14359 15899 14365
rect 16206 14356 16212 14368
rect 16264 14356 16270 14408
rect 16482 14396 16488 14408
rect 16443 14368 16488 14396
rect 16482 14356 16488 14368
rect 16540 14356 16546 14408
rect 16666 14396 16672 14408
rect 16627 14368 16672 14396
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 18230 14396 18236 14408
rect 18191 14368 18236 14396
rect 18230 14356 18236 14368
rect 18288 14356 18294 14408
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14396 18383 14399
rect 18414 14396 18420 14408
rect 18371 14368 18420 14396
rect 18371 14365 18383 14368
rect 18325 14359 18383 14365
rect 18414 14356 18420 14368
rect 18472 14356 18478 14408
rect 14458 14328 14464 14340
rect 11900 14300 14464 14328
rect 14458 14288 14464 14300
rect 14516 14288 14522 14340
rect 18874 14328 18880 14340
rect 14568 14300 18880 14328
rect 5074 14260 5080 14272
rect 2832 14232 2877 14260
rect 4264 14232 5080 14260
rect 2832 14220 2838 14232
rect 5074 14220 5080 14232
rect 5132 14220 5138 14272
rect 5534 14260 5540 14272
rect 5495 14232 5540 14260
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 6917 14263 6975 14269
rect 6917 14229 6929 14263
rect 6963 14260 6975 14263
rect 7466 14260 7472 14272
rect 6963 14232 7472 14260
rect 6963 14229 6975 14232
rect 6917 14223 6975 14229
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 9306 14260 9312 14272
rect 9267 14232 9312 14260
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 13078 14220 13084 14272
rect 13136 14260 13142 14272
rect 13173 14263 13231 14269
rect 13173 14260 13185 14263
rect 13136 14232 13185 14260
rect 13136 14220 13142 14232
rect 13173 14229 13185 14232
rect 13219 14229 13231 14263
rect 13173 14223 13231 14229
rect 13541 14263 13599 14269
rect 13541 14229 13553 14263
rect 13587 14260 13599 14263
rect 13722 14260 13728 14272
rect 13587 14232 13728 14260
rect 13587 14229 13599 14232
rect 13541 14223 13599 14229
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 13998 14220 14004 14272
rect 14056 14260 14062 14272
rect 14568 14260 14596 14300
rect 18874 14288 18880 14300
rect 18932 14288 18938 14340
rect 14056 14232 14596 14260
rect 14056 14220 14062 14232
rect 14642 14220 14648 14272
rect 14700 14260 14706 14272
rect 15286 14260 15292 14272
rect 14700 14232 15292 14260
rect 14700 14220 14706 14232
rect 15286 14220 15292 14232
rect 15344 14220 15350 14272
rect 15378 14220 15384 14272
rect 15436 14260 15442 14272
rect 16025 14263 16083 14269
rect 16025 14260 16037 14263
rect 15436 14232 16037 14260
rect 15436 14220 15442 14232
rect 16025 14229 16037 14232
rect 16071 14229 16083 14263
rect 16025 14223 16083 14229
rect 18046 14220 18052 14272
rect 18104 14260 18110 14272
rect 18509 14263 18567 14269
rect 18509 14260 18521 14263
rect 18104 14232 18521 14260
rect 18104 14220 18110 14232
rect 18509 14229 18521 14232
rect 18555 14229 18567 14263
rect 18509 14223 18567 14229
rect 1104 14170 21043 14192
rect 1104 14118 5894 14170
rect 5946 14118 5958 14170
rect 6010 14118 6022 14170
rect 6074 14118 6086 14170
rect 6138 14118 6150 14170
rect 6202 14118 10839 14170
rect 10891 14118 10903 14170
rect 10955 14118 10967 14170
rect 11019 14118 11031 14170
rect 11083 14118 11095 14170
rect 11147 14118 15784 14170
rect 15836 14118 15848 14170
rect 15900 14118 15912 14170
rect 15964 14118 15976 14170
rect 16028 14118 16040 14170
rect 16092 14118 20729 14170
rect 20781 14118 20793 14170
rect 20845 14118 20857 14170
rect 20909 14118 20921 14170
rect 20973 14118 20985 14170
rect 21037 14118 21043 14170
rect 1104 14096 21043 14118
rect 1946 14016 1952 14068
rect 2004 14056 2010 14068
rect 2041 14059 2099 14065
rect 2041 14056 2053 14059
rect 2004 14028 2053 14056
rect 2004 14016 2010 14028
rect 2041 14025 2053 14028
rect 2087 14025 2099 14059
rect 2041 14019 2099 14025
rect 2967 14059 3025 14065
rect 2967 14025 2979 14059
rect 3013 14056 3025 14059
rect 3326 14056 3332 14068
rect 3013 14028 3332 14056
rect 3013 14025 3025 14028
rect 2967 14019 3025 14025
rect 3326 14016 3332 14028
rect 3384 14016 3390 14068
rect 5166 14016 5172 14068
rect 5224 14056 5230 14068
rect 5353 14059 5411 14065
rect 5353 14056 5365 14059
rect 5224 14028 5365 14056
rect 5224 14016 5230 14028
rect 5353 14025 5365 14028
rect 5399 14025 5411 14059
rect 7006 14056 7012 14068
rect 5353 14019 5411 14025
rect 5460 14028 7012 14056
rect 2406 13948 2412 14000
rect 2464 13988 2470 14000
rect 3053 13991 3111 13997
rect 3053 13988 3065 13991
rect 2464 13960 3065 13988
rect 2464 13948 2470 13960
rect 3053 13957 3065 13960
rect 3099 13988 3111 13991
rect 5460 13988 5488 14028
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 7098 14016 7104 14068
rect 7156 14056 7162 14068
rect 9309 14059 9367 14065
rect 7156 14028 9168 14056
rect 7156 14016 7162 14028
rect 3099 13960 5488 13988
rect 3099 13957 3111 13960
rect 3053 13951 3111 13957
rect 6822 13948 6828 14000
rect 6880 13948 6886 14000
rect 6918 13991 6976 13997
rect 6918 13966 6930 13991
rect 6964 13966 6976 13991
rect 7282 13988 7288 14000
rect 6826 13945 6884 13948
rect 1949 13923 2007 13929
rect 1949 13889 1961 13923
rect 1995 13920 2007 13923
rect 2038 13920 2044 13932
rect 1995 13892 2044 13920
rect 1995 13889 2007 13892
rect 1949 13883 2007 13889
rect 2038 13880 2044 13892
rect 2096 13920 2102 13932
rect 2869 13923 2927 13929
rect 2096 13892 2544 13920
rect 2096 13880 2102 13892
rect 2225 13855 2283 13861
rect 2225 13821 2237 13855
rect 2271 13821 2283 13855
rect 2516 13852 2544 13892
rect 2869 13889 2881 13923
rect 2915 13920 2927 13923
rect 2915 13892 3096 13920
rect 2915 13889 2927 13892
rect 2869 13883 2927 13889
rect 2958 13852 2964 13864
rect 2516 13824 2964 13852
rect 2225 13815 2283 13821
rect 2240 13784 2268 13815
rect 2958 13812 2964 13824
rect 3016 13812 3022 13864
rect 3068 13852 3096 13892
rect 3142 13880 3148 13932
rect 3200 13920 3206 13932
rect 4985 13923 5043 13929
rect 3200 13892 3245 13920
rect 3200 13880 3206 13892
rect 4985 13889 4997 13923
rect 5031 13889 5043 13923
rect 4985 13883 5043 13889
rect 5169 13923 5227 13929
rect 5169 13889 5181 13923
rect 5215 13920 5227 13923
rect 5626 13920 5632 13932
rect 5215 13892 5632 13920
rect 5215 13889 5227 13892
rect 5169 13883 5227 13889
rect 3234 13852 3240 13864
rect 3068 13824 3240 13852
rect 3234 13812 3240 13824
rect 3292 13812 3298 13864
rect 5000 13852 5028 13883
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 5736 13892 6776 13920
rect 6826 13911 6838 13945
rect 6872 13911 6884 13945
rect 6914 13914 6920 13966
rect 6972 13914 6978 13966
rect 7024 13960 7288 13988
rect 7024 13929 7052 13960
rect 7282 13948 7288 13960
rect 7340 13948 7346 14000
rect 7190 13929 7196 13932
rect 7009 13923 7067 13929
rect 6826 13905 6884 13911
rect 5736 13864 5764 13892
rect 5718 13852 5724 13864
rect 5000 13824 5724 13852
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 6638 13852 6644 13864
rect 6599 13824 6644 13852
rect 6638 13812 6644 13824
rect 6696 13812 6702 13864
rect 6748 13852 6776 13892
rect 7009 13889 7021 13923
rect 7055 13889 7067 13923
rect 7009 13883 7067 13889
rect 7147 13923 7196 13929
rect 7147 13889 7159 13923
rect 7193 13889 7196 13923
rect 7147 13883 7196 13889
rect 7190 13880 7196 13883
rect 7248 13880 7254 13932
rect 7834 13920 7840 13932
rect 7795 13892 7840 13920
rect 7834 13880 7840 13892
rect 7892 13880 7898 13932
rect 8018 13920 8024 13932
rect 7979 13892 8024 13920
rect 8018 13880 8024 13892
rect 8076 13880 8082 13932
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13920 8999 13923
rect 9030 13920 9036 13932
rect 8987 13892 9036 13920
rect 8987 13889 8999 13892
rect 8941 13883 8999 13889
rect 9030 13880 9036 13892
rect 9088 13880 9094 13932
rect 7285 13855 7343 13861
rect 6748 13824 7236 13852
rect 2866 13784 2872 13796
rect 2240 13756 2872 13784
rect 2866 13744 2872 13756
rect 2924 13744 2930 13796
rect 7208 13784 7236 13824
rect 7285 13821 7297 13855
rect 7331 13852 7343 13855
rect 8849 13855 8907 13861
rect 7331 13824 7972 13852
rect 7331 13821 7343 13824
rect 7285 13815 7343 13821
rect 7944 13796 7972 13824
rect 8849 13821 8861 13855
rect 8895 13821 8907 13855
rect 9140 13852 9168 14028
rect 9309 14025 9321 14059
rect 9355 14056 9367 14059
rect 10686 14056 10692 14068
rect 9355 14028 10692 14056
rect 9355 14025 9367 14028
rect 9309 14019 9367 14025
rect 9876 13997 9904 14028
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 11885 14059 11943 14065
rect 11885 14025 11897 14059
rect 11931 14056 11943 14059
rect 12066 14056 12072 14068
rect 11931 14028 12072 14056
rect 11931 14025 11943 14028
rect 11885 14019 11943 14025
rect 12066 14016 12072 14028
rect 12124 14056 12130 14068
rect 13354 14056 13360 14068
rect 12124 14028 13360 14056
rect 12124 14016 12130 14028
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 15470 14016 15476 14068
rect 15528 14056 15534 14068
rect 15749 14059 15807 14065
rect 15749 14056 15761 14059
rect 15528 14028 15761 14056
rect 15528 14016 15534 14028
rect 15749 14025 15761 14028
rect 15795 14025 15807 14059
rect 15749 14019 15807 14025
rect 16482 14016 16488 14068
rect 16540 14056 16546 14068
rect 17313 14059 17371 14065
rect 17313 14056 17325 14059
rect 16540 14028 17325 14056
rect 16540 14016 16546 14028
rect 17313 14025 17325 14028
rect 17359 14025 17371 14059
rect 17313 14019 17371 14025
rect 9861 13991 9919 13997
rect 9861 13957 9873 13991
rect 9907 13957 9919 13991
rect 9861 13951 9919 13957
rect 10413 13991 10471 13997
rect 10413 13957 10425 13991
rect 10459 13988 10471 13991
rect 14001 13991 14059 13997
rect 10459 13960 13952 13988
rect 10459 13957 10471 13960
rect 10413 13951 10471 13957
rect 11900 13932 11928 13960
rect 9214 13880 9220 13932
rect 9272 13920 9278 13932
rect 10045 13923 10103 13929
rect 10045 13920 10057 13923
rect 9272 13892 10057 13920
rect 9272 13880 9278 13892
rect 10045 13889 10057 13892
rect 10091 13889 10103 13923
rect 10045 13883 10103 13889
rect 11882 13880 11888 13932
rect 11940 13880 11946 13932
rect 12894 13920 12900 13932
rect 12176 13892 12756 13920
rect 12855 13892 12900 13920
rect 11701 13855 11759 13861
rect 9140 13824 11652 13852
rect 8849 13815 8907 13821
rect 7837 13787 7895 13793
rect 7837 13784 7849 13787
rect 7208 13756 7849 13784
rect 7837 13753 7849 13756
rect 7883 13753 7895 13787
rect 7837 13747 7895 13753
rect 7926 13744 7932 13796
rect 7984 13744 7990 13796
rect 8864 13784 8892 13815
rect 8938 13784 8944 13796
rect 8864 13756 8944 13784
rect 8938 13744 8944 13756
rect 8996 13744 9002 13796
rect 11624 13784 11652 13824
rect 11701 13821 11713 13855
rect 11747 13852 11759 13855
rect 11790 13852 11796 13864
rect 11747 13824 11796 13852
rect 11747 13821 11759 13824
rect 11701 13815 11759 13821
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 12176 13861 12204 13892
rect 12161 13855 12219 13861
rect 12161 13852 12173 13855
rect 11900 13824 12173 13852
rect 11900 13784 11928 13824
rect 12161 13821 12173 13824
rect 12207 13821 12219 13855
rect 12161 13815 12219 13821
rect 12253 13855 12311 13861
rect 12253 13821 12265 13855
rect 12299 13852 12311 13855
rect 12342 13852 12348 13864
rect 12299 13824 12348 13852
rect 12299 13821 12311 13824
rect 12253 13815 12311 13821
rect 12342 13812 12348 13824
rect 12400 13812 12406 13864
rect 12728 13852 12756 13892
rect 12894 13880 12900 13892
rect 12952 13880 12958 13932
rect 13924 13920 13952 13960
rect 14001 13957 14013 13991
rect 14047 13988 14059 13991
rect 14047 13960 15240 13988
rect 14047 13957 14059 13960
rect 14001 13951 14059 13957
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 13924 13892 14289 13920
rect 14277 13889 14289 13892
rect 14323 13920 14335 13923
rect 14550 13920 14556 13932
rect 14323 13892 14556 13920
rect 14323 13889 14335 13892
rect 14277 13883 14335 13889
rect 14550 13880 14556 13892
rect 14608 13880 14614 13932
rect 14734 13920 14740 13932
rect 14695 13892 14740 13920
rect 14734 13880 14740 13892
rect 14792 13880 14798 13932
rect 15212 13929 15240 13960
rect 15286 13948 15292 14000
rect 15344 13988 15350 14000
rect 15381 13991 15439 13997
rect 15381 13988 15393 13991
rect 15344 13960 15393 13988
rect 15344 13948 15350 13960
rect 15381 13957 15393 13960
rect 15427 13957 15439 13991
rect 15654 13988 15660 14000
rect 15381 13951 15439 13957
rect 15488 13960 15660 13988
rect 15488 13929 15516 13960
rect 15654 13948 15660 13960
rect 15712 13948 15718 14000
rect 16390 13948 16396 14000
rect 16448 13988 16454 14000
rect 16853 13991 16911 13997
rect 16853 13988 16865 13991
rect 16448 13960 16865 13988
rect 16448 13948 16454 13960
rect 16853 13957 16865 13960
rect 16899 13957 16911 13991
rect 17328 13988 17356 14019
rect 17954 14016 17960 14068
rect 18012 14056 18018 14068
rect 18782 14056 18788 14068
rect 18012 14028 18788 14056
rect 18012 14016 18018 14028
rect 18782 14016 18788 14028
rect 18840 14016 18846 14068
rect 19429 14059 19487 14065
rect 19429 14025 19441 14059
rect 19475 14025 19487 14059
rect 19610 14056 19616 14068
rect 19571 14028 19616 14056
rect 19429 14019 19487 14025
rect 18966 13988 18972 14000
rect 17328 13960 17724 13988
rect 16853 13951 16911 13957
rect 15197 13923 15255 13929
rect 15197 13889 15209 13923
rect 15243 13889 15255 13923
rect 15197 13883 15255 13889
rect 15473 13923 15531 13929
rect 15473 13889 15485 13923
rect 15519 13889 15531 13923
rect 15473 13883 15531 13889
rect 15565 13923 15623 13929
rect 15565 13889 15577 13923
rect 15611 13920 15623 13923
rect 17494 13920 17500 13932
rect 15611 13892 17500 13920
rect 15611 13889 15623 13892
rect 15565 13883 15623 13889
rect 17494 13880 17500 13892
rect 17552 13880 17558 13932
rect 13998 13852 14004 13864
rect 12728 13824 14004 13852
rect 13998 13812 14004 13824
rect 14056 13812 14062 13864
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13852 14427 13855
rect 17696 13852 17724 13960
rect 18524 13960 18972 13988
rect 17954 13880 17960 13932
rect 18012 13920 18018 13932
rect 18230 13920 18236 13932
rect 18012 13892 18236 13920
rect 18012 13880 18018 13892
rect 18230 13880 18236 13892
rect 18288 13920 18294 13932
rect 18325 13923 18383 13929
rect 18325 13920 18337 13923
rect 18288 13892 18337 13920
rect 18288 13880 18294 13892
rect 18325 13889 18337 13892
rect 18371 13889 18383 13923
rect 18325 13883 18383 13889
rect 18414 13880 18420 13932
rect 18472 13920 18478 13932
rect 18524 13920 18552 13960
rect 18966 13948 18972 13960
rect 19024 13988 19030 14000
rect 19444 13988 19472 14019
rect 19610 14016 19616 14028
rect 19668 14016 19674 14068
rect 19024 13960 19472 13988
rect 19024 13948 19030 13960
rect 18637 13923 18695 13929
rect 18472 13892 18565 13920
rect 18472 13880 18478 13892
rect 18637 13889 18649 13923
rect 18683 13920 18695 13923
rect 18782 13920 18788 13932
rect 18683 13892 18788 13920
rect 18683 13889 18695 13892
rect 18637 13883 18695 13889
rect 18782 13880 18788 13892
rect 18840 13880 18846 13932
rect 19554 13923 19612 13929
rect 19554 13920 19566 13923
rect 19306 13892 19566 13920
rect 18509 13855 18567 13861
rect 18509 13852 18521 13855
rect 14415 13824 14596 13852
rect 17696 13824 18521 13852
rect 14415 13821 14427 13824
rect 14369 13815 14427 13821
rect 14458 13784 14464 13796
rect 11624 13756 11928 13784
rect 13004 13756 14044 13784
rect 14419 13756 14464 13784
rect 1578 13716 1584 13728
rect 1539 13688 1584 13716
rect 1578 13676 1584 13688
rect 1636 13676 1642 13728
rect 10410 13676 10416 13728
rect 10468 13716 10474 13728
rect 13004 13716 13032 13756
rect 10468 13688 13032 13716
rect 13081 13719 13139 13725
rect 10468 13676 10474 13688
rect 13081 13685 13093 13719
rect 13127 13716 13139 13719
rect 13170 13716 13176 13728
rect 13127 13688 13176 13716
rect 13127 13685 13139 13688
rect 13081 13679 13139 13685
rect 13170 13676 13176 13688
rect 13228 13676 13234 13728
rect 14016 13716 14044 13756
rect 14458 13744 14464 13756
rect 14516 13744 14522 13796
rect 14568 13784 14596 13824
rect 18509 13821 18521 13824
rect 18555 13821 18567 13855
rect 18509 13815 18567 13821
rect 15194 13784 15200 13796
rect 14568 13756 15200 13784
rect 15194 13744 15200 13756
rect 15252 13784 15258 13796
rect 16298 13784 16304 13796
rect 15252 13756 16304 13784
rect 15252 13744 15258 13756
rect 16298 13744 16304 13756
rect 16356 13744 16362 13796
rect 17126 13784 17132 13796
rect 17039 13756 17132 13784
rect 17126 13744 17132 13756
rect 17184 13784 17190 13796
rect 19306 13784 19334 13892
rect 19554 13889 19566 13892
rect 19600 13920 19612 13923
rect 19794 13920 19800 13932
rect 19600 13892 19800 13920
rect 19600 13889 19612 13892
rect 19554 13883 19612 13889
rect 19794 13880 19800 13892
rect 19852 13880 19858 13932
rect 20070 13852 20076 13864
rect 20031 13824 20076 13852
rect 20070 13812 20076 13824
rect 20128 13812 20134 13864
rect 19978 13784 19984 13796
rect 17184 13756 19334 13784
rect 19939 13756 19984 13784
rect 17184 13744 17190 13756
rect 19978 13744 19984 13756
rect 20036 13744 20042 13796
rect 14182 13716 14188 13728
rect 14016 13688 14188 13716
rect 14182 13676 14188 13688
rect 14240 13716 14246 13728
rect 14550 13716 14556 13728
rect 14240 13688 14556 13716
rect 14240 13676 14246 13688
rect 14550 13676 14556 13688
rect 14608 13676 14614 13728
rect 14642 13676 14648 13728
rect 14700 13716 14706 13728
rect 15010 13716 15016 13728
rect 14700 13688 15016 13716
rect 14700 13676 14706 13688
rect 15010 13676 15016 13688
rect 15068 13716 15074 13728
rect 17144 13716 17172 13744
rect 18138 13716 18144 13728
rect 15068 13688 17172 13716
rect 18099 13688 18144 13716
rect 15068 13676 15074 13688
rect 18138 13676 18144 13688
rect 18196 13676 18202 13728
rect 1104 13626 20884 13648
rect 1104 13574 3422 13626
rect 3474 13574 3486 13626
rect 3538 13574 3550 13626
rect 3602 13574 3614 13626
rect 3666 13574 3678 13626
rect 3730 13574 8367 13626
rect 8419 13574 8431 13626
rect 8483 13574 8495 13626
rect 8547 13574 8559 13626
rect 8611 13574 8623 13626
rect 8675 13574 13312 13626
rect 13364 13574 13376 13626
rect 13428 13574 13440 13626
rect 13492 13574 13504 13626
rect 13556 13574 13568 13626
rect 13620 13574 18257 13626
rect 18309 13574 18321 13626
rect 18373 13574 18385 13626
rect 18437 13574 18449 13626
rect 18501 13574 18513 13626
rect 18565 13574 20884 13626
rect 1104 13552 20884 13574
rect 7558 13512 7564 13524
rect 7519 13484 7564 13512
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 9217 13515 9275 13521
rect 9217 13481 9229 13515
rect 9263 13512 9275 13515
rect 9306 13512 9312 13524
rect 9263 13484 9312 13512
rect 9263 13481 9275 13484
rect 9217 13475 9275 13481
rect 9306 13472 9312 13484
rect 9364 13472 9370 13524
rect 12894 13472 12900 13524
rect 12952 13512 12958 13524
rect 13541 13515 13599 13521
rect 13541 13512 13553 13515
rect 12952 13484 13553 13512
rect 12952 13472 12958 13484
rect 13541 13481 13553 13484
rect 13587 13481 13599 13515
rect 13541 13475 13599 13481
rect 14277 13515 14335 13521
rect 14277 13481 14289 13515
rect 14323 13512 14335 13515
rect 14458 13512 14464 13524
rect 14323 13484 14464 13512
rect 14323 13481 14335 13484
rect 14277 13475 14335 13481
rect 14458 13472 14464 13484
rect 14516 13472 14522 13524
rect 17494 13512 17500 13524
rect 17455 13484 17500 13512
rect 17494 13472 17500 13484
rect 17552 13472 17558 13524
rect 2958 13404 2964 13456
rect 3016 13444 3022 13456
rect 3234 13444 3240 13456
rect 3016 13416 3240 13444
rect 3016 13404 3022 13416
rect 3234 13404 3240 13416
rect 3292 13444 3298 13456
rect 11606 13444 11612 13456
rect 3292 13416 4936 13444
rect 11567 13416 11612 13444
rect 3292 13404 3298 13416
rect 4908 13388 4936 13416
rect 11606 13404 11612 13416
rect 11664 13404 11670 13456
rect 4706 13376 4712 13388
rect 4667 13348 4712 13376
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 4890 13376 4896 13388
rect 4851 13348 4896 13376
rect 4890 13336 4896 13348
rect 4948 13336 4954 13388
rect 8938 13336 8944 13388
rect 8996 13376 9002 13388
rect 12342 13376 12348 13388
rect 8996 13348 12348 13376
rect 8996 13336 9002 13348
rect 2038 13268 2044 13320
rect 2096 13308 2102 13320
rect 2225 13311 2283 13317
rect 2225 13308 2237 13311
rect 2096 13280 2237 13308
rect 2096 13268 2102 13280
rect 2225 13277 2237 13280
rect 2271 13277 2283 13311
rect 2225 13271 2283 13277
rect 5626 13268 5632 13320
rect 5684 13308 5690 13320
rect 6822 13308 6828 13320
rect 5684 13280 6828 13308
rect 5684 13268 5690 13280
rect 6822 13268 6828 13280
rect 6880 13308 6886 13320
rect 7469 13311 7527 13317
rect 7469 13308 7481 13311
rect 6880 13280 7481 13308
rect 6880 13268 6886 13280
rect 7469 13277 7481 13280
rect 7515 13277 7527 13311
rect 9122 13308 9128 13320
rect 9083 13280 9128 13308
rect 7469 13271 7527 13277
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 11256 13317 11284 13348
rect 12342 13336 12348 13348
rect 12400 13336 12406 13388
rect 14918 13376 14924 13388
rect 14292 13348 14924 13376
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13277 9367 13311
rect 9309 13271 9367 13277
rect 11241 13311 11299 13317
rect 11241 13277 11253 13311
rect 11287 13277 11299 13311
rect 11241 13271 11299 13277
rect 11395 13311 11453 13317
rect 11395 13277 11407 13311
rect 11441 13308 11453 13311
rect 11790 13308 11796 13320
rect 11441 13280 11796 13308
rect 11441 13277 11453 13280
rect 11395 13271 11453 13277
rect 2685 13243 2743 13249
rect 2685 13209 2697 13243
rect 2731 13240 2743 13243
rect 2866 13240 2872 13252
rect 2731 13212 2872 13240
rect 2731 13209 2743 13212
rect 2685 13203 2743 13209
rect 2866 13200 2872 13212
rect 2924 13240 2930 13252
rect 4062 13240 4068 13252
rect 2924 13212 4068 13240
rect 2924 13200 2930 13212
rect 4062 13200 4068 13212
rect 4120 13200 4126 13252
rect 8202 13200 8208 13252
rect 8260 13240 8266 13252
rect 9324 13240 9352 13271
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 12066 13268 12072 13320
rect 12124 13308 12130 13320
rect 14292 13317 14320 13348
rect 14918 13336 14924 13348
rect 14976 13376 14982 13388
rect 15378 13376 15384 13388
rect 14976 13348 15384 13376
rect 14976 13336 14982 13348
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 18138 13376 18144 13388
rect 18099 13348 18144 13376
rect 18138 13336 18144 13348
rect 18196 13336 18202 13388
rect 13449 13311 13507 13317
rect 13449 13308 13461 13311
rect 12124 13280 13461 13308
rect 12124 13268 12130 13280
rect 13449 13277 13461 13280
rect 13495 13277 13507 13311
rect 13449 13271 13507 13277
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 14461 13311 14519 13317
rect 14461 13277 14473 13311
rect 14507 13277 14519 13311
rect 14461 13271 14519 13277
rect 10686 13240 10692 13252
rect 8260 13212 10692 13240
rect 8260 13200 8266 13212
rect 10686 13200 10692 13212
rect 10744 13200 10750 13252
rect 14476 13240 14504 13271
rect 16850 13268 16856 13320
rect 16908 13308 16914 13320
rect 17681 13311 17739 13317
rect 17681 13308 17693 13311
rect 16908 13280 17693 13308
rect 16908 13268 16914 13280
rect 17681 13277 17693 13280
rect 17727 13277 17739 13311
rect 17681 13271 17739 13277
rect 17770 13268 17776 13320
rect 17828 13308 17834 13320
rect 18046 13308 18052 13320
rect 17828 13280 17873 13308
rect 18007 13280 18052 13308
rect 17828 13268 17834 13280
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 19886 13308 19892 13320
rect 19847 13280 19892 13308
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 19981 13243 20039 13249
rect 19981 13240 19993 13243
rect 14476 13212 19993 13240
rect 19981 13209 19993 13212
rect 20027 13240 20039 13243
rect 20070 13240 20076 13252
rect 20027 13212 20076 13240
rect 20027 13209 20039 13212
rect 19981 13203 20039 13209
rect 20070 13200 20076 13212
rect 20128 13200 20134 13252
rect 4154 13132 4160 13184
rect 4212 13172 4218 13184
rect 4249 13175 4307 13181
rect 4249 13172 4261 13175
rect 4212 13144 4261 13172
rect 4212 13132 4218 13144
rect 4249 13141 4261 13144
rect 4295 13141 4307 13175
rect 4614 13172 4620 13184
rect 4575 13144 4620 13172
rect 4249 13135 4307 13141
rect 4614 13132 4620 13144
rect 4672 13132 4678 13184
rect 1104 13082 21043 13104
rect 1104 13030 5894 13082
rect 5946 13030 5958 13082
rect 6010 13030 6022 13082
rect 6074 13030 6086 13082
rect 6138 13030 6150 13082
rect 6202 13030 10839 13082
rect 10891 13030 10903 13082
rect 10955 13030 10967 13082
rect 11019 13030 11031 13082
rect 11083 13030 11095 13082
rect 11147 13030 15784 13082
rect 15836 13030 15848 13082
rect 15900 13030 15912 13082
rect 15964 13030 15976 13082
rect 16028 13030 16040 13082
rect 16092 13030 20729 13082
rect 20781 13030 20793 13082
rect 20845 13030 20857 13082
rect 20909 13030 20921 13082
rect 20973 13030 20985 13082
rect 21037 13030 21043 13082
rect 1104 13008 21043 13030
rect 4154 12968 4160 12980
rect 4115 12940 4160 12968
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 5353 12971 5411 12977
rect 5353 12937 5365 12971
rect 5399 12968 5411 12971
rect 5534 12968 5540 12980
rect 5399 12940 5540 12968
rect 5399 12937 5411 12940
rect 5353 12931 5411 12937
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 6825 12971 6883 12977
rect 6825 12937 6837 12971
rect 6871 12968 6883 12971
rect 7098 12968 7104 12980
rect 6871 12940 7104 12968
rect 6871 12937 6883 12940
rect 6825 12931 6883 12937
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 13170 12928 13176 12980
rect 13228 12928 13234 12980
rect 15562 12928 15568 12980
rect 15620 12968 15626 12980
rect 15841 12971 15899 12977
rect 15841 12968 15853 12971
rect 15620 12940 15853 12968
rect 15620 12928 15626 12940
rect 15841 12937 15853 12940
rect 15887 12937 15899 12971
rect 16850 12968 16856 12980
rect 16811 12940 16856 12968
rect 15841 12931 15899 12937
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 18601 12971 18659 12977
rect 18601 12937 18613 12971
rect 18647 12968 18659 12971
rect 20073 12971 20131 12977
rect 20073 12968 20085 12971
rect 18647 12940 20085 12968
rect 18647 12937 18659 12940
rect 18601 12931 18659 12937
rect 20073 12937 20085 12940
rect 20119 12937 20131 12971
rect 20073 12931 20131 12937
rect 4246 12860 4252 12912
rect 4304 12860 4310 12912
rect 4338 12860 4344 12912
rect 4396 12900 4402 12912
rect 9214 12900 9220 12912
rect 4396 12872 9220 12900
rect 4396 12860 4402 12872
rect 9214 12860 9220 12872
rect 9272 12860 9278 12912
rect 10686 12860 10692 12912
rect 10744 12900 10750 12912
rect 13188 12900 13216 12928
rect 18616 12900 18644 12931
rect 10744 12872 13400 12900
rect 10744 12860 10750 12872
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12832 2559 12835
rect 3326 12832 3332 12844
rect 2547 12804 3332 12832
rect 2547 12801 2559 12804
rect 2501 12795 2559 12801
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 4065 12835 4123 12841
rect 4065 12801 4077 12835
rect 4111 12832 4123 12835
rect 4264 12832 4292 12860
rect 5261 12835 5319 12841
rect 5261 12832 5273 12835
rect 4111 12804 5273 12832
rect 4111 12801 4123 12804
rect 4065 12795 4123 12801
rect 5261 12801 5273 12804
rect 5307 12832 5319 12835
rect 5350 12832 5356 12844
rect 5307 12804 5356 12832
rect 5307 12801 5319 12804
rect 5261 12795 5319 12801
rect 5350 12792 5356 12804
rect 5408 12792 5414 12844
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 6641 12835 6699 12841
rect 6641 12832 6653 12835
rect 5776 12804 6653 12832
rect 5776 12792 5782 12804
rect 6641 12801 6653 12804
rect 6687 12801 6699 12835
rect 6641 12795 6699 12801
rect 6914 12792 6920 12844
rect 6972 12832 6978 12844
rect 7009 12835 7067 12841
rect 7009 12832 7021 12835
rect 6972 12804 7021 12832
rect 6972 12792 6978 12804
rect 7009 12801 7021 12804
rect 7055 12801 7067 12835
rect 7190 12832 7196 12844
rect 7151 12804 7196 12832
rect 7009 12795 7067 12801
rect 7190 12792 7196 12804
rect 7248 12832 7254 12844
rect 7374 12832 7380 12844
rect 7248 12804 7380 12832
rect 7248 12792 7254 12804
rect 7374 12792 7380 12804
rect 7432 12792 7438 12844
rect 9030 12832 9036 12844
rect 8991 12804 9036 12832
rect 9030 12792 9036 12804
rect 9088 12832 9094 12844
rect 9398 12832 9404 12844
rect 9088 12804 9404 12832
rect 9088 12792 9094 12804
rect 9398 12792 9404 12804
rect 9456 12792 9462 12844
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12832 11759 12835
rect 13170 12832 13176 12844
rect 11747 12804 13176 12832
rect 11747 12801 11759 12804
rect 11701 12795 11759 12801
rect 13170 12792 13176 12804
rect 13228 12792 13234 12844
rect 13372 12841 13400 12872
rect 17236 12872 18644 12900
rect 17236 12844 17264 12872
rect 13357 12835 13415 12841
rect 13357 12801 13369 12835
rect 13403 12801 13415 12835
rect 13357 12795 13415 12801
rect 14918 12792 14924 12844
rect 14976 12832 14982 12844
rect 15749 12835 15807 12841
rect 15749 12832 15761 12835
rect 14976 12804 15761 12832
rect 14976 12792 14982 12804
rect 15749 12801 15761 12804
rect 15795 12801 15807 12835
rect 16022 12832 16028 12844
rect 15983 12804 16028 12832
rect 15749 12795 15807 12801
rect 16022 12792 16028 12804
rect 16080 12792 16086 12844
rect 16666 12792 16672 12844
rect 16724 12832 16730 12844
rect 17129 12835 17187 12841
rect 17129 12832 17141 12835
rect 16724 12804 17141 12832
rect 16724 12792 16730 12804
rect 17129 12801 17141 12804
rect 17175 12801 17187 12835
rect 17129 12795 17187 12801
rect 17218 12792 17224 12844
rect 17276 12832 17282 12844
rect 17276 12804 17369 12832
rect 17276 12792 17282 12804
rect 17954 12792 17960 12844
rect 18012 12832 18018 12844
rect 18417 12835 18475 12841
rect 18417 12832 18429 12835
rect 18012 12804 18429 12832
rect 18012 12792 18018 12804
rect 18417 12801 18429 12804
rect 18463 12801 18475 12835
rect 18417 12795 18475 12801
rect 18598 12792 18604 12844
rect 18656 12832 18662 12844
rect 18693 12835 18751 12841
rect 18693 12832 18705 12835
rect 18656 12804 18705 12832
rect 18656 12792 18662 12804
rect 18693 12801 18705 12804
rect 18739 12801 18751 12835
rect 18693 12795 18751 12801
rect 19518 12792 19524 12844
rect 19576 12832 19582 12844
rect 19705 12835 19763 12841
rect 19705 12832 19717 12835
rect 19576 12804 19717 12832
rect 19576 12792 19582 12804
rect 19705 12801 19717 12804
rect 19751 12801 19763 12835
rect 19886 12832 19892 12844
rect 19847 12804 19892 12832
rect 19705 12795 19763 12801
rect 19886 12792 19892 12804
rect 19944 12792 19950 12844
rect 2038 12724 2044 12776
rect 2096 12764 2102 12776
rect 3053 12767 3111 12773
rect 3053 12764 3065 12767
rect 2096 12736 3065 12764
rect 2096 12724 2102 12736
rect 3053 12733 3065 12736
rect 3099 12764 3111 12767
rect 4249 12767 4307 12773
rect 4249 12764 4261 12767
rect 3099 12736 4016 12764
rect 3099 12733 3111 12736
rect 3053 12727 3111 12733
rect 3050 12588 3056 12640
rect 3108 12628 3114 12640
rect 3697 12631 3755 12637
rect 3697 12628 3709 12631
rect 3108 12600 3709 12628
rect 3108 12588 3114 12600
rect 3697 12597 3709 12600
rect 3743 12597 3755 12631
rect 3988 12628 4016 12736
rect 4080 12736 4261 12764
rect 4080 12708 4108 12736
rect 4249 12733 4261 12736
rect 4295 12733 4307 12767
rect 4249 12727 4307 12733
rect 4890 12724 4896 12776
rect 4948 12764 4954 12776
rect 5445 12767 5503 12773
rect 5445 12764 5457 12767
rect 4948 12736 5457 12764
rect 4948 12724 4954 12736
rect 5445 12733 5457 12736
rect 5491 12764 5503 12767
rect 7282 12764 7288 12776
rect 5491 12736 7288 12764
rect 5491 12733 5503 12736
rect 5445 12727 5503 12733
rect 7282 12724 7288 12736
rect 7340 12724 7346 12776
rect 8938 12764 8944 12776
rect 8899 12736 8944 12764
rect 8938 12724 8944 12736
rect 8996 12724 9002 12776
rect 9125 12767 9183 12773
rect 9125 12733 9137 12767
rect 9171 12733 9183 12767
rect 9125 12727 9183 12733
rect 4062 12656 4068 12708
rect 4120 12656 4126 12708
rect 4338 12628 4344 12640
rect 3988 12600 4344 12628
rect 3697 12591 3755 12597
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 4890 12628 4896 12640
rect 4851 12600 4896 12628
rect 4890 12588 4896 12600
rect 4948 12588 4954 12640
rect 7006 12628 7012 12640
rect 6967 12600 7012 12628
rect 7006 12588 7012 12600
rect 7064 12588 7070 12640
rect 8754 12628 8760 12640
rect 8715 12600 8760 12628
rect 8754 12588 8760 12600
rect 8812 12588 8818 12640
rect 9140 12628 9168 12727
rect 9214 12724 9220 12776
rect 9272 12764 9278 12776
rect 9272 12736 9317 12764
rect 9272 12724 9278 12736
rect 10502 12724 10508 12776
rect 10560 12764 10566 12776
rect 11977 12767 12035 12773
rect 11977 12764 11989 12767
rect 10560 12736 11989 12764
rect 10560 12724 10566 12736
rect 11977 12733 11989 12736
rect 12023 12733 12035 12767
rect 11977 12727 12035 12733
rect 12986 12724 12992 12776
rect 13044 12764 13050 12776
rect 13541 12767 13599 12773
rect 13541 12764 13553 12767
rect 13044 12736 13553 12764
rect 13044 12724 13050 12736
rect 13541 12733 13553 12736
rect 13587 12733 13599 12767
rect 13541 12727 13599 12733
rect 16574 12724 16580 12776
rect 16632 12764 16638 12776
rect 17037 12767 17095 12773
rect 17037 12764 17049 12767
rect 16632 12736 17049 12764
rect 16632 12724 16638 12736
rect 17037 12733 17049 12736
rect 17083 12733 17095 12767
rect 17037 12727 17095 12733
rect 17313 12767 17371 12773
rect 17313 12733 17325 12767
rect 17359 12764 17371 12767
rect 17862 12764 17868 12776
rect 17359 12736 17868 12764
rect 17359 12733 17371 12736
rect 17313 12727 17371 12733
rect 11793 12699 11851 12705
rect 11793 12665 11805 12699
rect 11839 12696 11851 12699
rect 12066 12696 12072 12708
rect 11839 12668 12072 12696
rect 11839 12665 11851 12668
rect 11793 12659 11851 12665
rect 12066 12656 12072 12668
rect 12124 12656 12130 12708
rect 14550 12656 14556 12708
rect 14608 12696 14614 12708
rect 17328 12696 17356 12727
rect 17862 12724 17868 12736
rect 17920 12724 17926 12776
rect 14608 12668 17356 12696
rect 18417 12699 18475 12705
rect 14608 12656 14614 12668
rect 18417 12665 18429 12699
rect 18463 12696 18475 12699
rect 18690 12696 18696 12708
rect 18463 12668 18696 12696
rect 18463 12665 18475 12668
rect 18417 12659 18475 12665
rect 18690 12656 18696 12668
rect 18748 12656 18754 12708
rect 9214 12628 9220 12640
rect 9140 12600 9220 12628
rect 9214 12588 9220 12600
rect 9272 12588 9278 12640
rect 11698 12628 11704 12640
rect 11659 12600 11704 12628
rect 11698 12588 11704 12600
rect 11756 12588 11762 12640
rect 14734 12588 14740 12640
rect 14792 12628 14798 12640
rect 15286 12628 15292 12640
rect 14792 12600 15292 12628
rect 14792 12588 14798 12600
rect 15286 12588 15292 12600
rect 15344 12588 15350 12640
rect 19702 12628 19708 12640
rect 19663 12600 19708 12628
rect 19702 12588 19708 12600
rect 19760 12588 19766 12640
rect 1104 12538 20884 12560
rect 1104 12486 3422 12538
rect 3474 12486 3486 12538
rect 3538 12486 3550 12538
rect 3602 12486 3614 12538
rect 3666 12486 3678 12538
rect 3730 12486 8367 12538
rect 8419 12486 8431 12538
rect 8483 12486 8495 12538
rect 8547 12486 8559 12538
rect 8611 12486 8623 12538
rect 8675 12486 13312 12538
rect 13364 12486 13376 12538
rect 13428 12486 13440 12538
rect 13492 12486 13504 12538
rect 13556 12486 13568 12538
rect 13620 12486 18257 12538
rect 18309 12486 18321 12538
rect 18373 12486 18385 12538
rect 18437 12486 18449 12538
rect 18501 12486 18513 12538
rect 18565 12486 20884 12538
rect 1104 12464 20884 12486
rect 4062 12384 4068 12436
rect 4120 12424 4126 12436
rect 5442 12424 5448 12436
rect 4120 12396 5448 12424
rect 4120 12384 4126 12396
rect 5442 12384 5448 12396
rect 5500 12384 5506 12436
rect 9122 12424 9128 12436
rect 9083 12396 9128 12424
rect 9122 12384 9128 12396
rect 9180 12384 9186 12436
rect 9398 12384 9404 12436
rect 9456 12424 9462 12436
rect 10502 12424 10508 12436
rect 9456 12396 10508 12424
rect 9456 12384 9462 12396
rect 10502 12384 10508 12396
rect 10560 12384 10566 12436
rect 10686 12384 10692 12436
rect 10744 12424 10750 12436
rect 11241 12427 11299 12433
rect 11241 12424 11253 12427
rect 10744 12396 11253 12424
rect 10744 12384 10750 12396
rect 11241 12393 11253 12396
rect 11287 12393 11299 12427
rect 11790 12424 11796 12436
rect 11751 12396 11796 12424
rect 11241 12387 11299 12393
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 13262 12424 13268 12436
rect 12636 12396 13268 12424
rect 6638 12356 6644 12368
rect 2332 12328 6644 12356
rect 2332 12297 2360 12328
rect 6638 12316 6644 12328
rect 6696 12316 6702 12368
rect 12636 12356 12664 12396
rect 13262 12384 13268 12396
rect 13320 12424 13326 12436
rect 14829 12427 14887 12433
rect 14829 12424 14841 12427
rect 13320 12396 14841 12424
rect 13320 12384 13326 12396
rect 14829 12393 14841 12396
rect 14875 12393 14887 12427
rect 14829 12387 14887 12393
rect 15286 12384 15292 12436
rect 15344 12424 15350 12436
rect 15381 12427 15439 12433
rect 15381 12424 15393 12427
rect 15344 12396 15393 12424
rect 15344 12384 15350 12396
rect 15381 12393 15393 12396
rect 15427 12393 15439 12427
rect 15381 12387 15439 12393
rect 17589 12427 17647 12433
rect 17589 12393 17601 12427
rect 17635 12424 17647 12427
rect 17770 12424 17776 12436
rect 17635 12396 17776 12424
rect 17635 12393 17647 12396
rect 17589 12387 17647 12393
rect 17770 12384 17776 12396
rect 17828 12384 17834 12436
rect 19518 12384 19524 12436
rect 19576 12424 19582 12436
rect 19705 12427 19763 12433
rect 19705 12424 19717 12427
rect 19576 12396 19717 12424
rect 19576 12384 19582 12396
rect 19705 12393 19717 12396
rect 19751 12393 19763 12427
rect 19705 12387 19763 12393
rect 19794 12384 19800 12436
rect 19852 12424 19858 12436
rect 20162 12424 20168 12436
rect 19852 12396 20168 12424
rect 19852 12384 19858 12396
rect 20162 12384 20168 12396
rect 20220 12384 20226 12436
rect 15102 12356 15108 12368
rect 10980 12328 12664 12356
rect 12728 12328 15108 12356
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12257 2375 12291
rect 2317 12251 2375 12257
rect 2501 12291 2559 12297
rect 2501 12257 2513 12291
rect 2547 12288 2559 12291
rect 2547 12260 2774 12288
rect 2547 12257 2559 12260
rect 2501 12251 2559 12257
rect 2746 12152 2774 12260
rect 2958 12248 2964 12300
rect 3016 12288 3022 12300
rect 3145 12291 3203 12297
rect 3145 12288 3157 12291
rect 3016 12260 3157 12288
rect 3016 12248 3022 12260
rect 3145 12257 3157 12260
rect 3191 12257 3203 12291
rect 3145 12251 3203 12257
rect 3329 12291 3387 12297
rect 3329 12257 3341 12291
rect 3375 12288 3387 12291
rect 4062 12288 4068 12300
rect 3375 12260 4068 12288
rect 3375 12257 3387 12260
rect 3329 12251 3387 12257
rect 2866 12180 2872 12232
rect 2924 12220 2930 12232
rect 3053 12223 3111 12229
rect 3053 12220 3065 12223
rect 2924 12192 3065 12220
rect 2924 12180 2930 12192
rect 3053 12189 3065 12192
rect 3099 12189 3111 12223
rect 3053 12183 3111 12189
rect 3344 12152 3372 12251
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 4890 12248 4896 12300
rect 4948 12288 4954 12300
rect 5261 12291 5319 12297
rect 5261 12288 5273 12291
rect 4948 12260 5273 12288
rect 4948 12248 4954 12260
rect 5261 12257 5273 12260
rect 5307 12257 5319 12291
rect 5442 12288 5448 12300
rect 5403 12260 5448 12288
rect 5261 12251 5319 12257
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 5626 12248 5632 12300
rect 5684 12288 5690 12300
rect 7282 12288 7288 12300
rect 5684 12260 6776 12288
rect 7243 12260 7288 12288
rect 5684 12248 5690 12260
rect 4614 12180 4620 12232
rect 4672 12220 4678 12232
rect 6748 12229 6776 12260
rect 7282 12248 7288 12260
rect 7340 12248 7346 12300
rect 9030 12288 9036 12300
rect 8312 12260 9036 12288
rect 6365 12223 6423 12229
rect 6365 12220 6377 12223
rect 4672 12192 6377 12220
rect 4672 12180 4678 12192
rect 6365 12189 6377 12192
rect 6411 12189 6423 12223
rect 6365 12183 6423 12189
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12189 6791 12223
rect 7098 12220 7104 12232
rect 7059 12192 7104 12220
rect 6733 12183 6791 12189
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 7837 12223 7895 12229
rect 7837 12189 7849 12223
rect 7883 12220 7895 12223
rect 7926 12220 7932 12232
rect 7883 12192 7932 12220
rect 7883 12189 7895 12192
rect 7837 12183 7895 12189
rect 7926 12180 7932 12192
rect 7984 12180 7990 12232
rect 8312 12229 8340 12260
rect 9030 12248 9036 12260
rect 9088 12248 9094 12300
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12189 8355 12223
rect 8297 12183 8355 12189
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12220 8631 12223
rect 8938 12220 8944 12232
rect 8619 12192 8944 12220
rect 8619 12189 8631 12192
rect 8573 12183 8631 12189
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 9122 12180 9128 12232
rect 9180 12220 9186 12232
rect 9306 12220 9312 12232
rect 9180 12192 9312 12220
rect 9180 12180 9186 12192
rect 9306 12180 9312 12192
rect 9364 12180 9370 12232
rect 9401 12223 9459 12229
rect 9401 12189 9413 12223
rect 9447 12220 9459 12223
rect 9858 12220 9864 12232
rect 9447 12192 9864 12220
rect 9447 12189 9459 12192
rect 9401 12183 9459 12189
rect 9858 12180 9864 12192
rect 9916 12220 9922 12232
rect 10778 12220 10784 12232
rect 9916 12192 10784 12220
rect 9916 12180 9922 12192
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 10879 12223 10937 12229
rect 10879 12189 10891 12223
rect 10925 12222 10937 12223
rect 10980 12222 11008 12328
rect 12161 12291 12219 12297
rect 12161 12288 12173 12291
rect 11624 12260 12173 12288
rect 11624 12232 11652 12260
rect 12161 12257 12173 12260
rect 12207 12288 12219 12291
rect 12728 12288 12756 12328
rect 15102 12316 15108 12328
rect 15160 12316 15166 12368
rect 17494 12316 17500 12368
rect 17552 12356 17558 12368
rect 17552 12328 18000 12356
rect 17552 12316 17558 12328
rect 14366 12288 14372 12300
rect 12207 12260 12756 12288
rect 13372 12260 14372 12288
rect 12207 12257 12219 12260
rect 12161 12251 12219 12257
rect 10925 12194 11008 12222
rect 11333 12223 11391 12229
rect 10925 12189 10937 12194
rect 10879 12183 10937 12189
rect 11333 12189 11345 12223
rect 11379 12220 11391 12223
rect 11606 12220 11612 12232
rect 11379 12192 11612 12220
rect 11379 12189 11391 12192
rect 11333 12183 11391 12189
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 11974 12220 11980 12232
rect 11935 12192 11980 12220
rect 11974 12180 11980 12192
rect 12032 12180 12038 12232
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 12124 12192 12169 12220
rect 12124 12180 12130 12192
rect 12250 12180 12256 12232
rect 12308 12220 12314 12232
rect 13081 12223 13139 12229
rect 12308 12192 12353 12220
rect 12308 12180 12314 12192
rect 13081 12189 13093 12223
rect 13127 12189 13139 12223
rect 13262 12220 13268 12232
rect 13223 12192 13268 12220
rect 13081 12183 13139 12189
rect 2746 12124 3372 12152
rect 4430 12112 4436 12164
rect 4488 12152 4494 12164
rect 5258 12152 5264 12164
rect 4488 12124 5264 12152
rect 4488 12112 4494 12124
rect 5258 12112 5264 12124
rect 5316 12112 5322 12164
rect 8481 12155 8539 12161
rect 8481 12121 8493 12155
rect 8527 12152 8539 12155
rect 9140 12152 9168 12180
rect 9674 12152 9680 12164
rect 8527 12124 9168 12152
rect 9635 12124 9680 12152
rect 8527 12121 8539 12124
rect 8481 12115 8539 12121
rect 9674 12112 9680 12124
rect 9732 12112 9738 12164
rect 9766 12112 9772 12164
rect 9824 12152 9830 12164
rect 9824 12124 9869 12152
rect 9824 12112 9830 12124
rect 10502 12112 10508 12164
rect 10560 12152 10566 12164
rect 10965 12155 11023 12161
rect 10965 12152 10977 12155
rect 10560 12124 10977 12152
rect 10560 12112 10566 12124
rect 10965 12121 10977 12124
rect 11011 12121 11023 12155
rect 10965 12115 11023 12121
rect 11057 12155 11115 12161
rect 11057 12121 11069 12155
rect 11103 12152 11115 12155
rect 12434 12152 12440 12164
rect 11103 12124 12440 12152
rect 11103 12121 11115 12124
rect 11057 12115 11115 12121
rect 12434 12112 12440 12124
rect 12492 12152 12498 12164
rect 13096 12152 13124 12183
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 12492 12124 13124 12152
rect 12492 12112 12498 12124
rect 1854 12084 1860 12096
rect 1815 12056 1860 12084
rect 1854 12044 1860 12056
rect 1912 12044 1918 12096
rect 2222 12084 2228 12096
rect 2183 12056 2228 12084
rect 2222 12044 2228 12056
rect 2280 12044 2286 12096
rect 3326 12084 3332 12096
rect 3287 12056 3332 12084
rect 3326 12044 3332 12056
rect 3384 12044 3390 12096
rect 4801 12087 4859 12093
rect 4801 12053 4813 12087
rect 4847 12084 4859 12087
rect 4890 12084 4896 12096
rect 4847 12056 4896 12084
rect 4847 12053 4859 12056
rect 4801 12047 4859 12053
rect 4890 12044 4896 12056
rect 4948 12044 4954 12096
rect 5169 12087 5227 12093
rect 5169 12053 5181 12087
rect 5215 12084 5227 12087
rect 6914 12084 6920 12096
rect 5215 12056 6920 12084
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 8386 12084 8392 12096
rect 8444 12093 8450 12096
rect 8353 12056 8392 12084
rect 8386 12044 8392 12056
rect 8444 12047 8453 12093
rect 10597 12087 10655 12093
rect 10597 12053 10609 12087
rect 10643 12084 10655 12087
rect 10686 12084 10692 12096
rect 10643 12056 10692 12084
rect 10643 12053 10655 12056
rect 10597 12047 10655 12053
rect 8444 12044 8450 12047
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 10778 12044 10784 12096
rect 10836 12084 10842 12096
rect 13372 12084 13400 12260
rect 14366 12248 14372 12260
rect 14424 12248 14430 12300
rect 16574 12288 16580 12300
rect 15396 12260 16344 12288
rect 16535 12260 16580 12288
rect 13630 12180 13636 12232
rect 13688 12220 13694 12232
rect 14274 12220 14280 12232
rect 13688 12192 14280 12220
rect 13688 12180 13694 12192
rect 14274 12180 14280 12192
rect 14332 12220 14338 12232
rect 14553 12223 14611 12229
rect 14553 12220 14565 12223
rect 14332 12192 14565 12220
rect 14332 12180 14338 12192
rect 14553 12189 14565 12192
rect 14599 12189 14611 12223
rect 14553 12183 14611 12189
rect 14642 12180 14648 12232
rect 14700 12220 14706 12232
rect 14918 12220 14924 12232
rect 14700 12192 14793 12220
rect 14879 12192 14924 12220
rect 14700 12180 14706 12192
rect 14918 12180 14924 12192
rect 14976 12180 14982 12232
rect 15010 12180 15016 12232
rect 15068 12220 15074 12232
rect 15396 12229 15424 12260
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 15068 12192 15393 12220
rect 15068 12180 15074 12192
rect 15381 12189 15393 12192
rect 15427 12189 15439 12223
rect 15565 12223 15623 12229
rect 15565 12220 15577 12223
rect 15381 12183 15439 12189
rect 15488 12192 15577 12220
rect 14458 12112 14464 12164
rect 14516 12152 14522 12164
rect 14660 12152 14688 12180
rect 14516 12124 14688 12152
rect 14516 12112 14522 12124
rect 15102 12112 15108 12164
rect 15160 12152 15166 12164
rect 15488 12152 15516 12192
rect 15565 12189 15577 12192
rect 15611 12220 15623 12223
rect 16206 12220 16212 12232
rect 15611 12192 16212 12220
rect 15611 12189 15623 12192
rect 15565 12183 15623 12189
rect 16206 12180 16212 12192
rect 16264 12180 16270 12232
rect 16316 12229 16344 12260
rect 16574 12248 16580 12260
rect 16632 12248 16638 12300
rect 16301 12223 16359 12229
rect 16301 12189 16313 12223
rect 16347 12220 16359 12223
rect 17586 12220 17592 12232
rect 16347 12192 17592 12220
rect 16347 12189 16359 12192
rect 16301 12183 16359 12189
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 17862 12229 17868 12232
rect 17845 12223 17868 12229
rect 17845 12189 17857 12223
rect 17845 12183 17868 12189
rect 17862 12180 17868 12183
rect 17920 12180 17926 12232
rect 17972 12229 18000 12328
rect 19610 12316 19616 12368
rect 19668 12356 19674 12368
rect 20073 12359 20131 12365
rect 20073 12356 20085 12359
rect 19668 12328 20085 12356
rect 19668 12316 19674 12328
rect 20073 12325 20085 12328
rect 20119 12325 20131 12359
rect 20073 12319 20131 12325
rect 18874 12248 18880 12300
rect 18932 12288 18938 12300
rect 19797 12291 19855 12297
rect 19797 12288 19809 12291
rect 18932 12260 19809 12288
rect 18932 12248 18938 12260
rect 19797 12257 19809 12260
rect 19843 12257 19855 12291
rect 19797 12251 19855 12257
rect 17954 12223 18012 12229
rect 17954 12189 17966 12223
rect 18000 12189 18012 12223
rect 17954 12183 18012 12189
rect 18046 12180 18052 12232
rect 18104 12220 18110 12232
rect 18233 12223 18291 12229
rect 18104 12192 18149 12220
rect 18104 12180 18110 12192
rect 18233 12189 18245 12223
rect 18279 12220 18291 12223
rect 18598 12220 18604 12232
rect 18279 12192 18604 12220
rect 18279 12189 18291 12192
rect 18233 12183 18291 12189
rect 15160 12124 15516 12152
rect 15160 12112 15166 12124
rect 16022 12112 16028 12164
rect 16080 12152 16086 12164
rect 16117 12155 16175 12161
rect 16117 12152 16129 12155
rect 16080 12124 16129 12152
rect 16080 12112 16086 12124
rect 16117 12121 16129 12124
rect 16163 12121 16175 12155
rect 16117 12115 16175 12121
rect 10836 12056 13400 12084
rect 13449 12087 13507 12093
rect 10836 12044 10842 12056
rect 13449 12053 13461 12087
rect 13495 12084 13507 12087
rect 15194 12084 15200 12096
rect 13495 12056 15200 12084
rect 13495 12053 13507 12056
rect 13449 12047 13507 12053
rect 15194 12044 15200 12056
rect 15252 12044 15258 12096
rect 16132 12084 16160 12115
rect 18248 12084 18276 12183
rect 18598 12180 18604 12192
rect 18656 12220 18662 12232
rect 19242 12220 19248 12232
rect 18656 12192 19248 12220
rect 18656 12180 18662 12192
rect 19242 12180 19248 12192
rect 19300 12180 19306 12232
rect 19705 12223 19763 12229
rect 19705 12189 19717 12223
rect 19751 12220 19763 12223
rect 19886 12220 19892 12232
rect 19751 12192 19892 12220
rect 19751 12189 19763 12192
rect 19705 12183 19763 12189
rect 19886 12180 19892 12192
rect 19944 12180 19950 12232
rect 16132 12056 18276 12084
rect 1104 11994 21043 12016
rect 1104 11942 5894 11994
rect 5946 11942 5958 11994
rect 6010 11942 6022 11994
rect 6074 11942 6086 11994
rect 6138 11942 6150 11994
rect 6202 11942 10839 11994
rect 10891 11942 10903 11994
rect 10955 11942 10967 11994
rect 11019 11942 11031 11994
rect 11083 11942 11095 11994
rect 11147 11942 15784 11994
rect 15836 11942 15848 11994
rect 15900 11942 15912 11994
rect 15964 11942 15976 11994
rect 16028 11942 16040 11994
rect 16092 11942 20729 11994
rect 20781 11942 20793 11994
rect 20845 11942 20857 11994
rect 20909 11942 20921 11994
rect 20973 11942 20985 11994
rect 21037 11942 21043 11994
rect 1104 11920 21043 11942
rect 2314 11840 2320 11892
rect 2372 11880 2378 11892
rect 2409 11883 2467 11889
rect 2409 11880 2421 11883
rect 2372 11852 2421 11880
rect 2372 11840 2378 11852
rect 2409 11849 2421 11852
rect 2455 11849 2467 11883
rect 2409 11843 2467 11849
rect 2774 11840 2780 11892
rect 2832 11880 2838 11892
rect 2869 11883 2927 11889
rect 2869 11880 2881 11883
rect 2832 11852 2881 11880
rect 2832 11840 2838 11852
rect 2869 11849 2881 11852
rect 2915 11849 2927 11883
rect 2869 11843 2927 11849
rect 7561 11883 7619 11889
rect 7561 11849 7573 11883
rect 7607 11880 7619 11883
rect 7650 11880 7656 11892
rect 7607 11852 7656 11880
rect 7607 11849 7619 11852
rect 7561 11843 7619 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 11238 11880 11244 11892
rect 9824 11852 11244 11880
rect 9824 11840 9830 11852
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 11974 11840 11980 11892
rect 12032 11880 12038 11892
rect 12161 11883 12219 11889
rect 12161 11880 12173 11883
rect 12032 11852 12173 11880
rect 12032 11840 12038 11852
rect 12161 11849 12173 11852
rect 12207 11849 12219 11883
rect 12342 11880 12348 11892
rect 12303 11852 12348 11880
rect 12161 11843 12219 11849
rect 4338 11772 4344 11824
rect 4396 11812 4402 11824
rect 4525 11815 4583 11821
rect 4525 11812 4537 11815
rect 4396 11784 4537 11812
rect 4396 11772 4402 11784
rect 4525 11781 4537 11784
rect 4571 11781 4583 11815
rect 4525 11775 4583 11781
rect 8754 11772 8760 11824
rect 8812 11812 8818 11824
rect 8849 11815 8907 11821
rect 8849 11812 8861 11815
rect 8812 11784 8861 11812
rect 8812 11772 8818 11784
rect 8849 11781 8861 11784
rect 8895 11781 8907 11815
rect 8849 11775 8907 11781
rect 9401 11815 9459 11821
rect 9401 11781 9413 11815
rect 9447 11812 9459 11815
rect 9950 11812 9956 11824
rect 9447 11784 9956 11812
rect 9447 11781 9459 11784
rect 9401 11775 9459 11781
rect 9950 11772 9956 11784
rect 10008 11772 10014 11824
rect 10594 11772 10600 11824
rect 10652 11812 10658 11824
rect 12176 11812 12204 11843
rect 12342 11840 12348 11852
rect 12400 11840 12406 11892
rect 13446 11840 13452 11892
rect 13504 11880 13510 11892
rect 13541 11883 13599 11889
rect 13541 11880 13553 11883
rect 13504 11852 13553 11880
rect 13504 11840 13510 11852
rect 13541 11849 13553 11852
rect 13587 11849 13599 11883
rect 13541 11843 13599 11849
rect 13630 11840 13636 11892
rect 13688 11880 13694 11892
rect 16666 11880 16672 11892
rect 13688 11852 16672 11880
rect 13688 11840 13694 11852
rect 10652 11784 10824 11812
rect 12176 11784 12434 11812
rect 10652 11772 10658 11784
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11744 2283 11747
rect 2774 11744 2780 11756
rect 2271 11716 2780 11744
rect 2271 11713 2283 11716
rect 2225 11707 2283 11713
rect 2774 11704 2780 11716
rect 2832 11704 2838 11756
rect 3234 11744 3240 11756
rect 3147 11716 3240 11744
rect 3234 11704 3240 11716
rect 3292 11744 3298 11756
rect 3878 11744 3884 11756
rect 3292 11716 3884 11744
rect 3292 11704 3298 11716
rect 3878 11704 3884 11716
rect 3936 11704 3942 11756
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11713 4307 11747
rect 4430 11744 4436 11756
rect 4391 11716 4436 11744
rect 4249 11707 4307 11713
rect 2041 11679 2099 11685
rect 2041 11645 2053 11679
rect 2087 11676 2099 11679
rect 2866 11676 2872 11688
rect 2087 11648 2872 11676
rect 2087 11645 2099 11648
rect 2041 11639 2099 11645
rect 2866 11636 2872 11648
rect 2924 11636 2930 11688
rect 3329 11679 3387 11685
rect 3329 11645 3341 11679
rect 3375 11645 3387 11679
rect 4264 11676 4292 11707
rect 4430 11704 4436 11716
rect 4488 11704 4494 11756
rect 4614 11744 4620 11756
rect 4575 11716 4620 11744
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 5442 11744 5448 11756
rect 5355 11716 5448 11744
rect 5442 11704 5448 11716
rect 5500 11744 5506 11756
rect 5500 11716 5948 11744
rect 5500 11704 5506 11716
rect 5261 11679 5319 11685
rect 5261 11676 5273 11679
rect 4264 11648 5273 11676
rect 3329 11639 3387 11645
rect 5261 11645 5273 11648
rect 5307 11645 5319 11679
rect 5261 11639 5319 11645
rect 5721 11679 5779 11685
rect 5721 11645 5733 11679
rect 5767 11676 5779 11679
rect 5810 11676 5816 11688
rect 5767 11648 5816 11676
rect 5767 11645 5779 11648
rect 5721 11639 5779 11645
rect 3344 11608 3372 11639
rect 5810 11636 5816 11648
rect 5868 11636 5874 11688
rect 5534 11608 5540 11620
rect 3344 11580 5540 11608
rect 5534 11568 5540 11580
rect 5592 11608 5598 11620
rect 5629 11611 5687 11617
rect 5629 11608 5641 11611
rect 5592 11580 5641 11608
rect 5592 11568 5598 11580
rect 5629 11577 5641 11580
rect 5675 11577 5687 11611
rect 5920 11608 5948 11716
rect 6914 11704 6920 11756
rect 6972 11744 6978 11756
rect 7469 11747 7527 11753
rect 7469 11744 7481 11747
rect 6972 11716 7481 11744
rect 6972 11704 6978 11716
rect 7469 11713 7481 11716
rect 7515 11713 7527 11747
rect 7469 11707 7527 11713
rect 8386 11704 8392 11756
rect 8444 11744 8450 11756
rect 9033 11747 9091 11753
rect 9033 11744 9045 11747
rect 8444 11716 9045 11744
rect 8444 11704 8450 11716
rect 9033 11713 9045 11716
rect 9079 11713 9091 11747
rect 10502 11744 10508 11756
rect 10463 11716 10508 11744
rect 9033 11707 9091 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10686 11744 10692 11756
rect 10647 11716 10692 11744
rect 10686 11704 10692 11716
rect 10744 11704 10750 11756
rect 10796 11753 10824 11784
rect 10781 11747 10839 11753
rect 10781 11713 10793 11747
rect 10827 11713 10839 11747
rect 10781 11707 10839 11713
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 11977 11747 12035 11753
rect 11977 11744 11989 11747
rect 11664 11716 11989 11744
rect 11664 11704 11670 11716
rect 11977 11713 11989 11716
rect 12023 11713 12035 11747
rect 11977 11707 12035 11713
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 12124 11716 12217 11744
rect 12124 11704 12130 11716
rect 7282 11636 7288 11688
rect 7340 11676 7346 11688
rect 7653 11679 7711 11685
rect 7653 11676 7665 11679
rect 7340 11648 7665 11676
rect 7340 11636 7346 11648
rect 7653 11645 7665 11648
rect 7699 11645 7711 11679
rect 7653 11639 7711 11645
rect 10597 11679 10655 11685
rect 10597 11645 10609 11679
rect 10643 11676 10655 11679
rect 11698 11676 11704 11688
rect 10643 11648 11704 11676
rect 10643 11645 10655 11648
rect 10597 11639 10655 11645
rect 11698 11636 11704 11648
rect 11756 11636 11762 11688
rect 7558 11608 7564 11620
rect 5920 11580 7564 11608
rect 5629 11571 5687 11577
rect 7558 11568 7564 11580
rect 7616 11568 7622 11620
rect 11514 11568 11520 11620
rect 11572 11608 11578 11620
rect 11793 11611 11851 11617
rect 11793 11608 11805 11611
rect 11572 11580 11805 11608
rect 11572 11568 11578 11580
rect 11793 11577 11805 11580
rect 11839 11577 11851 11611
rect 12084 11608 12112 11704
rect 12406 11676 12434 11784
rect 13170 11772 13176 11824
rect 13228 11812 13234 11824
rect 15948 11821 15976 11852
rect 16666 11840 16672 11852
rect 16724 11840 16730 11892
rect 19242 11880 19248 11892
rect 19203 11852 19248 11880
rect 19242 11840 19248 11852
rect 19300 11840 19306 11892
rect 19978 11840 19984 11892
rect 20036 11880 20042 11892
rect 20073 11883 20131 11889
rect 20073 11880 20085 11883
rect 20036 11852 20085 11880
rect 20036 11840 20042 11852
rect 20073 11849 20085 11852
rect 20119 11849 20131 11883
rect 20073 11843 20131 11849
rect 14185 11815 14243 11821
rect 14185 11812 14197 11815
rect 13228 11784 14197 11812
rect 13228 11772 13234 11784
rect 12986 11704 12992 11756
rect 13044 11744 13050 11756
rect 13357 11747 13415 11753
rect 13357 11744 13369 11747
rect 13044 11716 13369 11744
rect 13044 11704 13050 11716
rect 13357 11713 13369 11716
rect 13403 11744 13415 11747
rect 13538 11744 13544 11756
rect 13403 11716 13544 11744
rect 13403 11713 13415 11716
rect 13357 11707 13415 11713
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 13648 11753 13676 11784
rect 14185 11781 14197 11784
rect 14231 11781 14243 11815
rect 14185 11775 14243 11781
rect 15933 11815 15991 11821
rect 15933 11781 15945 11815
rect 15979 11781 15991 11815
rect 16206 11812 16212 11824
rect 15933 11775 15991 11781
rect 16040 11784 16212 11812
rect 13633 11747 13691 11753
rect 13633 11713 13645 11747
rect 13679 11713 13691 11747
rect 14090 11744 14096 11756
rect 14051 11716 14096 11744
rect 13633 11707 13691 11713
rect 14090 11704 14096 11716
rect 14148 11704 14154 11756
rect 14274 11704 14280 11756
rect 14332 11744 14338 11756
rect 15013 11747 15071 11753
rect 14332 11716 14425 11744
rect 14332 11704 14338 11716
rect 15013 11713 15025 11747
rect 15059 11744 15071 11747
rect 15102 11744 15108 11756
rect 15059 11716 15108 11744
rect 15059 11713 15071 11716
rect 15013 11707 15071 11713
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 15197 11747 15255 11753
rect 15197 11713 15209 11747
rect 15243 11744 15255 11747
rect 15286 11744 15292 11756
rect 15243 11716 15292 11744
rect 15243 11713 15255 11716
rect 15197 11707 15255 11713
rect 15286 11704 15292 11716
rect 15344 11704 15350 11756
rect 15654 11744 15660 11756
rect 15615 11716 15660 11744
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 15746 11704 15752 11756
rect 15804 11744 15810 11756
rect 16040 11753 16068 11784
rect 16206 11772 16212 11784
rect 16264 11812 16270 11824
rect 17034 11812 17040 11824
rect 16264 11784 17040 11812
rect 16264 11772 16270 11784
rect 17034 11772 17040 11784
rect 17092 11772 17098 11824
rect 17862 11772 17868 11824
rect 17920 11812 17926 11824
rect 17920 11784 19288 11812
rect 17920 11772 17926 11784
rect 16025 11747 16083 11753
rect 15804 11716 15849 11744
rect 15804 11704 15810 11716
rect 16025 11713 16037 11747
rect 16071 11713 16083 11747
rect 16025 11707 16083 11713
rect 16122 11747 16180 11753
rect 16122 11713 16134 11747
rect 16168 11744 16180 11747
rect 16390 11744 16396 11756
rect 16168 11716 16396 11744
rect 16168 11713 16180 11716
rect 16122 11707 16180 11713
rect 14182 11676 14188 11688
rect 12406 11648 14188 11676
rect 14182 11636 14188 11648
rect 14240 11636 14246 11688
rect 12342 11608 12348 11620
rect 12084 11580 12348 11608
rect 11793 11571 11851 11577
rect 3234 11500 3240 11552
rect 3292 11540 3298 11552
rect 3513 11543 3571 11549
rect 3513 11540 3525 11543
rect 3292 11512 3525 11540
rect 3292 11500 3298 11512
rect 3513 11509 3525 11512
rect 3559 11509 3571 11543
rect 3513 11503 3571 11509
rect 3786 11500 3792 11552
rect 3844 11540 3850 11552
rect 4801 11543 4859 11549
rect 4801 11540 4813 11543
rect 3844 11512 4813 11540
rect 3844 11500 3850 11512
rect 4801 11509 4813 11512
rect 4847 11509 4859 11543
rect 4801 11503 4859 11509
rect 7101 11543 7159 11549
rect 7101 11509 7113 11543
rect 7147 11540 7159 11543
rect 7190 11540 7196 11552
rect 7147 11512 7196 11540
rect 7147 11509 7159 11512
rect 7101 11503 7159 11509
rect 7190 11500 7196 11512
rect 7248 11500 7254 11552
rect 10318 11540 10324 11552
rect 10279 11512 10324 11540
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 11808 11540 11836 11571
rect 12342 11568 12348 11580
rect 12400 11568 12406 11620
rect 14292 11608 14320 11704
rect 15120 11676 15148 11704
rect 16132 11676 16160 11707
rect 16390 11704 16396 11716
rect 16448 11704 16454 11756
rect 17494 11744 17500 11756
rect 17455 11716 17500 11744
rect 17494 11704 17500 11716
rect 17552 11704 17558 11756
rect 18601 11747 18659 11753
rect 18601 11713 18613 11747
rect 18647 11744 18659 11747
rect 19150 11744 19156 11756
rect 18647 11716 19156 11744
rect 18647 11713 18659 11716
rect 18601 11707 18659 11713
rect 19150 11704 19156 11716
rect 19208 11704 19214 11756
rect 19260 11744 19288 11784
rect 19426 11772 19432 11824
rect 19484 11812 19490 11824
rect 19797 11815 19855 11821
rect 19797 11812 19809 11815
rect 19484 11784 19809 11812
rect 19484 11772 19490 11784
rect 19797 11781 19809 11784
rect 19843 11781 19855 11815
rect 19797 11775 19855 11781
rect 19702 11744 19708 11756
rect 19260 11716 19708 11744
rect 19702 11704 19708 11716
rect 19760 11744 19766 11756
rect 19981 11747 20039 11753
rect 19981 11744 19993 11747
rect 19760 11716 19993 11744
rect 19760 11704 19766 11716
rect 19981 11713 19993 11716
rect 20027 11713 20039 11747
rect 19981 11707 20039 11713
rect 17310 11676 17316 11688
rect 15120 11648 16160 11676
rect 17271 11648 17316 11676
rect 17310 11636 17316 11648
rect 17368 11636 17374 11688
rect 18874 11636 18880 11688
rect 18932 11676 18938 11688
rect 18969 11679 19027 11685
rect 18969 11676 18981 11679
rect 18932 11648 18981 11676
rect 18932 11636 18938 11648
rect 18969 11645 18981 11648
rect 19015 11645 19027 11679
rect 18969 11639 19027 11645
rect 18766 11611 18824 11617
rect 14292 11580 16436 11608
rect 16408 11552 16436 11580
rect 18766 11577 18778 11611
rect 18812 11608 18824 11611
rect 19242 11608 19248 11620
rect 18812 11580 19248 11608
rect 18812 11577 18824 11580
rect 18766 11571 18824 11577
rect 19242 11568 19248 11580
rect 19300 11568 19306 11620
rect 12250 11540 12256 11552
rect 11808 11512 12256 11540
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 13357 11543 13415 11549
rect 13357 11509 13369 11543
rect 13403 11540 13415 11543
rect 13814 11540 13820 11552
rect 13403 11512 13820 11540
rect 13403 11509 13415 11512
rect 13357 11503 13415 11509
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 14090 11500 14096 11552
rect 14148 11540 14154 11552
rect 14274 11540 14280 11552
rect 14148 11512 14280 11540
rect 14148 11500 14154 11512
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 15013 11543 15071 11549
rect 15013 11509 15025 11543
rect 15059 11540 15071 11543
rect 15562 11540 15568 11552
rect 15059 11512 15568 11540
rect 15059 11509 15071 11512
rect 15013 11503 15071 11509
rect 15562 11500 15568 11512
rect 15620 11500 15626 11552
rect 16298 11540 16304 11552
rect 16259 11512 16304 11540
rect 16298 11500 16304 11512
rect 16356 11500 16362 11552
rect 16390 11500 16396 11552
rect 16448 11540 16454 11552
rect 17681 11543 17739 11549
rect 17681 11540 17693 11543
rect 16448 11512 17693 11540
rect 16448 11500 16454 11512
rect 17681 11509 17693 11512
rect 17727 11509 17739 11543
rect 17681 11503 17739 11509
rect 18877 11543 18935 11549
rect 18877 11509 18889 11543
rect 18923 11540 18935 11543
rect 19886 11540 19892 11552
rect 18923 11512 19892 11540
rect 18923 11509 18935 11512
rect 18877 11503 18935 11509
rect 19886 11500 19892 11512
rect 19944 11500 19950 11552
rect 1104 11450 20884 11472
rect 1104 11398 3422 11450
rect 3474 11398 3486 11450
rect 3538 11398 3550 11450
rect 3602 11398 3614 11450
rect 3666 11398 3678 11450
rect 3730 11398 8367 11450
rect 8419 11398 8431 11450
rect 8483 11398 8495 11450
rect 8547 11398 8559 11450
rect 8611 11398 8623 11450
rect 8675 11398 13312 11450
rect 13364 11398 13376 11450
rect 13428 11398 13440 11450
rect 13492 11398 13504 11450
rect 13556 11398 13568 11450
rect 13620 11398 18257 11450
rect 18309 11398 18321 11450
rect 18373 11398 18385 11450
rect 18437 11398 18449 11450
rect 18501 11398 18513 11450
rect 18565 11398 20884 11450
rect 1104 11376 20884 11398
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 14645 11339 14703 11345
rect 12492 11308 12537 11336
rect 12492 11296 12498 11308
rect 14645 11305 14657 11339
rect 14691 11336 14703 11339
rect 15010 11336 15016 11348
rect 14691 11308 15016 11336
rect 14691 11305 14703 11308
rect 14645 11299 14703 11305
rect 15010 11296 15016 11308
rect 15068 11296 15074 11348
rect 15746 11296 15752 11348
rect 15804 11336 15810 11348
rect 16117 11339 16175 11345
rect 16117 11336 16129 11339
rect 15804 11308 16129 11336
rect 15804 11296 15810 11308
rect 16117 11305 16129 11308
rect 16163 11305 16175 11339
rect 16117 11299 16175 11305
rect 1857 11271 1915 11277
rect 1857 11237 1869 11271
rect 1903 11268 1915 11271
rect 1946 11268 1952 11280
rect 1903 11240 1952 11268
rect 1903 11237 1915 11240
rect 1857 11231 1915 11237
rect 1946 11228 1952 11240
rect 2004 11228 2010 11280
rect 6733 11271 6791 11277
rect 6733 11237 6745 11271
rect 6779 11268 6791 11271
rect 7098 11268 7104 11280
rect 6779 11240 7104 11268
rect 6779 11237 6791 11240
rect 6733 11231 6791 11237
rect 7098 11228 7104 11240
rect 7156 11228 7162 11280
rect 13078 11228 13084 11280
rect 13136 11268 13142 11280
rect 14277 11271 14335 11277
rect 14277 11268 14289 11271
rect 13136 11240 14289 11268
rect 13136 11228 13142 11240
rect 14277 11237 14289 11240
rect 14323 11237 14335 11271
rect 14277 11231 14335 11237
rect 14458 11228 14464 11280
rect 14516 11268 14522 11280
rect 16025 11271 16083 11277
rect 16025 11268 16037 11271
rect 14516 11240 16037 11268
rect 14516 11228 14522 11240
rect 16025 11237 16037 11240
rect 16071 11237 16083 11271
rect 18046 11268 18052 11280
rect 16025 11231 16083 11237
rect 16132 11240 18052 11268
rect 3326 11200 3332 11212
rect 1872 11172 3332 11200
rect 1872 11141 1900 11172
rect 3326 11160 3332 11172
rect 3384 11160 3390 11212
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 4157 11203 4215 11209
rect 4157 11200 4169 11203
rect 3936 11172 4169 11200
rect 3936 11160 3942 11172
rect 4157 11169 4169 11172
rect 4203 11169 4215 11203
rect 7190 11200 7196 11212
rect 7151 11172 7196 11200
rect 4157 11163 4215 11169
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7377 11203 7435 11209
rect 7377 11169 7389 11203
rect 7423 11200 7435 11203
rect 7558 11200 7564 11212
rect 7423 11172 7564 11200
rect 7423 11169 7435 11172
rect 7377 11163 7435 11169
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 14182 11160 14188 11212
rect 14240 11200 14246 11212
rect 16132 11200 16160 11240
rect 18046 11228 18052 11240
rect 18104 11228 18110 11280
rect 18874 11228 18880 11280
rect 18932 11268 18938 11280
rect 18932 11240 19748 11268
rect 18932 11228 18938 11240
rect 14240 11172 16160 11200
rect 16209 11203 16267 11209
rect 14240 11160 14246 11172
rect 16209 11169 16221 11203
rect 16255 11200 16267 11203
rect 17218 11200 17224 11212
rect 16255 11172 17224 11200
rect 16255 11169 16267 11172
rect 16209 11163 16267 11169
rect 17218 11160 17224 11172
rect 17276 11160 17282 11212
rect 19242 11160 19248 11212
rect 19300 11200 19306 11212
rect 19521 11203 19579 11209
rect 19521 11200 19533 11203
rect 19300 11172 19533 11200
rect 19300 11160 19306 11172
rect 19521 11169 19533 11172
rect 19567 11169 19579 11203
rect 19521 11163 19579 11169
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11101 1915 11135
rect 1857 11095 1915 11101
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11132 2191 11135
rect 2958 11132 2964 11144
rect 2179 11104 2964 11132
rect 2179 11101 2191 11104
rect 2133 11095 2191 11101
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 3970 11132 3976 11144
rect 3931 11104 3976 11132
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 12342 11132 12348 11144
rect 12303 11104 12348 11132
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11132 13599 11135
rect 14458 11132 14464 11144
rect 13587 11104 14464 11132
rect 13587 11101 13599 11104
rect 13541 11095 13599 11101
rect 14458 11092 14464 11104
rect 14516 11092 14522 11144
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11132 15991 11135
rect 16390 11132 16396 11144
rect 15979 11104 16396 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 17586 11132 17592 11144
rect 17499 11104 17592 11132
rect 17586 11092 17592 11104
rect 17644 11092 17650 11144
rect 19150 11092 19156 11144
rect 19208 11132 19214 11144
rect 19720 11141 19748 11240
rect 20162 11200 20168 11212
rect 20123 11172 20168 11200
rect 20162 11160 20168 11172
rect 20220 11160 20226 11212
rect 19429 11135 19487 11141
rect 19429 11132 19441 11135
rect 19208 11104 19441 11132
rect 19208 11092 19214 11104
rect 19429 11101 19441 11104
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 19705 11135 19763 11141
rect 19705 11101 19717 11135
rect 19751 11101 19763 11135
rect 19705 11095 19763 11101
rect 2041 11067 2099 11073
rect 2041 11033 2053 11067
rect 2087 11064 2099 11067
rect 2866 11064 2872 11076
rect 2087 11036 2872 11064
rect 2087 11033 2099 11036
rect 2041 11027 2099 11033
rect 2866 11024 2872 11036
rect 2924 11024 2930 11076
rect 7101 11067 7159 11073
rect 7101 11033 7113 11067
rect 7147 11064 7159 11067
rect 7190 11064 7196 11076
rect 7147 11036 7196 11064
rect 7147 11033 7159 11036
rect 7101 11027 7159 11033
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 11330 11024 11336 11076
rect 11388 11064 11394 11076
rect 13633 11067 13691 11073
rect 13633 11064 13645 11067
rect 11388 11036 13645 11064
rect 11388 11024 11394 11036
rect 13633 11033 13645 11036
rect 13679 11064 13691 11067
rect 14645 11067 14703 11073
rect 14645 11064 14657 11067
rect 13679 11036 14657 11064
rect 13679 11033 13691 11036
rect 13633 11027 13691 11033
rect 14645 11033 14657 11036
rect 14691 11033 14703 11067
rect 17604 11064 17632 11092
rect 19978 11064 19984 11076
rect 17604 11036 19984 11064
rect 14645 11027 14703 11033
rect 19978 11024 19984 11036
rect 20036 11024 20042 11076
rect 2774 10956 2780 11008
rect 2832 10996 2838 11008
rect 2958 10996 2964 11008
rect 2832 10968 2964 10996
rect 2832 10956 2838 10968
rect 2958 10956 2964 10968
rect 3016 10956 3022 11008
rect 13998 10956 14004 11008
rect 14056 10996 14062 11008
rect 14829 10999 14887 11005
rect 14829 10996 14841 10999
rect 14056 10968 14841 10996
rect 14056 10956 14062 10968
rect 14829 10965 14841 10968
rect 14875 10965 14887 10999
rect 14829 10959 14887 10965
rect 16850 10956 16856 11008
rect 16908 10996 16914 11008
rect 17681 10999 17739 11005
rect 17681 10996 17693 10999
rect 16908 10968 17693 10996
rect 16908 10956 16914 10968
rect 17681 10965 17693 10968
rect 17727 10996 17739 10999
rect 17770 10996 17776 11008
rect 17727 10968 17776 10996
rect 17727 10965 17739 10968
rect 17681 10959 17739 10965
rect 17770 10956 17776 10968
rect 17828 10956 17834 11008
rect 1104 10906 21043 10928
rect 1104 10854 5894 10906
rect 5946 10854 5958 10906
rect 6010 10854 6022 10906
rect 6074 10854 6086 10906
rect 6138 10854 6150 10906
rect 6202 10854 10839 10906
rect 10891 10854 10903 10906
rect 10955 10854 10967 10906
rect 11019 10854 11031 10906
rect 11083 10854 11095 10906
rect 11147 10854 15784 10906
rect 15836 10854 15848 10906
rect 15900 10854 15912 10906
rect 15964 10854 15976 10906
rect 16028 10854 16040 10906
rect 16092 10854 20729 10906
rect 20781 10854 20793 10906
rect 20845 10854 20857 10906
rect 20909 10854 20921 10906
rect 20973 10854 20985 10906
rect 21037 10854 21043 10906
rect 1104 10832 21043 10854
rect 6822 10752 6828 10804
rect 6880 10792 6886 10804
rect 15470 10792 15476 10804
rect 6880 10764 15476 10792
rect 6880 10752 6886 10764
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 19150 10792 19156 10804
rect 18432 10764 19156 10792
rect 1670 10724 1676 10736
rect 1631 10696 1676 10724
rect 1670 10684 1676 10696
rect 1728 10684 1734 10736
rect 1857 10727 1915 10733
rect 1857 10693 1869 10727
rect 1903 10724 1915 10727
rect 3970 10724 3976 10736
rect 1903 10696 3976 10724
rect 1903 10693 1915 10696
rect 1857 10687 1915 10693
rect 3970 10684 3976 10696
rect 4028 10684 4034 10736
rect 10036 10727 10094 10733
rect 10036 10693 10048 10727
rect 10082 10724 10094 10727
rect 10318 10724 10324 10736
rect 10082 10696 10324 10724
rect 10082 10693 10094 10696
rect 10036 10687 10094 10693
rect 10318 10684 10324 10696
rect 10376 10684 10382 10736
rect 18432 10733 18460 10764
rect 19150 10752 19156 10764
rect 19208 10792 19214 10804
rect 19613 10795 19671 10801
rect 19613 10792 19625 10795
rect 19208 10764 19625 10792
rect 19208 10752 19214 10764
rect 19613 10761 19625 10764
rect 19659 10761 19671 10795
rect 19613 10755 19671 10761
rect 18417 10727 18475 10733
rect 18417 10693 18429 10727
rect 18463 10693 18475 10727
rect 19426 10724 19432 10736
rect 18417 10687 18475 10693
rect 18524 10696 19432 10724
rect 8012 10659 8070 10665
rect 8012 10625 8024 10659
rect 8058 10656 8070 10659
rect 13814 10656 13820 10668
rect 8058 10628 11284 10656
rect 13775 10628 13820 10656
rect 8058 10625 8070 10628
rect 8012 10619 8070 10625
rect 11256 10600 11284 10628
rect 13814 10616 13820 10628
rect 13872 10616 13878 10668
rect 14918 10616 14924 10668
rect 14976 10656 14982 10668
rect 16850 10656 16856 10668
rect 14976 10628 16856 10656
rect 14976 10616 14982 10628
rect 16850 10616 16856 10628
rect 16908 10616 16914 10668
rect 17034 10656 17040 10668
rect 16995 10628 17040 10656
rect 17034 10616 17040 10628
rect 17092 10656 17098 10668
rect 18524 10656 18552 10696
rect 19426 10684 19432 10696
rect 19484 10724 19490 10736
rect 19794 10724 19800 10736
rect 19484 10696 19800 10724
rect 19484 10684 19490 10696
rect 19794 10684 19800 10696
rect 19852 10724 19858 10736
rect 19852 10696 20024 10724
rect 19852 10684 19858 10696
rect 17092 10628 18552 10656
rect 18601 10659 18659 10665
rect 17092 10616 17098 10628
rect 18601 10625 18613 10659
rect 18647 10656 18659 10659
rect 19242 10656 19248 10668
rect 18647 10628 19248 10656
rect 18647 10625 18659 10628
rect 18601 10619 18659 10625
rect 19242 10616 19248 10628
rect 19300 10616 19306 10668
rect 19610 10656 19616 10668
rect 19571 10628 19616 10656
rect 19610 10616 19616 10628
rect 19668 10616 19674 10668
rect 19996 10665 20024 10696
rect 19981 10659 20039 10665
rect 19981 10625 19993 10659
rect 20027 10625 20039 10659
rect 19981 10619 20039 10625
rect 7006 10548 7012 10600
rect 7064 10588 7070 10600
rect 7745 10591 7803 10597
rect 7745 10588 7757 10591
rect 7064 10560 7757 10588
rect 7064 10548 7070 10560
rect 7745 10557 7757 10560
rect 7791 10557 7803 10591
rect 9766 10588 9772 10600
rect 9727 10560 9772 10588
rect 7745 10551 7803 10557
rect 9766 10548 9772 10560
rect 9824 10548 9830 10600
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 13170 10588 13176 10600
rect 11296 10560 13176 10588
rect 11296 10548 11302 10560
rect 13170 10548 13176 10560
rect 13228 10588 13234 10600
rect 13909 10591 13967 10597
rect 13909 10588 13921 10591
rect 13228 10560 13921 10588
rect 13228 10548 13234 10560
rect 13909 10557 13921 10560
rect 13955 10557 13967 10591
rect 13909 10551 13967 10557
rect 18046 10548 18052 10600
rect 18104 10588 18110 10600
rect 19429 10591 19487 10597
rect 19429 10588 19441 10591
rect 18104 10560 19441 10588
rect 18104 10548 18110 10560
rect 19429 10557 19441 10560
rect 19475 10557 19487 10591
rect 19429 10551 19487 10557
rect 9122 10520 9128 10532
rect 9083 10492 9128 10520
rect 9122 10480 9128 10492
rect 9180 10480 9186 10532
rect 14274 10480 14280 10532
rect 14332 10520 14338 10532
rect 15286 10520 15292 10532
rect 14332 10492 15292 10520
rect 14332 10480 14338 10492
rect 15286 10480 15292 10492
rect 15344 10480 15350 10532
rect 11149 10455 11207 10461
rect 11149 10421 11161 10455
rect 11195 10452 11207 10455
rect 13722 10452 13728 10464
rect 11195 10424 13728 10452
rect 11195 10421 11207 10424
rect 11149 10415 11207 10421
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 13998 10452 14004 10464
rect 13959 10424 14004 10452
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 14185 10455 14243 10461
rect 14185 10421 14197 10455
rect 14231 10452 14243 10455
rect 14550 10452 14556 10464
rect 14231 10424 14556 10452
rect 14231 10421 14243 10424
rect 14185 10415 14243 10421
rect 14550 10412 14556 10424
rect 14608 10412 14614 10464
rect 16945 10455 17003 10461
rect 16945 10421 16957 10455
rect 16991 10452 17003 10455
rect 17126 10452 17132 10464
rect 16991 10424 17132 10452
rect 16991 10421 17003 10424
rect 16945 10415 17003 10421
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 18690 10452 18696 10464
rect 18651 10424 18696 10452
rect 18690 10412 18696 10424
rect 18748 10412 18754 10464
rect 1104 10362 20884 10384
rect 1104 10310 3422 10362
rect 3474 10310 3486 10362
rect 3538 10310 3550 10362
rect 3602 10310 3614 10362
rect 3666 10310 3678 10362
rect 3730 10310 8367 10362
rect 8419 10310 8431 10362
rect 8483 10310 8495 10362
rect 8547 10310 8559 10362
rect 8611 10310 8623 10362
rect 8675 10310 13312 10362
rect 13364 10310 13376 10362
rect 13428 10310 13440 10362
rect 13492 10310 13504 10362
rect 13556 10310 13568 10362
rect 13620 10310 18257 10362
rect 18309 10310 18321 10362
rect 18373 10310 18385 10362
rect 18437 10310 18449 10362
rect 18501 10310 18513 10362
rect 18565 10310 20884 10362
rect 1104 10288 20884 10310
rect 2222 10208 2228 10260
rect 2280 10248 2286 10260
rect 2961 10251 3019 10257
rect 2961 10248 2973 10251
rect 2280 10220 2973 10248
rect 2280 10208 2286 10220
rect 2961 10217 2973 10220
rect 3007 10217 3019 10251
rect 2961 10211 3019 10217
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 8389 10251 8447 10257
rect 8389 10248 8401 10251
rect 7248 10220 8401 10248
rect 7248 10208 7254 10220
rect 8389 10217 8401 10220
rect 8435 10217 8447 10251
rect 11606 10248 11612 10260
rect 11567 10220 11612 10248
rect 8389 10211 8447 10217
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 14918 10248 14924 10260
rect 12820 10220 14924 10248
rect 10321 10115 10379 10121
rect 10321 10081 10333 10115
rect 10367 10112 10379 10115
rect 11330 10112 11336 10124
rect 10367 10084 11336 10112
rect 10367 10081 10379 10084
rect 10321 10075 10379 10081
rect 11330 10072 11336 10084
rect 11388 10072 11394 10124
rect 1578 10044 1584 10056
rect 1539 10016 1584 10044
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 1854 10053 1860 10056
rect 1848 10044 1860 10053
rect 1815 10016 1860 10044
rect 1848 10007 1860 10016
rect 1854 10004 1860 10007
rect 1912 10004 1918 10056
rect 3878 10004 3884 10056
rect 3936 10044 3942 10056
rect 5077 10047 5135 10053
rect 5077 10044 5089 10047
rect 3936 10016 5089 10044
rect 3936 10004 3942 10016
rect 5077 10013 5089 10016
rect 5123 10013 5135 10047
rect 5077 10007 5135 10013
rect 5344 10047 5402 10053
rect 5344 10013 5356 10047
rect 5390 10044 5402 10047
rect 6822 10044 6828 10056
rect 5390 10016 6828 10044
rect 5390 10013 5402 10016
rect 5344 10007 5402 10013
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 7006 10044 7012 10056
rect 6967 10016 7012 10044
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 7098 10004 7104 10056
rect 7156 10044 7162 10056
rect 7265 10047 7323 10053
rect 7265 10044 7277 10047
rect 7156 10016 7277 10044
rect 7156 10004 7162 10016
rect 7265 10013 7277 10016
rect 7311 10013 7323 10047
rect 7265 10007 7323 10013
rect 9766 10004 9772 10056
rect 9824 10044 9830 10056
rect 10045 10047 10103 10053
rect 10045 10044 10057 10047
rect 9824 10016 10057 10044
rect 9824 10004 9830 10016
rect 10045 10013 10057 10016
rect 10091 10013 10103 10047
rect 10045 10007 10103 10013
rect 11422 10004 11428 10056
rect 11480 10044 11486 10056
rect 12820 10053 12848 10220
rect 14918 10208 14924 10220
rect 14976 10208 14982 10260
rect 15286 10208 15292 10260
rect 15344 10248 15350 10260
rect 16669 10251 16727 10257
rect 16669 10248 16681 10251
rect 15344 10220 16681 10248
rect 15344 10208 15350 10220
rect 16669 10217 16681 10220
rect 16715 10248 16727 10251
rect 18690 10248 18696 10260
rect 16715 10220 18696 10248
rect 16715 10217 16727 10220
rect 16669 10211 16727 10217
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 18874 10208 18880 10260
rect 18932 10248 18938 10260
rect 19610 10248 19616 10260
rect 18932 10220 19616 10248
rect 18932 10208 18938 10220
rect 19610 10208 19616 10220
rect 19668 10208 19674 10260
rect 12894 10140 12900 10192
rect 12952 10189 12958 10192
rect 12952 10183 13001 10189
rect 12952 10149 12955 10183
rect 12989 10180 13001 10183
rect 13078 10180 13084 10192
rect 12989 10152 13084 10180
rect 12989 10149 13001 10152
rect 12952 10143 13001 10149
rect 12952 10140 12958 10143
rect 13078 10140 13084 10152
rect 13136 10140 13142 10192
rect 13814 10140 13820 10192
rect 13872 10180 13878 10192
rect 15657 10183 15715 10189
rect 15657 10180 15669 10183
rect 13872 10152 15669 10180
rect 13872 10140 13878 10152
rect 15657 10149 15669 10152
rect 15703 10149 15715 10183
rect 15657 10143 15715 10149
rect 15749 10183 15807 10189
rect 15749 10149 15761 10183
rect 15795 10180 15807 10183
rect 16850 10180 16856 10192
rect 15795 10152 16856 10180
rect 15795 10149 15807 10152
rect 15749 10143 15807 10149
rect 16850 10140 16856 10152
rect 16908 10140 16914 10192
rect 19242 10140 19248 10192
rect 19300 10180 19306 10192
rect 19797 10183 19855 10189
rect 19797 10180 19809 10183
rect 19300 10152 19809 10180
rect 19300 10140 19306 10152
rect 19797 10149 19809 10152
rect 19843 10149 19855 10183
rect 19797 10143 19855 10149
rect 13170 10072 13176 10124
rect 13228 10112 13234 10124
rect 14550 10112 14556 10124
rect 13228 10084 13308 10112
rect 14511 10084 14556 10112
rect 13228 10072 13234 10084
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 11480 10016 12817 10044
rect 11480 10004 11486 10016
rect 12805 10013 12817 10016
rect 12851 10013 12863 10047
rect 12805 10007 12863 10013
rect 13078 10004 13084 10056
rect 13136 10044 13142 10056
rect 13280 10053 13308 10084
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 14645 10115 14703 10121
rect 14645 10081 14657 10115
rect 14691 10112 14703 10115
rect 14826 10112 14832 10124
rect 14691 10084 14832 10112
rect 14691 10081 14703 10084
rect 14645 10075 14703 10081
rect 14826 10072 14832 10084
rect 14884 10072 14890 10124
rect 13265 10047 13323 10053
rect 13136 10016 13181 10044
rect 13136 10004 13142 10016
rect 13265 10013 13277 10047
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 14737 10047 14795 10053
rect 14737 10013 14749 10047
rect 14783 10044 14795 10047
rect 15381 10047 15439 10053
rect 15381 10044 15393 10047
rect 14783 10016 15393 10044
rect 14783 10013 14795 10016
rect 14737 10007 14795 10013
rect 15381 10013 15393 10016
rect 15427 10013 15439 10047
rect 15562 10044 15568 10056
rect 15523 10016 15568 10044
rect 15381 10007 15439 10013
rect 13173 9979 13231 9985
rect 13173 9945 13185 9979
rect 13219 9976 13231 9979
rect 14476 9976 14504 10007
rect 15562 10004 15568 10016
rect 15620 10004 15626 10056
rect 15841 10047 15899 10053
rect 15841 10013 15853 10047
rect 15887 10013 15899 10047
rect 15841 10007 15899 10013
rect 16025 10047 16083 10053
rect 16025 10013 16037 10047
rect 16071 10044 16083 10047
rect 16298 10044 16304 10056
rect 16071 10016 16304 10044
rect 16071 10013 16083 10016
rect 16025 10007 16083 10013
rect 13219 9948 14504 9976
rect 13219 9945 13231 9948
rect 13173 9939 13231 9945
rect 14642 9936 14648 9988
rect 14700 9976 14706 9988
rect 15856 9976 15884 10007
rect 16298 10004 16304 10016
rect 16356 10004 16362 10056
rect 17405 10047 17463 10053
rect 17405 10013 17417 10047
rect 17451 10013 17463 10047
rect 17862 10044 17868 10056
rect 17823 10016 17868 10044
rect 17405 10007 17463 10013
rect 14700 9948 15884 9976
rect 16485 9979 16543 9985
rect 14700 9936 14706 9948
rect 16485 9945 16497 9979
rect 16531 9945 16543 9979
rect 16485 9939 16543 9945
rect 6457 9911 6515 9917
rect 6457 9877 6469 9911
rect 6503 9908 6515 9911
rect 7834 9908 7840 9920
rect 6503 9880 7840 9908
rect 6503 9877 6515 9880
rect 6457 9871 6515 9877
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 14274 9908 14280 9920
rect 14235 9880 14280 9908
rect 14274 9868 14280 9880
rect 14332 9868 14338 9920
rect 15378 9868 15384 9920
rect 15436 9908 15442 9920
rect 16500 9908 16528 9939
rect 16666 9936 16672 9988
rect 16724 9985 16730 9988
rect 16724 9979 16743 9985
rect 16731 9945 16743 9979
rect 17420 9976 17448 10007
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 18046 10044 18052 10056
rect 18007 10016 18052 10044
rect 18046 10004 18052 10016
rect 18104 10044 18110 10056
rect 18104 10016 19564 10044
rect 18104 10004 18110 10016
rect 17954 9976 17960 9988
rect 17420 9948 17960 9976
rect 16724 9939 16743 9945
rect 16724 9936 16730 9939
rect 17954 9936 17960 9948
rect 18012 9936 18018 9988
rect 19426 9976 19432 9988
rect 19387 9948 19432 9976
rect 19426 9936 19432 9948
rect 19484 9936 19490 9988
rect 19536 9976 19564 10016
rect 19629 9979 19687 9985
rect 19629 9976 19641 9979
rect 19536 9948 19641 9976
rect 19629 9945 19641 9948
rect 19675 9945 19687 9979
rect 19629 9939 19687 9945
rect 17586 9908 17592 9920
rect 15436 9880 16528 9908
rect 17547 9880 17592 9908
rect 15436 9868 15442 9880
rect 17586 9868 17592 9880
rect 17644 9868 17650 9920
rect 1104 9818 21043 9840
rect 1104 9766 5894 9818
rect 5946 9766 5958 9818
rect 6010 9766 6022 9818
rect 6074 9766 6086 9818
rect 6138 9766 6150 9818
rect 6202 9766 10839 9818
rect 10891 9766 10903 9818
rect 10955 9766 10967 9818
rect 11019 9766 11031 9818
rect 11083 9766 11095 9818
rect 11147 9766 15784 9818
rect 15836 9766 15848 9818
rect 15900 9766 15912 9818
rect 15964 9766 15976 9818
rect 16028 9766 16040 9818
rect 16092 9766 20729 9818
rect 20781 9766 20793 9818
rect 20845 9766 20857 9818
rect 20909 9766 20921 9818
rect 20973 9766 20985 9818
rect 21037 9766 21043 9818
rect 1104 9744 21043 9766
rect 13078 9704 13084 9716
rect 13039 9676 13084 9704
rect 13078 9664 13084 9676
rect 13136 9664 13142 9716
rect 17310 9704 17316 9716
rect 16684 9676 17316 9704
rect 3044 9639 3102 9645
rect 3044 9605 3056 9639
rect 3090 9636 3102 9639
rect 3786 9636 3792 9648
rect 3090 9608 3792 9636
rect 3090 9605 3102 9608
rect 3044 9599 3102 9605
rect 3786 9596 3792 9608
rect 3844 9596 3850 9648
rect 14182 9636 14188 9648
rect 13188 9608 14188 9636
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 8846 9568 8852 9580
rect 8067 9540 8852 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 8846 9528 8852 9540
rect 8904 9528 8910 9580
rect 12986 9568 12992 9580
rect 12947 9540 12992 9568
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 13188 9577 13216 9608
rect 14182 9596 14188 9608
rect 14240 9596 14246 9648
rect 15378 9596 15384 9648
rect 15436 9636 15442 9648
rect 15473 9639 15531 9645
rect 15473 9636 15485 9639
rect 15436 9608 15485 9636
rect 15436 9596 15442 9608
rect 15473 9605 15485 9608
rect 15519 9605 15531 9639
rect 16684 9636 16712 9676
rect 17310 9664 17316 9676
rect 17368 9704 17374 9716
rect 17368 9676 18644 9704
rect 17368 9664 17374 9676
rect 16850 9636 16856 9648
rect 15473 9599 15531 9605
rect 15948 9608 16712 9636
rect 16811 9608 16856 9636
rect 13173 9571 13231 9577
rect 13173 9537 13185 9571
rect 13219 9537 13231 9571
rect 13173 9531 13231 9537
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 13780 9540 14289 9568
rect 13780 9528 13786 9540
rect 14277 9537 14289 9540
rect 14323 9537 14335 9571
rect 14458 9568 14464 9580
rect 14419 9540 14464 9568
rect 14277 9531 14335 9537
rect 14458 9528 14464 9540
rect 14516 9528 14522 9580
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9537 15163 9571
rect 15286 9568 15292 9580
rect 15247 9540 15292 9568
rect 15105 9531 15163 9537
rect 1578 9460 1584 9512
rect 1636 9500 1642 9512
rect 2774 9500 2780 9512
rect 1636 9472 2780 9500
rect 1636 9460 1642 9472
rect 2774 9460 2780 9472
rect 2832 9500 2838 9512
rect 2832 9472 2877 9500
rect 2832 9460 2838 9472
rect 7006 9460 7012 9512
rect 7064 9500 7070 9512
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 7064 9472 7757 9500
rect 7064 9460 7070 9472
rect 7745 9469 7757 9472
rect 7791 9469 7803 9503
rect 7745 9463 7803 9469
rect 12894 9460 12900 9512
rect 12952 9500 12958 9512
rect 15120 9500 15148 9531
rect 15286 9528 15292 9540
rect 15344 9568 15350 9580
rect 15948 9568 15976 9608
rect 16850 9596 16856 9608
rect 16908 9596 16914 9648
rect 17586 9636 17592 9648
rect 17052 9608 17592 9636
rect 15344 9540 15976 9568
rect 16117 9571 16175 9577
rect 15344 9528 15350 9540
rect 16117 9537 16129 9571
rect 16163 9568 16175 9571
rect 16206 9568 16212 9580
rect 16163 9540 16212 9568
rect 16163 9537 16175 9540
rect 16117 9531 16175 9537
rect 16206 9528 16212 9540
rect 16264 9528 16270 9580
rect 17052 9577 17080 9608
rect 17586 9596 17592 9608
rect 17644 9596 17650 9648
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 17052 9500 17080 9531
rect 17126 9528 17132 9580
rect 17184 9568 17190 9580
rect 17184 9540 17229 9568
rect 17184 9528 17190 9540
rect 18046 9528 18052 9580
rect 18104 9568 18110 9580
rect 18509 9571 18567 9577
rect 18509 9568 18521 9571
rect 18104 9540 18521 9568
rect 18104 9528 18110 9540
rect 18509 9537 18521 9540
rect 18555 9537 18567 9571
rect 18616 9568 18644 9676
rect 18874 9568 18880 9580
rect 18616 9540 18880 9568
rect 18509 9531 18567 9537
rect 18874 9528 18880 9540
rect 18932 9528 18938 9580
rect 12952 9472 17080 9500
rect 12952 9460 12958 9472
rect 4157 9435 4215 9441
rect 4157 9401 4169 9435
rect 4203 9432 4215 9435
rect 4614 9432 4620 9444
rect 4203 9404 4620 9432
rect 4203 9401 4215 9404
rect 4157 9395 4215 9401
rect 4614 9392 4620 9404
rect 4672 9392 4678 9444
rect 16853 9435 16911 9441
rect 16853 9401 16865 9435
rect 16899 9432 16911 9435
rect 16942 9432 16948 9444
rect 16899 9404 16948 9432
rect 16899 9401 16911 9404
rect 16853 9395 16911 9401
rect 16942 9392 16948 9404
rect 17000 9392 17006 9444
rect 19518 9392 19524 9444
rect 19576 9432 19582 9444
rect 19705 9435 19763 9441
rect 19705 9432 19717 9435
rect 19576 9404 19717 9432
rect 19576 9392 19582 9404
rect 19705 9401 19717 9404
rect 19751 9401 19763 9435
rect 19705 9395 19763 9401
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 9125 9367 9183 9373
rect 9125 9364 9137 9367
rect 6788 9336 9137 9364
rect 6788 9324 6794 9336
rect 9125 9333 9137 9336
rect 9171 9333 9183 9367
rect 9125 9327 9183 9333
rect 14090 9324 14096 9376
rect 14148 9364 14154 9376
rect 14369 9367 14427 9373
rect 14369 9364 14381 9367
rect 14148 9336 14381 9364
rect 14148 9324 14154 9336
rect 14369 9333 14381 9336
rect 14415 9333 14427 9367
rect 14369 9327 14427 9333
rect 16209 9367 16267 9373
rect 16209 9333 16221 9367
rect 16255 9364 16267 9367
rect 16666 9364 16672 9376
rect 16255 9336 16672 9364
rect 16255 9333 16267 9336
rect 16209 9327 16267 9333
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 1104 9274 20884 9296
rect 1104 9222 3422 9274
rect 3474 9222 3486 9274
rect 3538 9222 3550 9274
rect 3602 9222 3614 9274
rect 3666 9222 3678 9274
rect 3730 9222 8367 9274
rect 8419 9222 8431 9274
rect 8483 9222 8495 9274
rect 8547 9222 8559 9274
rect 8611 9222 8623 9274
rect 8675 9222 13312 9274
rect 13364 9222 13376 9274
rect 13428 9222 13440 9274
rect 13492 9222 13504 9274
rect 13556 9222 13568 9274
rect 13620 9222 18257 9274
rect 18309 9222 18321 9274
rect 18373 9222 18385 9274
rect 18437 9222 18449 9274
rect 18501 9222 18513 9274
rect 18565 9222 20884 9274
rect 1104 9200 20884 9222
rect 2866 9120 2872 9172
rect 2924 9160 2930 9172
rect 2961 9163 3019 9169
rect 2961 9160 2973 9163
rect 2924 9132 2973 9160
rect 2924 9120 2930 9132
rect 2961 9129 2973 9132
rect 3007 9129 3019 9163
rect 2961 9123 3019 9129
rect 5997 9163 6055 9169
rect 5997 9129 6009 9163
rect 6043 9160 6055 9163
rect 6914 9160 6920 9172
rect 6043 9132 6920 9160
rect 6043 9129 6055 9132
rect 5997 9123 6055 9129
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 8481 9163 8539 9169
rect 8481 9129 8493 9163
rect 8527 9160 8539 9163
rect 11514 9160 11520 9172
rect 8527 9132 11520 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 11701 9163 11759 9169
rect 11701 9129 11713 9163
rect 11747 9160 11759 9163
rect 12342 9160 12348 9172
rect 11747 9132 12348 9160
rect 11747 9129 11759 9132
rect 11701 9123 11759 9129
rect 12342 9120 12348 9132
rect 12400 9160 12406 9172
rect 15286 9160 15292 9172
rect 12400 9132 15292 9160
rect 12400 9120 12406 9132
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 17865 9163 17923 9169
rect 17865 9129 17877 9163
rect 17911 9160 17923 9163
rect 18046 9160 18052 9172
rect 17911 9132 18052 9160
rect 17911 9129 17923 9132
rect 17865 9123 17923 9129
rect 18046 9120 18052 9132
rect 18104 9120 18110 9172
rect 19886 9160 19892 9172
rect 19847 9132 19892 9160
rect 19886 9120 19892 9132
rect 19944 9120 19950 9172
rect 17954 9052 17960 9104
rect 18012 9092 18018 9104
rect 19705 9095 19763 9101
rect 19705 9092 19717 9095
rect 18012 9064 19717 9092
rect 18012 9052 18018 9064
rect 19705 9061 19717 9064
rect 19751 9061 19763 9095
rect 19705 9055 19763 9061
rect 1578 9024 1584 9036
rect 1539 8996 1584 9024
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 7006 8984 7012 9036
rect 7064 9024 7070 9036
rect 7101 9027 7159 9033
rect 7101 9024 7113 9027
rect 7064 8996 7113 9024
rect 7064 8984 7070 8996
rect 7101 8993 7113 8996
rect 7147 8993 7159 9027
rect 7101 8987 7159 8993
rect 10413 9027 10471 9033
rect 10413 8993 10425 9027
rect 10459 9024 10471 9027
rect 11422 9024 11428 9036
rect 10459 8996 11428 9024
rect 10459 8993 10471 8996
rect 10413 8987 10471 8993
rect 11422 8984 11428 8996
rect 11480 8984 11486 9036
rect 16206 8984 16212 9036
rect 16264 9024 16270 9036
rect 16264 8996 17448 9024
rect 16264 8984 16270 8996
rect 1854 8965 1860 8968
rect 1848 8956 1860 8965
rect 1815 8928 1860 8956
rect 1848 8919 1860 8928
rect 1854 8916 1860 8919
rect 1912 8916 1918 8968
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 4890 8965 4896 8968
rect 4617 8959 4675 8965
rect 4617 8956 4629 8959
rect 3936 8928 4629 8956
rect 3936 8916 3942 8928
rect 4617 8925 4629 8928
rect 4663 8925 4675 8959
rect 4884 8956 4896 8965
rect 4851 8928 4896 8956
rect 4617 8919 4675 8925
rect 4884 8919 4896 8928
rect 4890 8916 4896 8919
rect 4948 8916 4954 8968
rect 7368 8959 7426 8965
rect 7368 8925 7380 8959
rect 7414 8956 7426 8959
rect 8202 8956 8208 8968
rect 7414 8928 8208 8956
rect 7414 8925 7426 8928
rect 7368 8919 7426 8925
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 9766 8916 9772 8968
rect 9824 8956 9830 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9824 8928 10149 8956
rect 9824 8916 9830 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 14369 8959 14427 8965
rect 14369 8956 14381 8959
rect 13780 8928 14381 8956
rect 13780 8916 13786 8928
rect 14369 8925 14381 8928
rect 14415 8925 14427 8959
rect 16574 8956 16580 8968
rect 16535 8928 16580 8956
rect 14369 8919 14427 8925
rect 16574 8916 16580 8928
rect 16632 8916 16638 8968
rect 16942 8956 16948 8968
rect 16903 8928 16948 8956
rect 16942 8916 16948 8928
rect 17000 8916 17006 8968
rect 17034 8916 17040 8968
rect 17092 8956 17098 8968
rect 17420 8965 17448 8996
rect 18046 8984 18052 9036
rect 18104 9024 18110 9036
rect 19429 9027 19487 9033
rect 19429 9024 19441 9027
rect 18104 8996 19441 9024
rect 18104 8984 18110 8996
rect 19429 8993 19441 8996
rect 19475 8993 19487 9027
rect 19429 8987 19487 8993
rect 17405 8959 17463 8965
rect 17092 8928 17137 8956
rect 17092 8916 17098 8928
rect 17405 8925 17417 8959
rect 17451 8925 17463 8959
rect 17405 8919 17463 8925
rect 17497 8959 17555 8965
rect 17497 8925 17509 8959
rect 17543 8956 17555 8959
rect 18598 8956 18604 8968
rect 17543 8928 18604 8956
rect 17543 8925 17555 8928
rect 17497 8919 17555 8925
rect 14458 8848 14464 8900
rect 14516 8888 14522 8900
rect 14553 8891 14611 8897
rect 14553 8888 14565 8891
rect 14516 8860 14565 8888
rect 14516 8848 14522 8860
rect 14553 8857 14565 8860
rect 14599 8857 14611 8891
rect 17420 8888 17448 8919
rect 18598 8916 18604 8928
rect 18656 8916 18662 8968
rect 18874 8888 18880 8900
rect 17420 8860 18880 8888
rect 14553 8851 14611 8857
rect 18874 8848 18880 8860
rect 18932 8848 18938 8900
rect 13998 8780 14004 8832
rect 14056 8820 14062 8832
rect 14737 8823 14795 8829
rect 14737 8820 14749 8823
rect 14056 8792 14749 8820
rect 14056 8780 14062 8792
rect 14737 8789 14749 8792
rect 14783 8789 14795 8823
rect 14737 8783 14795 8789
rect 1104 8730 21043 8752
rect 1104 8678 5894 8730
rect 5946 8678 5958 8730
rect 6010 8678 6022 8730
rect 6074 8678 6086 8730
rect 6138 8678 6150 8730
rect 6202 8678 10839 8730
rect 10891 8678 10903 8730
rect 10955 8678 10967 8730
rect 11019 8678 11031 8730
rect 11083 8678 11095 8730
rect 11147 8678 15784 8730
rect 15836 8678 15848 8730
rect 15900 8678 15912 8730
rect 15964 8678 15976 8730
rect 16028 8678 16040 8730
rect 16092 8678 20729 8730
rect 20781 8678 20793 8730
rect 20845 8678 20857 8730
rect 20909 8678 20921 8730
rect 20973 8678 20985 8730
rect 21037 8678 21043 8730
rect 1104 8656 21043 8678
rect 4341 8619 4399 8625
rect 4341 8585 4353 8619
rect 4387 8616 4399 8619
rect 5534 8616 5540 8628
rect 4387 8588 5540 8616
rect 4387 8585 4399 8588
rect 4341 8579 4399 8585
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8616 11207 8619
rect 16574 8616 16580 8628
rect 11195 8588 16580 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 16574 8576 16580 8588
rect 16632 8616 16638 8628
rect 16632 8588 17908 8616
rect 16632 8576 16638 8588
rect 3234 8557 3240 8560
rect 3228 8548 3240 8557
rect 3195 8520 3240 8548
rect 3228 8511 3240 8520
rect 3234 8508 3240 8511
rect 3292 8508 3298 8560
rect 10036 8551 10094 8557
rect 10036 8517 10048 8551
rect 10082 8548 10094 8551
rect 12894 8548 12900 8560
rect 10082 8520 12900 8548
rect 10082 8517 10094 8520
rect 10036 8511 10094 8517
rect 12894 8508 12900 8520
rect 12952 8508 12958 8560
rect 13630 8548 13636 8560
rect 13188 8520 13636 8548
rect 7926 8440 7932 8492
rect 7984 8480 7990 8492
rect 13188 8489 13216 8520
rect 13630 8508 13636 8520
rect 13688 8548 13694 8560
rect 14185 8551 14243 8557
rect 14185 8548 14197 8551
rect 13688 8520 14197 8548
rect 13688 8508 13694 8520
rect 14185 8517 14197 8520
rect 14231 8548 14243 8551
rect 16942 8548 16948 8560
rect 14231 8520 16948 8548
rect 14231 8517 14243 8520
rect 14185 8511 14243 8517
rect 16942 8508 16948 8520
rect 17000 8548 17006 8560
rect 17221 8551 17279 8557
rect 17221 8548 17233 8551
rect 17000 8520 17233 8548
rect 17000 8508 17006 8520
rect 17221 8517 17233 8520
rect 17267 8517 17279 8551
rect 17880 8548 17908 8588
rect 17954 8576 17960 8628
rect 18012 8616 18018 8628
rect 18233 8619 18291 8625
rect 18233 8616 18245 8619
rect 18012 8588 18245 8616
rect 18012 8576 18018 8588
rect 18233 8585 18245 8588
rect 18279 8585 18291 8619
rect 18233 8579 18291 8585
rect 18432 8588 19012 8616
rect 18432 8548 18460 8588
rect 17880 8520 18460 8548
rect 18509 8551 18567 8557
rect 17221 8511 17279 8517
rect 18509 8517 18521 8551
rect 18555 8548 18567 8551
rect 18690 8548 18696 8560
rect 18555 8520 18696 8548
rect 18555 8517 18567 8520
rect 18509 8511 18567 8517
rect 18690 8508 18696 8520
rect 18748 8508 18754 8560
rect 13173 8483 13231 8489
rect 7984 8452 12434 8480
rect 7984 8440 7990 8452
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 2961 8415 3019 8421
rect 2961 8412 2973 8415
rect 2832 8384 2973 8412
rect 2832 8372 2838 8384
rect 2961 8381 2973 8384
rect 3007 8381 3019 8415
rect 9766 8412 9772 8424
rect 9727 8384 9772 8412
rect 2961 8375 3019 8381
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 12406 8412 12434 8452
rect 13173 8449 13185 8483
rect 13219 8449 13231 8483
rect 13173 8443 13231 8449
rect 13357 8483 13415 8489
rect 13357 8449 13369 8483
rect 13403 8480 13415 8483
rect 13722 8480 13728 8492
rect 13403 8452 13728 8480
rect 13403 8449 13415 8452
rect 13357 8443 13415 8449
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 13998 8480 14004 8492
rect 13959 8452 14004 8480
rect 13998 8440 14004 8452
rect 14056 8440 14062 8492
rect 14090 8440 14096 8492
rect 14148 8480 14154 8492
rect 14323 8483 14381 8489
rect 14148 8452 14193 8480
rect 14148 8440 14154 8452
rect 14323 8449 14335 8483
rect 14369 8480 14381 8483
rect 15194 8480 15200 8492
rect 14369 8452 15200 8480
rect 14369 8449 14381 8452
rect 14323 8443 14381 8449
rect 15194 8440 15200 8452
rect 15252 8440 15258 8492
rect 16850 8480 16856 8492
rect 16811 8452 16856 8480
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8449 17095 8483
rect 17037 8443 17095 8449
rect 18417 8483 18475 8489
rect 18417 8449 18429 8483
rect 18463 8449 18475 8483
rect 18417 8443 18475 8449
rect 14461 8415 14519 8421
rect 14461 8412 14473 8415
rect 12406 8384 14473 8412
rect 14461 8381 14473 8384
rect 14507 8412 14519 8415
rect 16666 8412 16672 8424
rect 14507 8384 16672 8412
rect 14507 8381 14519 8384
rect 14461 8375 14519 8381
rect 16666 8372 16672 8384
rect 16724 8412 16730 8424
rect 17052 8412 17080 8443
rect 17126 8412 17132 8424
rect 16724 8384 17132 8412
rect 16724 8372 16730 8384
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 18432 8412 18460 8443
rect 18598 8440 18604 8492
rect 18656 8480 18662 8492
rect 18785 8483 18843 8489
rect 18656 8452 18749 8480
rect 18656 8440 18662 8452
rect 18432 8384 18644 8412
rect 18616 8356 18644 8384
rect 13170 8304 13176 8356
rect 13228 8344 13234 8356
rect 13265 8347 13323 8353
rect 13265 8344 13277 8347
rect 13228 8316 13277 8344
rect 13228 8304 13234 8316
rect 13265 8313 13277 8316
rect 13311 8313 13323 8347
rect 13265 8307 13323 8313
rect 18598 8304 18604 8356
rect 18656 8304 18662 8356
rect 13814 8276 13820 8288
rect 13775 8248 13820 8276
rect 13814 8236 13820 8248
rect 13872 8236 13878 8288
rect 18708 8276 18736 8452
rect 18785 8449 18797 8483
rect 18831 8449 18843 8483
rect 18785 8443 18843 8449
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8480 18935 8483
rect 18984 8480 19012 8588
rect 18923 8452 19012 8480
rect 18923 8449 18935 8452
rect 18877 8443 18935 8449
rect 18800 8344 18828 8443
rect 18874 8344 18880 8356
rect 18800 8316 18880 8344
rect 18874 8304 18880 8316
rect 18932 8304 18938 8356
rect 19610 8276 19616 8288
rect 18708 8248 19616 8276
rect 19610 8236 19616 8248
rect 19668 8236 19674 8288
rect 1104 8186 20884 8208
rect 1104 8134 3422 8186
rect 3474 8134 3486 8186
rect 3538 8134 3550 8186
rect 3602 8134 3614 8186
rect 3666 8134 3678 8186
rect 3730 8134 8367 8186
rect 8419 8134 8431 8186
rect 8483 8134 8495 8186
rect 8547 8134 8559 8186
rect 8611 8134 8623 8186
rect 8675 8134 13312 8186
rect 13364 8134 13376 8186
rect 13428 8134 13440 8186
rect 13492 8134 13504 8186
rect 13556 8134 13568 8186
rect 13620 8134 18257 8186
rect 18309 8134 18321 8186
rect 18373 8134 18385 8186
rect 18437 8134 18449 8186
rect 18501 8134 18513 8186
rect 18565 8134 20884 8186
rect 1104 8112 20884 8134
rect 6181 8075 6239 8081
rect 6181 8041 6193 8075
rect 6227 8072 6239 8075
rect 7374 8072 7380 8084
rect 6227 8044 7380 8072
rect 6227 8041 6239 8044
rect 6181 8035 6239 8041
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 8018 8032 8024 8084
rect 8076 8072 8082 8084
rect 8389 8075 8447 8081
rect 8389 8072 8401 8075
rect 8076 8044 8401 8072
rect 8076 8032 8082 8044
rect 8389 8041 8401 8044
rect 8435 8041 8447 8075
rect 8389 8035 8447 8041
rect 11333 8075 11391 8081
rect 11333 8041 11345 8075
rect 11379 8072 11391 8075
rect 14458 8072 14464 8084
rect 11379 8044 14464 8072
rect 11379 8041 11391 8044
rect 11333 8035 11391 8041
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 15194 8032 15200 8084
rect 15252 8072 15258 8084
rect 15565 8075 15623 8081
rect 15565 8072 15577 8075
rect 15252 8044 15577 8072
rect 15252 8032 15258 8044
rect 15565 8041 15577 8044
rect 15611 8041 15623 8075
rect 15565 8035 15623 8041
rect 16945 8075 17003 8081
rect 16945 8041 16957 8075
rect 16991 8072 17003 8075
rect 17034 8072 17040 8084
rect 16991 8044 17040 8072
rect 16991 8041 17003 8044
rect 16945 8035 17003 8041
rect 17034 8032 17040 8044
rect 17092 8032 17098 8084
rect 16114 8004 16120 8016
rect 12406 7976 16120 8004
rect 7006 7936 7012 7948
rect 6967 7908 7012 7936
rect 7006 7896 7012 7908
rect 7064 7896 7070 7948
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 9953 7939 10011 7945
rect 9953 7936 9965 7939
rect 9824 7908 9965 7936
rect 9824 7896 9830 7908
rect 9953 7905 9965 7908
rect 9999 7905 10011 7939
rect 9953 7899 10011 7905
rect 3878 7828 3884 7880
rect 3936 7868 3942 7880
rect 4801 7871 4859 7877
rect 4801 7868 4813 7871
rect 3936 7840 4813 7868
rect 3936 7828 3942 7840
rect 4801 7837 4813 7840
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 7276 7871 7334 7877
rect 7276 7837 7288 7871
rect 7322 7868 7334 7871
rect 12406 7868 12434 7976
rect 16114 7964 16120 7976
rect 16172 7964 16178 8016
rect 18690 8004 18696 8016
rect 18616 7976 18696 8004
rect 13262 7896 13268 7948
rect 13320 7936 13326 7948
rect 18616 7945 18644 7976
rect 18690 7964 18696 7976
rect 18748 7964 18754 8016
rect 18874 7964 18880 8016
rect 18932 8004 18938 8016
rect 18932 7976 19564 8004
rect 18932 7964 18938 7976
rect 17589 7939 17647 7945
rect 13320 7908 13365 7936
rect 13320 7896 13326 7908
rect 17589 7905 17601 7939
rect 17635 7936 17647 7939
rect 18601 7939 18659 7945
rect 18601 7936 18613 7939
rect 17635 7908 18613 7936
rect 17635 7905 17647 7908
rect 17589 7899 17647 7905
rect 18601 7905 18613 7908
rect 18647 7936 18659 7939
rect 18647 7908 19472 7936
rect 18647 7905 18659 7908
rect 18601 7899 18659 7905
rect 7322 7840 12434 7868
rect 13081 7871 13139 7877
rect 7322 7837 7334 7840
rect 7276 7831 7334 7837
rect 13081 7837 13093 7871
rect 13127 7868 13139 7871
rect 13814 7868 13820 7880
rect 13127 7840 13820 7868
rect 13127 7837 13139 7840
rect 13081 7831 13139 7837
rect 13814 7828 13820 7840
rect 13872 7828 13878 7880
rect 15197 7871 15255 7877
rect 15197 7837 15209 7871
rect 15243 7868 15255 7871
rect 15286 7868 15292 7880
rect 15243 7840 15292 7868
rect 15243 7837 15255 7840
rect 15197 7831 15255 7837
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 15562 7868 15568 7880
rect 15523 7840 15568 7868
rect 15562 7828 15568 7840
rect 15620 7828 15626 7880
rect 16853 7871 16911 7877
rect 16853 7837 16865 7871
rect 16899 7868 16911 7871
rect 16942 7868 16948 7880
rect 16899 7840 16948 7868
rect 16899 7837 16911 7840
rect 16853 7831 16911 7837
rect 16942 7828 16948 7840
rect 17000 7828 17006 7880
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7868 17095 7871
rect 17126 7868 17132 7880
rect 17083 7840 17132 7868
rect 17083 7837 17095 7840
rect 17037 7831 17095 7837
rect 17126 7828 17132 7840
rect 17184 7828 17190 7880
rect 17497 7871 17555 7877
rect 17497 7837 17509 7871
rect 17543 7837 17555 7871
rect 18506 7868 18512 7880
rect 18467 7840 18512 7868
rect 17497 7831 17555 7837
rect 5068 7803 5126 7809
rect 5068 7769 5080 7803
rect 5114 7800 5126 7803
rect 9490 7800 9496 7812
rect 5114 7772 9496 7800
rect 5114 7769 5126 7772
rect 5068 7763 5126 7769
rect 9490 7760 9496 7772
rect 9548 7760 9554 7812
rect 10220 7803 10278 7809
rect 10220 7769 10232 7803
rect 10266 7800 10278 7803
rect 14274 7800 14280 7812
rect 10266 7772 14280 7800
rect 10266 7769 10278 7772
rect 10220 7763 10278 7769
rect 14274 7760 14280 7772
rect 14332 7760 14338 7812
rect 17512 7800 17540 7831
rect 18506 7828 18512 7840
rect 18564 7828 18570 7880
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7868 18843 7871
rect 18874 7868 18880 7880
rect 18831 7840 18880 7868
rect 18831 7837 18843 7840
rect 18785 7831 18843 7837
rect 16868 7772 17540 7800
rect 18708 7800 18736 7831
rect 18874 7828 18880 7840
rect 18932 7828 18938 7880
rect 19444 7877 19472 7908
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7837 19487 7871
rect 19536 7868 19564 7976
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 19536 7840 19625 7868
rect 19429 7831 19487 7837
rect 19613 7837 19625 7840
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 18708 7772 19656 7800
rect 16868 7744 16896 7772
rect 19628 7744 19656 7772
rect 12618 7732 12624 7744
rect 12579 7704 12624 7732
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 12989 7735 13047 7741
rect 12989 7701 13001 7735
rect 13035 7732 13047 7735
rect 13722 7732 13728 7744
rect 13035 7704 13728 7732
rect 13035 7701 13047 7704
rect 12989 7695 13047 7701
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 15381 7735 15439 7741
rect 15381 7701 15393 7735
rect 15427 7732 15439 7735
rect 16850 7732 16856 7744
rect 15427 7704 16856 7732
rect 15427 7701 15439 7704
rect 15381 7695 15439 7701
rect 16850 7692 16856 7704
rect 16908 7692 16914 7744
rect 18325 7735 18383 7741
rect 18325 7701 18337 7735
rect 18371 7732 18383 7735
rect 18598 7732 18604 7744
rect 18371 7704 18604 7732
rect 18371 7701 18383 7704
rect 18325 7695 18383 7701
rect 18598 7692 18604 7704
rect 18656 7692 18662 7744
rect 18782 7692 18788 7744
rect 18840 7732 18846 7744
rect 19521 7735 19579 7741
rect 19521 7732 19533 7735
rect 18840 7704 19533 7732
rect 18840 7692 18846 7704
rect 19521 7701 19533 7704
rect 19567 7701 19579 7735
rect 19521 7695 19579 7701
rect 19610 7692 19616 7744
rect 19668 7692 19674 7744
rect 1104 7642 21043 7664
rect 1104 7590 5894 7642
rect 5946 7590 5958 7642
rect 6010 7590 6022 7642
rect 6074 7590 6086 7642
rect 6138 7590 6150 7642
rect 6202 7590 10839 7642
rect 10891 7590 10903 7642
rect 10955 7590 10967 7642
rect 11019 7590 11031 7642
rect 11083 7590 11095 7642
rect 11147 7590 15784 7642
rect 15836 7590 15848 7642
rect 15900 7590 15912 7642
rect 15964 7590 15976 7642
rect 16028 7590 16040 7642
rect 16092 7590 20729 7642
rect 20781 7590 20793 7642
rect 20845 7590 20857 7642
rect 20909 7590 20921 7642
rect 20973 7590 20985 7642
rect 21037 7590 21043 7642
rect 1104 7568 21043 7590
rect 7006 7488 7012 7540
rect 7064 7528 7070 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 7064 7500 9137 7528
rect 7064 7488 7070 7500
rect 9125 7497 9137 7500
rect 9171 7528 9183 7531
rect 9766 7528 9772 7540
rect 9171 7500 9772 7528
rect 9171 7497 9183 7500
rect 9125 7491 9183 7497
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 17773 7531 17831 7537
rect 17773 7497 17785 7531
rect 17819 7528 17831 7531
rect 18506 7528 18512 7540
rect 17819 7500 18512 7528
rect 17819 7497 17831 7500
rect 17773 7491 17831 7497
rect 18506 7488 18512 7500
rect 18564 7488 18570 7540
rect 15286 7460 15292 7472
rect 13004 7432 15292 7460
rect 2590 7392 2596 7404
rect 2551 7364 2596 7392
rect 2590 7352 2596 7364
rect 2648 7352 2654 7404
rect 7834 7392 7840 7404
rect 7795 7364 7840 7392
rect 7834 7352 7840 7364
rect 7892 7352 7898 7404
rect 12894 7352 12900 7404
rect 12952 7392 12958 7404
rect 13004 7401 13032 7432
rect 15286 7420 15292 7432
rect 15344 7420 15350 7472
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12952 7364 13001 7392
rect 12952 7352 12958 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 14274 7392 14280 7404
rect 13127 7364 14280 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 15194 7392 15200 7404
rect 15155 7364 15200 7392
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 16942 7352 16948 7404
rect 17000 7392 17006 7404
rect 17681 7395 17739 7401
rect 17681 7392 17693 7395
rect 17000 7364 17693 7392
rect 17000 7352 17006 7364
rect 17681 7361 17693 7364
rect 17727 7361 17739 7395
rect 17681 7355 17739 7361
rect 13173 7327 13231 7333
rect 13173 7293 13185 7327
rect 13219 7324 13231 7327
rect 13262 7324 13268 7336
rect 13219 7296 13268 7324
rect 13219 7293 13231 7296
rect 13173 7287 13231 7293
rect 13078 7216 13084 7268
rect 13136 7256 13142 7268
rect 13188 7256 13216 7287
rect 13262 7284 13268 7296
rect 13320 7284 13326 7336
rect 15286 7324 15292 7336
rect 15247 7296 15292 7324
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 15470 7324 15476 7336
rect 15431 7296 15476 7324
rect 15470 7284 15476 7296
rect 15528 7284 15534 7336
rect 13136 7228 13216 7256
rect 13136 7216 13142 7228
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 3878 7188 3884 7200
rect 2832 7160 3884 7188
rect 2832 7148 2838 7160
rect 3878 7148 3884 7160
rect 3936 7148 3942 7200
rect 11698 7148 11704 7200
rect 11756 7188 11762 7200
rect 12621 7191 12679 7197
rect 12621 7188 12633 7191
rect 11756 7160 12633 7188
rect 11756 7148 11762 7160
rect 12621 7157 12633 7160
rect 12667 7157 12679 7191
rect 14826 7188 14832 7200
rect 14787 7160 14832 7188
rect 12621 7151 12679 7157
rect 14826 7148 14832 7160
rect 14884 7148 14890 7200
rect 1104 7098 20884 7120
rect 1104 7046 3422 7098
rect 3474 7046 3486 7098
rect 3538 7046 3550 7098
rect 3602 7046 3614 7098
rect 3666 7046 3678 7098
rect 3730 7046 8367 7098
rect 8419 7046 8431 7098
rect 8483 7046 8495 7098
rect 8547 7046 8559 7098
rect 8611 7046 8623 7098
rect 8675 7046 13312 7098
rect 13364 7046 13376 7098
rect 13428 7046 13440 7098
rect 13492 7046 13504 7098
rect 13556 7046 13568 7098
rect 13620 7046 18257 7098
rect 18309 7046 18321 7098
rect 18373 7046 18385 7098
rect 18437 7046 18449 7098
rect 18501 7046 18513 7098
rect 18565 7046 20884 7098
rect 1104 7024 20884 7046
rect 14274 6984 14280 6996
rect 14235 6956 14280 6984
rect 14274 6944 14280 6956
rect 14332 6944 14338 6996
rect 15286 6944 15292 6996
rect 15344 6984 15350 6996
rect 15473 6987 15531 6993
rect 15473 6984 15485 6987
rect 15344 6956 15485 6984
rect 15344 6944 15350 6956
rect 15473 6953 15485 6956
rect 15519 6953 15531 6987
rect 17402 6984 17408 6996
rect 17363 6956 17408 6984
rect 15473 6947 15531 6953
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 2590 6876 2596 6928
rect 2648 6916 2654 6928
rect 7285 6919 7343 6925
rect 7285 6916 7297 6919
rect 2648 6888 7297 6916
rect 2648 6876 2654 6888
rect 7285 6885 7297 6888
rect 7331 6916 7343 6919
rect 7834 6916 7840 6928
rect 7331 6888 7840 6916
rect 7331 6885 7343 6888
rect 7285 6879 7343 6885
rect 7834 6876 7840 6888
rect 7892 6876 7898 6928
rect 14458 6876 14464 6928
rect 14516 6916 14522 6928
rect 14516 6888 14964 6916
rect 14516 6876 14522 6888
rect 9766 6848 9772 6860
rect 9727 6820 9772 6848
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 14826 6848 14832 6860
rect 12406 6820 14832 6848
rect 1578 6780 1584 6792
rect 1539 6752 1584 6780
rect 1578 6740 1584 6752
rect 1636 6740 1642 6792
rect 1670 6740 1676 6792
rect 1728 6780 1734 6792
rect 1837 6783 1895 6789
rect 1837 6780 1849 6783
rect 1728 6752 1849 6780
rect 1728 6740 1734 6752
rect 1837 6749 1849 6752
rect 1883 6749 1895 6783
rect 1837 6743 1895 6749
rect 10036 6783 10094 6789
rect 10036 6749 10048 6783
rect 10082 6780 10094 6783
rect 12406 6780 12434 6820
rect 14826 6808 14832 6820
rect 14884 6808 14890 6860
rect 14936 6848 14964 6888
rect 15378 6876 15384 6928
rect 15436 6916 15442 6928
rect 15933 6919 15991 6925
rect 15933 6916 15945 6919
rect 15436 6888 15945 6916
rect 15436 6876 15442 6888
rect 15933 6885 15945 6888
rect 15979 6885 15991 6919
rect 15933 6879 15991 6885
rect 17313 6851 17371 6857
rect 14936 6820 15700 6848
rect 10082 6752 12434 6780
rect 10082 6749 10094 6752
rect 10036 6743 10094 6749
rect 13170 6740 13176 6792
rect 13228 6780 13234 6792
rect 13449 6783 13507 6789
rect 13449 6780 13461 6783
rect 13228 6752 13461 6780
rect 13228 6740 13234 6752
rect 13449 6749 13461 6752
rect 13495 6749 13507 6783
rect 13630 6780 13636 6792
rect 13591 6752 13636 6780
rect 13449 6743 13507 6749
rect 5534 6672 5540 6724
rect 5592 6712 5598 6724
rect 5997 6715 6055 6721
rect 5997 6712 6009 6715
rect 5592 6684 6009 6712
rect 5592 6672 5598 6684
rect 5997 6681 6009 6684
rect 6043 6681 6055 6715
rect 13464 6712 13492 6743
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 13722 6740 13728 6792
rect 13780 6780 13786 6792
rect 14458 6780 14464 6792
rect 13780 6752 13825 6780
rect 14419 6752 14464 6780
rect 13780 6740 13786 6752
rect 14458 6740 14464 6752
rect 14516 6740 14522 6792
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6749 14611 6783
rect 15562 6780 15568 6792
rect 14553 6743 14611 6749
rect 14844 6752 15568 6780
rect 14568 6712 14596 6743
rect 14844 6721 14872 6752
rect 15562 6740 15568 6752
rect 15620 6740 15626 6792
rect 15672 6789 15700 6820
rect 17313 6817 17325 6851
rect 17359 6848 17371 6851
rect 18782 6848 18788 6860
rect 17359 6820 18788 6848
rect 17359 6817 17371 6820
rect 17313 6811 17371 6817
rect 15657 6783 15715 6789
rect 15657 6749 15669 6783
rect 15703 6749 15715 6783
rect 15657 6743 15715 6749
rect 15749 6783 15807 6789
rect 15749 6749 15761 6783
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 16025 6783 16083 6789
rect 16025 6749 16037 6783
rect 16071 6780 16083 6783
rect 16114 6780 16120 6792
rect 16071 6752 16120 6780
rect 16071 6749 16083 6752
rect 16025 6743 16083 6749
rect 5997 6675 6055 6681
rect 12912 6684 13400 6712
rect 13464 6684 14596 6712
rect 14829 6715 14887 6721
rect 2961 6647 3019 6653
rect 2961 6613 2973 6647
rect 3007 6644 3019 6647
rect 3142 6644 3148 6656
rect 3007 6616 3148 6644
rect 3007 6613 3019 6616
rect 2961 6607 3019 6613
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 9030 6604 9036 6656
rect 9088 6644 9094 6656
rect 10318 6644 10324 6656
rect 9088 6616 10324 6644
rect 9088 6604 9094 6616
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 11149 6647 11207 6653
rect 11149 6613 11161 6647
rect 11195 6644 11207 6647
rect 12912 6644 12940 6684
rect 11195 6616 12940 6644
rect 11195 6613 11207 6616
rect 11149 6607 11207 6613
rect 12986 6604 12992 6656
rect 13044 6644 13050 6656
rect 13265 6647 13323 6653
rect 13265 6644 13277 6647
rect 13044 6616 13277 6644
rect 13044 6604 13050 6616
rect 13265 6613 13277 6616
rect 13311 6613 13323 6647
rect 13372 6644 13400 6684
rect 14829 6681 14841 6715
rect 14875 6681 14887 6715
rect 14829 6675 14887 6681
rect 14918 6672 14924 6724
rect 14976 6712 14982 6724
rect 15764 6712 15792 6743
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 17034 6740 17040 6792
rect 17092 6780 17098 6792
rect 17129 6783 17187 6789
rect 17129 6780 17141 6783
rect 17092 6752 17141 6780
rect 17092 6740 17098 6752
rect 17129 6749 17141 6752
rect 17175 6749 17187 6783
rect 17129 6743 17187 6749
rect 17328 6712 17356 6811
rect 18782 6808 18788 6820
rect 18840 6808 18846 6860
rect 17405 6783 17463 6789
rect 17405 6749 17417 6783
rect 17451 6780 17463 6783
rect 17862 6780 17868 6792
rect 17451 6752 17868 6780
rect 17451 6749 17463 6752
rect 17405 6743 17463 6749
rect 14976 6684 15021 6712
rect 15764 6684 17356 6712
rect 14976 6672 14982 6684
rect 15194 6644 15200 6656
rect 13372 6616 15200 6644
rect 13265 6607 13323 6613
rect 15194 6604 15200 6616
rect 15252 6604 15258 6656
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 17420 6644 17448 6743
rect 17862 6740 17868 6752
rect 17920 6780 17926 6792
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 17920 6752 18245 6780
rect 17920 6740 17926 6752
rect 18233 6749 18245 6752
rect 18279 6749 18291 6783
rect 18598 6780 18604 6792
rect 18559 6752 18604 6780
rect 18233 6743 18291 6749
rect 18598 6740 18604 6752
rect 18656 6740 18662 6792
rect 18690 6740 18696 6792
rect 18748 6780 18754 6792
rect 18748 6752 18793 6780
rect 18748 6740 18754 6752
rect 17276 6616 17448 6644
rect 17589 6647 17647 6653
rect 17276 6604 17282 6616
rect 17589 6613 17601 6647
rect 17635 6644 17647 6647
rect 18046 6644 18052 6656
rect 17635 6616 18052 6644
rect 17635 6613 17647 6616
rect 17589 6607 17647 6613
rect 18046 6604 18052 6616
rect 18104 6604 18110 6656
rect 18322 6644 18328 6656
rect 18283 6616 18328 6644
rect 18322 6604 18328 6616
rect 18380 6604 18386 6656
rect 1104 6554 21043 6576
rect 1104 6502 5894 6554
rect 5946 6502 5958 6554
rect 6010 6502 6022 6554
rect 6074 6502 6086 6554
rect 6138 6502 6150 6554
rect 6202 6502 10839 6554
rect 10891 6502 10903 6554
rect 10955 6502 10967 6554
rect 11019 6502 11031 6554
rect 11083 6502 11095 6554
rect 11147 6502 15784 6554
rect 15836 6502 15848 6554
rect 15900 6502 15912 6554
rect 15964 6502 15976 6554
rect 16028 6502 16040 6554
rect 16092 6502 20729 6554
rect 20781 6502 20793 6554
rect 20845 6502 20857 6554
rect 20909 6502 20921 6554
rect 20973 6502 20985 6554
rect 21037 6502 21043 6554
rect 1104 6480 21043 6502
rect 4157 6443 4215 6449
rect 4157 6409 4169 6443
rect 4203 6440 4215 6443
rect 4246 6440 4252 6452
rect 4203 6412 4252 6440
rect 4203 6409 4215 6412
rect 4157 6403 4215 6409
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 8481 6443 8539 6449
rect 8481 6409 8493 6443
rect 8527 6440 8539 6443
rect 12986 6440 12992 6452
rect 8527 6412 12434 6440
rect 12947 6412 12992 6440
rect 8527 6409 8539 6412
rect 8481 6403 8539 6409
rect 3050 6381 3056 6384
rect 3044 6372 3056 6381
rect 3011 6344 3056 6372
rect 3044 6335 3056 6344
rect 3050 6332 3056 6335
rect 3108 6332 3114 6384
rect 9766 6372 9772 6384
rect 8956 6344 9772 6372
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 8956 6313 8984 6344
rect 9766 6332 9772 6344
rect 9824 6332 9830 6384
rect 12406 6372 12434 6412
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 14829 6443 14887 6449
rect 14829 6409 14841 6443
rect 14875 6440 14887 6443
rect 15562 6440 15568 6452
rect 14875 6412 15568 6440
rect 14875 6409 14887 6412
rect 14829 6403 14887 6409
rect 15562 6400 15568 6412
rect 15620 6400 15626 6452
rect 17037 6443 17095 6449
rect 17037 6409 17049 6443
rect 17083 6409 17095 6443
rect 17037 6403 17095 6409
rect 18325 6443 18383 6449
rect 18325 6409 18337 6443
rect 18371 6440 18383 6443
rect 18690 6440 18696 6452
rect 18371 6412 18696 6440
rect 18371 6409 18383 6412
rect 18325 6403 18383 6409
rect 12897 6375 12955 6381
rect 12897 6372 12909 6375
rect 12406 6344 12909 6372
rect 12897 6341 12909 6344
rect 12943 6372 12955 6375
rect 14458 6372 14464 6384
rect 12943 6344 14464 6372
rect 12943 6341 12955 6344
rect 12897 6335 12955 6341
rect 14458 6332 14464 6344
rect 14516 6332 14522 6384
rect 7368 6307 7426 6313
rect 2832 6276 2877 6304
rect 2832 6264 2838 6276
rect 7368 6273 7380 6307
rect 7414 6304 7426 6307
rect 8941 6307 8999 6313
rect 7414 6276 8892 6304
rect 7414 6273 7426 6276
rect 7368 6267 7426 6273
rect 7098 6236 7104 6248
rect 7059 6208 7104 6236
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 8864 6100 8892 6276
rect 8941 6273 8953 6307
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 9208 6307 9266 6313
rect 9208 6273 9220 6307
rect 9254 6304 9266 6307
rect 10502 6304 10508 6316
rect 9254 6276 10508 6304
rect 9254 6273 9266 6276
rect 9208 6267 9266 6273
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 13722 6264 13728 6316
rect 13780 6304 13786 6316
rect 14645 6307 14703 6313
rect 14645 6304 14657 6307
rect 13780 6276 14657 6304
rect 13780 6264 13786 6276
rect 14645 6273 14657 6276
rect 14691 6273 14703 6307
rect 14645 6267 14703 6273
rect 15470 6264 15476 6316
rect 15528 6304 15534 6316
rect 16025 6307 16083 6313
rect 16025 6304 16037 6307
rect 15528 6276 16037 6304
rect 15528 6264 15534 6276
rect 16025 6273 16037 6276
rect 16071 6304 16083 6307
rect 17052 6304 17080 6403
rect 18690 6400 18696 6412
rect 18748 6400 18754 6452
rect 17402 6332 17408 6384
rect 17460 6372 17466 6384
rect 17460 6344 19012 6372
rect 17460 6332 17466 6344
rect 17218 6304 17224 6316
rect 16071 6276 17080 6304
rect 17179 6276 17224 6304
rect 16071 6273 16083 6276
rect 16025 6267 16083 6273
rect 17218 6264 17224 6276
rect 17276 6264 17282 6316
rect 17512 6313 17540 6344
rect 18984 6316 19012 6344
rect 17497 6307 17555 6313
rect 17497 6273 17509 6307
rect 17543 6273 17555 6307
rect 17497 6267 17555 6273
rect 17954 6264 17960 6316
rect 18012 6304 18018 6316
rect 18509 6307 18567 6313
rect 18509 6304 18521 6307
rect 18012 6276 18521 6304
rect 18012 6264 18018 6276
rect 18509 6273 18521 6276
rect 18555 6273 18567 6307
rect 18782 6304 18788 6316
rect 18743 6276 18788 6304
rect 18509 6267 18567 6273
rect 18782 6264 18788 6276
rect 18840 6264 18846 6316
rect 18966 6304 18972 6316
rect 18927 6276 18972 6304
rect 18966 6264 18972 6276
rect 19024 6264 19030 6316
rect 13078 6196 13084 6248
rect 13136 6236 13142 6248
rect 13173 6239 13231 6245
rect 13173 6236 13185 6239
rect 13136 6208 13185 6236
rect 13136 6196 13142 6208
rect 13173 6205 13185 6208
rect 13219 6236 13231 6239
rect 15488 6236 15516 6264
rect 13219 6208 15516 6236
rect 15841 6239 15899 6245
rect 13219 6205 13231 6208
rect 13173 6199 13231 6205
rect 15841 6205 15853 6239
rect 15887 6205 15899 6239
rect 15841 6199 15899 6205
rect 12529 6171 12587 6177
rect 12529 6168 12541 6171
rect 9876 6140 12541 6168
rect 9876 6100 9904 6140
rect 12529 6137 12541 6140
rect 12575 6137 12587 6171
rect 12529 6131 12587 6137
rect 13630 6128 13636 6180
rect 13688 6168 13694 6180
rect 15856 6168 15884 6199
rect 18322 6168 18328 6180
rect 13688 6140 15884 6168
rect 15948 6140 18328 6168
rect 13688 6128 13694 6140
rect 10318 6100 10324 6112
rect 8864 6072 9904 6100
rect 10279 6072 10324 6100
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 11422 6060 11428 6112
rect 11480 6100 11486 6112
rect 15948 6100 15976 6140
rect 18322 6128 18328 6140
rect 18380 6128 18386 6180
rect 11480 6072 15976 6100
rect 16209 6103 16267 6109
rect 11480 6060 11486 6072
rect 16209 6069 16221 6103
rect 16255 6100 16267 6103
rect 16666 6100 16672 6112
rect 16255 6072 16672 6100
rect 16255 6069 16267 6072
rect 16209 6063 16267 6069
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 1104 6010 20884 6032
rect 1104 5958 3422 6010
rect 3474 5958 3486 6010
rect 3538 5958 3550 6010
rect 3602 5958 3614 6010
rect 3666 5958 3678 6010
rect 3730 5958 8367 6010
rect 8419 5958 8431 6010
rect 8483 5958 8495 6010
rect 8547 5958 8559 6010
rect 8611 5958 8623 6010
rect 8675 5958 13312 6010
rect 13364 5958 13376 6010
rect 13428 5958 13440 6010
rect 13492 5958 13504 6010
rect 13556 5958 13568 6010
rect 13620 5958 18257 6010
rect 18309 5958 18321 6010
rect 18373 5958 18385 6010
rect 18437 5958 18449 6010
rect 18501 5958 18513 6010
rect 18565 5958 20884 6010
rect 1104 5936 20884 5958
rect 6733 5899 6791 5905
rect 6733 5865 6745 5899
rect 6779 5896 6791 5899
rect 11149 5899 11207 5905
rect 6779 5868 10732 5896
rect 6779 5865 6791 5868
rect 6733 5859 6791 5865
rect 10704 5828 10732 5868
rect 11149 5865 11161 5899
rect 11195 5896 11207 5899
rect 12894 5896 12900 5908
rect 11195 5868 12900 5896
rect 11195 5865 11207 5868
rect 11149 5859 11207 5865
rect 12894 5856 12900 5868
rect 12952 5856 12958 5908
rect 14369 5899 14427 5905
rect 14369 5865 14381 5899
rect 14415 5896 14427 5899
rect 14918 5896 14924 5908
rect 14415 5868 14924 5896
rect 14415 5865 14427 5868
rect 14369 5859 14427 5865
rect 14918 5856 14924 5868
rect 14976 5856 14982 5908
rect 13722 5828 13728 5840
rect 10704 5800 13728 5828
rect 13722 5788 13728 5800
rect 13780 5788 13786 5840
rect 15010 5788 15016 5840
rect 15068 5828 15074 5840
rect 17218 5828 17224 5840
rect 15068 5800 17224 5828
rect 15068 5788 15074 5800
rect 17218 5788 17224 5800
rect 17276 5788 17282 5840
rect 18966 5788 18972 5840
rect 19024 5828 19030 5840
rect 19705 5831 19763 5837
rect 19705 5828 19717 5831
rect 19024 5800 19717 5828
rect 19024 5788 19030 5800
rect 19705 5797 19717 5800
rect 19751 5797 19763 5831
rect 19705 5791 19763 5797
rect 1578 5760 1584 5772
rect 1539 5732 1584 5760
rect 1578 5720 1584 5732
rect 1636 5720 1642 5772
rect 16666 5760 16672 5772
rect 16627 5732 16672 5760
rect 16666 5720 16672 5732
rect 16724 5720 16730 5772
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 1946 5692 1952 5704
rect 1903 5664 1952 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 1946 5652 1952 5664
rect 2004 5692 2010 5704
rect 2314 5692 2320 5704
rect 2004 5664 2320 5692
rect 2004 5652 2010 5664
rect 2314 5652 2320 5664
rect 2372 5652 2378 5704
rect 4522 5652 4528 5704
rect 4580 5692 4586 5704
rect 5353 5695 5411 5701
rect 5353 5692 5365 5695
rect 4580 5664 5365 5692
rect 4580 5652 4586 5664
rect 5353 5661 5365 5664
rect 5399 5661 5411 5695
rect 5353 5655 5411 5661
rect 9582 5652 9588 5704
rect 9640 5692 9646 5704
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 9640 5664 9781 5692
rect 9640 5652 9646 5664
rect 9769 5661 9781 5664
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 9968 5664 12434 5692
rect 5620 5627 5678 5633
rect 5620 5593 5632 5627
rect 5666 5624 5678 5627
rect 9968 5624 9996 5664
rect 5666 5596 9996 5624
rect 10036 5627 10094 5633
rect 5666 5593 5678 5596
rect 5620 5587 5678 5593
rect 10036 5593 10048 5627
rect 10082 5624 10094 5627
rect 11698 5624 11704 5636
rect 10082 5596 11704 5624
rect 10082 5593 10094 5596
rect 10036 5587 10094 5593
rect 11698 5584 11704 5596
rect 11756 5584 11762 5636
rect 12406 5624 12434 5664
rect 14458 5652 14464 5704
rect 14516 5692 14522 5704
rect 14645 5695 14703 5701
rect 14645 5692 14657 5695
rect 14516 5664 14657 5692
rect 14516 5652 14522 5664
rect 14645 5661 14657 5664
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 16114 5652 16120 5704
rect 16172 5692 16178 5704
rect 17313 5695 17371 5701
rect 17313 5692 17325 5695
rect 16172 5664 17325 5692
rect 16172 5652 16178 5664
rect 17313 5661 17325 5664
rect 17359 5661 17371 5695
rect 17494 5692 17500 5704
rect 17455 5664 17500 5692
rect 17313 5655 17371 5661
rect 12618 5624 12624 5636
rect 12406 5596 12624 5624
rect 12618 5584 12624 5596
rect 12676 5584 12682 5636
rect 14369 5627 14427 5633
rect 14369 5624 14381 5627
rect 13648 5596 14381 5624
rect 3145 5559 3203 5565
rect 3145 5525 3157 5559
rect 3191 5556 3203 5559
rect 5810 5556 5816 5568
rect 3191 5528 5816 5556
rect 3191 5525 3203 5528
rect 3145 5519 3203 5525
rect 5810 5516 5816 5528
rect 5868 5556 5874 5568
rect 13648 5556 13676 5596
rect 14369 5593 14381 5596
rect 14415 5624 14427 5627
rect 16132 5624 16160 5652
rect 14415 5596 16160 5624
rect 17328 5624 17356 5655
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 19429 5695 19487 5701
rect 19429 5661 19441 5695
rect 19475 5661 19487 5695
rect 19610 5692 19616 5704
rect 19571 5664 19616 5692
rect 19429 5655 19487 5661
rect 18874 5624 18880 5636
rect 17328 5596 18880 5624
rect 14415 5593 14427 5596
rect 14369 5587 14427 5593
rect 18874 5584 18880 5596
rect 18932 5624 18938 5636
rect 19444 5624 19472 5655
rect 19610 5652 19616 5664
rect 19668 5652 19674 5704
rect 18932 5596 19472 5624
rect 18932 5584 18938 5596
rect 5868 5528 13676 5556
rect 5868 5516 5874 5528
rect 13722 5516 13728 5568
rect 13780 5556 13786 5568
rect 14553 5559 14611 5565
rect 14553 5556 14565 5559
rect 13780 5528 14565 5556
rect 13780 5516 13786 5528
rect 14553 5525 14565 5528
rect 14599 5525 14611 5559
rect 14553 5519 14611 5525
rect 15470 5516 15476 5568
rect 15528 5556 15534 5568
rect 16117 5559 16175 5565
rect 16117 5556 16129 5559
rect 15528 5528 16129 5556
rect 15528 5516 15534 5528
rect 16117 5525 16129 5528
rect 16163 5525 16175 5559
rect 16482 5556 16488 5568
rect 16443 5528 16488 5556
rect 16117 5519 16175 5525
rect 16482 5516 16488 5528
rect 16540 5516 16546 5568
rect 16577 5559 16635 5565
rect 16577 5525 16589 5559
rect 16623 5556 16635 5559
rect 17405 5559 17463 5565
rect 17405 5556 17417 5559
rect 16623 5528 17417 5556
rect 16623 5525 16635 5528
rect 16577 5519 16635 5525
rect 17405 5525 17417 5528
rect 17451 5525 17463 5559
rect 17405 5519 17463 5525
rect 1104 5466 21043 5488
rect 1104 5414 5894 5466
rect 5946 5414 5958 5466
rect 6010 5414 6022 5466
rect 6074 5414 6086 5466
rect 6138 5414 6150 5466
rect 6202 5414 10839 5466
rect 10891 5414 10903 5466
rect 10955 5414 10967 5466
rect 11019 5414 11031 5466
rect 11083 5414 11095 5466
rect 11147 5414 15784 5466
rect 15836 5414 15848 5466
rect 15900 5414 15912 5466
rect 15964 5414 15976 5466
rect 16028 5414 16040 5466
rect 16092 5414 20729 5466
rect 20781 5414 20793 5466
rect 20845 5414 20857 5466
rect 20909 5414 20921 5466
rect 20973 5414 20985 5466
rect 21037 5414 21043 5466
rect 1104 5392 21043 5414
rect 7558 5312 7564 5364
rect 7616 5352 7622 5364
rect 17037 5355 17095 5361
rect 7616 5324 15608 5352
rect 7616 5312 7622 5324
rect 1578 5244 1584 5296
rect 1636 5284 1642 5296
rect 10036 5287 10094 5293
rect 1636 5256 4200 5284
rect 1636 5244 1642 5256
rect 4172 5225 4200 5256
rect 4724 5256 6408 5284
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5216 2559 5219
rect 3901 5219 3959 5225
rect 3901 5216 3913 5219
rect 2547 5188 3913 5216
rect 2547 5185 2559 5188
rect 2501 5179 2559 5185
rect 3901 5185 3913 5188
rect 3947 5216 3959 5219
rect 4157 5219 4215 5225
rect 3947 5188 4108 5216
rect 3947 5185 3959 5188
rect 3901 5179 3959 5185
rect 4080 5148 4108 5188
rect 4157 5185 4169 5219
rect 4203 5216 4215 5219
rect 4522 5216 4528 5228
rect 4203 5188 4528 5216
rect 4203 5185 4215 5188
rect 4157 5179 4215 5185
rect 4522 5176 4528 5188
rect 4580 5216 4586 5228
rect 4617 5219 4675 5225
rect 4617 5216 4629 5219
rect 4580 5188 4629 5216
rect 4580 5176 4586 5188
rect 4617 5185 4629 5188
rect 4663 5185 4675 5219
rect 4617 5179 4675 5185
rect 4724 5148 4752 5256
rect 4884 5219 4942 5225
rect 4884 5185 4896 5219
rect 4930 5216 4942 5219
rect 5626 5216 5632 5228
rect 4930 5188 5632 5216
rect 4930 5185 4942 5188
rect 4884 5179 4942 5185
rect 5626 5176 5632 5188
rect 5684 5176 5690 5228
rect 6380 5216 6408 5256
rect 10036 5253 10048 5287
rect 10082 5284 10094 5287
rect 15470 5284 15476 5296
rect 10082 5256 15476 5284
rect 10082 5253 10094 5256
rect 10036 5247 10094 5253
rect 15470 5244 15476 5256
rect 15528 5244 15534 5296
rect 11422 5216 11428 5228
rect 6380 5188 11428 5216
rect 11422 5176 11428 5188
rect 11480 5176 11486 5228
rect 12894 5216 12900 5228
rect 12855 5188 12900 5216
rect 12894 5176 12900 5188
rect 12952 5176 12958 5228
rect 13817 5219 13875 5225
rect 13817 5185 13829 5219
rect 13863 5216 13875 5219
rect 13906 5216 13912 5228
rect 13863 5188 13912 5216
rect 13863 5185 13875 5188
rect 13817 5179 13875 5185
rect 13906 5176 13912 5188
rect 13964 5176 13970 5228
rect 14369 5219 14427 5225
rect 14369 5185 14381 5219
rect 14415 5216 14427 5219
rect 15010 5216 15016 5228
rect 14415 5188 15016 5216
rect 14415 5185 14427 5188
rect 14369 5179 14427 5185
rect 4080 5120 4752 5148
rect 9582 5108 9588 5160
rect 9640 5148 9646 5160
rect 9769 5151 9827 5157
rect 9769 5148 9781 5151
rect 9640 5120 9781 5148
rect 9640 5108 9646 5120
rect 9769 5117 9781 5120
rect 9815 5117 9827 5151
rect 9769 5111 9827 5117
rect 12802 5108 12808 5160
rect 12860 5148 12866 5160
rect 12989 5151 13047 5157
rect 12989 5148 13001 5151
rect 12860 5120 13001 5148
rect 12860 5108 12866 5120
rect 12989 5117 13001 5120
rect 13035 5117 13047 5151
rect 12989 5111 13047 5117
rect 13173 5151 13231 5157
rect 13173 5117 13185 5151
rect 13219 5148 13231 5151
rect 14274 5148 14280 5160
rect 13219 5120 14280 5148
rect 13219 5117 13231 5120
rect 13173 5111 13231 5117
rect 14274 5108 14280 5120
rect 14332 5148 14338 5160
rect 14384 5148 14412 5179
rect 15010 5176 15016 5188
rect 15068 5176 15074 5228
rect 15194 5216 15200 5228
rect 15155 5188 15200 5216
rect 15194 5176 15200 5188
rect 15252 5176 15258 5228
rect 15289 5219 15347 5225
rect 15289 5185 15301 5219
rect 15335 5185 15347 5219
rect 15289 5179 15347 5185
rect 14332 5120 14412 5148
rect 14332 5108 14338 5120
rect 14826 5108 14832 5160
rect 14884 5148 14890 5160
rect 15304 5148 15332 5179
rect 15378 5176 15384 5228
rect 15436 5216 15442 5228
rect 15580 5225 15608 5324
rect 17037 5321 17049 5355
rect 17083 5352 17095 5355
rect 17494 5352 17500 5364
rect 17083 5324 17500 5352
rect 17083 5321 17095 5324
rect 17037 5315 17095 5321
rect 17494 5312 17500 5324
rect 17552 5312 17558 5364
rect 15565 5219 15623 5225
rect 15436 5188 15481 5216
rect 15436 5176 15442 5188
rect 15565 5185 15577 5219
rect 15611 5185 15623 5219
rect 15565 5179 15623 5185
rect 16945 5219 17003 5225
rect 16945 5185 16957 5219
rect 16991 5216 17003 5219
rect 17034 5216 17040 5228
rect 16991 5188 17040 5216
rect 16991 5185 17003 5188
rect 16945 5179 17003 5185
rect 17034 5176 17040 5188
rect 17092 5176 17098 5228
rect 14884 5120 15332 5148
rect 14884 5108 14890 5120
rect 2774 5040 2780 5092
rect 2832 5080 2838 5092
rect 11146 5080 11152 5092
rect 2832 5052 2877 5080
rect 11107 5052 11152 5080
rect 2832 5040 2838 5052
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 11238 5040 11244 5092
rect 11296 5080 11302 5092
rect 14921 5083 14979 5089
rect 14921 5080 14933 5083
rect 11296 5052 11928 5080
rect 11296 5040 11302 5052
rect 5810 4972 5816 5024
rect 5868 5012 5874 5024
rect 5997 5015 6055 5021
rect 5997 5012 6009 5015
rect 5868 4984 6009 5012
rect 5868 4972 5874 4984
rect 5997 4981 6009 4984
rect 6043 4981 6055 5015
rect 11900 5012 11928 5052
rect 14844 5052 14933 5080
rect 12529 5015 12587 5021
rect 12529 5012 12541 5015
rect 11900 4984 12541 5012
rect 5997 4975 6055 4981
rect 12529 4981 12541 4984
rect 12575 4981 12587 5015
rect 12529 4975 12587 4981
rect 12618 4972 12624 5024
rect 12676 5012 12682 5024
rect 14844 5012 14872 5052
rect 14921 5049 14933 5052
rect 14967 5049 14979 5083
rect 14921 5043 14979 5049
rect 12676 4984 14872 5012
rect 12676 4972 12682 4984
rect 1104 4922 20884 4944
rect 1104 4870 3422 4922
rect 3474 4870 3486 4922
rect 3538 4870 3550 4922
rect 3602 4870 3614 4922
rect 3666 4870 3678 4922
rect 3730 4870 8367 4922
rect 8419 4870 8431 4922
rect 8483 4870 8495 4922
rect 8547 4870 8559 4922
rect 8611 4870 8623 4922
rect 8675 4870 13312 4922
rect 13364 4870 13376 4922
rect 13428 4870 13440 4922
rect 13492 4870 13504 4922
rect 13556 4870 13568 4922
rect 13620 4870 18257 4922
rect 18309 4870 18321 4922
rect 18373 4870 18385 4922
rect 18437 4870 18449 4922
rect 18501 4870 18513 4922
rect 18565 4870 20884 4922
rect 1104 4848 20884 4870
rect 12618 4808 12624 4820
rect 8956 4780 12624 4808
rect 1578 4632 1584 4684
rect 1636 4672 1642 4684
rect 2041 4675 2099 4681
rect 2041 4672 2053 4675
rect 1636 4644 2053 4672
rect 1636 4632 1642 4644
rect 2041 4641 2053 4644
rect 2087 4641 2099 4675
rect 2041 4635 2099 4641
rect 4522 4632 4528 4684
rect 4580 4672 4586 4684
rect 5261 4675 5319 4681
rect 5261 4672 5273 4675
rect 4580 4644 5273 4672
rect 4580 4632 4586 4644
rect 5261 4641 5273 4644
rect 5307 4641 5319 4675
rect 7098 4672 7104 4684
rect 7059 4644 7104 4672
rect 5261 4635 5319 4641
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 5528 4607 5586 4613
rect 5528 4573 5540 4607
rect 5574 4604 5586 4607
rect 8956 4604 8984 4780
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 14642 4768 14648 4820
rect 14700 4808 14706 4820
rect 15378 4808 15384 4820
rect 14700 4780 15384 4808
rect 14700 4768 14706 4780
rect 15378 4768 15384 4780
rect 15436 4768 15442 4820
rect 14918 4740 14924 4752
rect 10888 4712 14924 4740
rect 5574 4576 8984 4604
rect 5574 4573 5586 4576
rect 5528 4567 5586 4573
rect 9582 4564 9588 4616
rect 9640 4604 9646 4616
rect 9769 4607 9827 4613
rect 9769 4604 9781 4607
rect 9640 4576 9781 4604
rect 9640 4564 9646 4576
rect 9769 4573 9781 4576
rect 9815 4573 9827 4607
rect 9769 4567 9827 4573
rect 10036 4607 10094 4613
rect 10036 4573 10048 4607
rect 10082 4604 10094 4607
rect 10888 4604 10916 4712
rect 14918 4700 14924 4712
rect 14976 4700 14982 4752
rect 15102 4700 15108 4752
rect 15160 4740 15166 4752
rect 16945 4743 17003 4749
rect 16945 4740 16957 4743
rect 15160 4712 16957 4740
rect 15160 4700 15166 4712
rect 16945 4709 16957 4712
rect 16991 4709 17003 4743
rect 19610 4740 19616 4752
rect 16945 4703 17003 4709
rect 17052 4712 19616 4740
rect 15194 4632 15200 4684
rect 15252 4672 15258 4684
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 15252 4644 15669 4672
rect 15252 4632 15258 4644
rect 15657 4641 15669 4644
rect 15703 4641 15715 4675
rect 17052 4672 17080 4712
rect 19610 4700 19616 4712
rect 19668 4700 19674 4752
rect 15657 4635 15715 4641
rect 16592 4644 17080 4672
rect 17129 4675 17187 4681
rect 10082 4576 10916 4604
rect 10082 4573 10094 4576
rect 10036 4567 10094 4573
rect 12802 4564 12808 4616
rect 12860 4604 12866 4616
rect 13541 4607 13599 4613
rect 13541 4604 13553 4607
rect 12860 4576 13553 4604
rect 12860 4564 12866 4576
rect 13541 4573 13553 4576
rect 13587 4573 13599 4607
rect 13541 4567 13599 4573
rect 13633 4607 13691 4613
rect 13633 4573 13645 4607
rect 13679 4604 13691 4607
rect 14461 4607 14519 4613
rect 14461 4604 14473 4607
rect 13679 4576 14473 4604
rect 13679 4573 13691 4576
rect 13633 4567 13691 4573
rect 14461 4573 14473 4576
rect 14507 4573 14519 4607
rect 14642 4604 14648 4616
rect 14603 4576 14648 4604
rect 14461 4567 14519 4573
rect 14642 4564 14648 4576
rect 14700 4564 14706 4616
rect 14863 4607 14921 4613
rect 14738 4585 14796 4591
rect 14738 4551 14750 4585
rect 14784 4551 14796 4585
rect 14863 4573 14875 4607
rect 14909 4604 14921 4607
rect 15212 4604 15240 4632
rect 14909 4576 15240 4604
rect 14909 4573 14921 4576
rect 14863 4567 14921 4573
rect 15378 4564 15384 4616
rect 15436 4604 15442 4616
rect 15565 4607 15623 4613
rect 15565 4604 15577 4607
rect 15436 4576 15577 4604
rect 15436 4564 15442 4576
rect 15565 4573 15577 4576
rect 15611 4573 15623 4607
rect 15565 4567 15623 4573
rect 14738 4548 14796 4551
rect 2308 4539 2366 4545
rect 2308 4505 2320 4539
rect 2354 4536 2366 4539
rect 3970 4536 3976 4548
rect 2354 4508 3976 4536
rect 2354 4505 2366 4508
rect 2308 4499 2366 4505
rect 3970 4496 3976 4508
rect 4028 4496 4034 4548
rect 7368 4539 7426 4545
rect 7368 4505 7380 4539
rect 7414 4536 7426 4539
rect 9858 4536 9864 4548
rect 7414 4508 9864 4536
rect 7414 4505 7426 4508
rect 7368 4499 7426 4505
rect 9858 4496 9864 4508
rect 9916 4496 9922 4548
rect 14734 4496 14740 4548
rect 14792 4496 14798 4548
rect 15105 4539 15163 4545
rect 15105 4505 15117 4539
rect 15151 4536 15163 4539
rect 16592 4536 16620 4644
rect 17129 4641 17141 4675
rect 17175 4672 17187 4675
rect 17494 4672 17500 4684
rect 17175 4644 17500 4672
rect 17175 4641 17187 4644
rect 17129 4635 17187 4641
rect 17494 4632 17500 4644
rect 17552 4632 17558 4684
rect 16666 4564 16672 4616
rect 16724 4604 16730 4616
rect 17218 4604 17224 4616
rect 16724 4576 17224 4604
rect 16724 4564 16730 4576
rect 17218 4564 17224 4576
rect 17276 4564 17282 4616
rect 18046 4604 18052 4616
rect 18007 4576 18052 4604
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 15151 4508 16620 4536
rect 15151 4505 15163 4508
rect 15105 4499 15163 4505
rect 16850 4496 16856 4548
rect 16908 4536 16914 4548
rect 17497 4539 17555 4545
rect 17497 4536 17509 4539
rect 16908 4508 17509 4536
rect 16908 4496 16914 4508
rect 17497 4505 17509 4508
rect 17543 4505 17555 4539
rect 17497 4499 17555 4505
rect 17589 4539 17647 4545
rect 17589 4505 17601 4539
rect 17635 4536 17647 4539
rect 18141 4539 18199 4545
rect 18141 4536 18153 4539
rect 17635 4508 18153 4536
rect 17635 4505 17647 4508
rect 17589 4499 17647 4505
rect 18141 4505 18153 4508
rect 18187 4505 18199 4539
rect 18141 4499 18199 4505
rect 3421 4471 3479 4477
rect 3421 4437 3433 4471
rect 3467 4468 3479 4471
rect 4798 4468 4804 4480
rect 3467 4440 4804 4468
rect 3467 4437 3479 4440
rect 3421 4431 3479 4437
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 6638 4468 6644 4480
rect 6599 4440 6644 4468
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 8481 4471 8539 4477
rect 8481 4437 8493 4471
rect 8527 4468 8539 4471
rect 10410 4468 10416 4480
rect 8527 4440 10416 4468
rect 8527 4437 8539 4440
rect 8481 4431 8539 4437
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 11149 4471 11207 4477
rect 11149 4437 11161 4471
rect 11195 4468 11207 4471
rect 17126 4468 17132 4480
rect 11195 4440 17132 4468
rect 11195 4437 11207 4440
rect 11149 4431 11207 4437
rect 17126 4428 17132 4440
rect 17184 4428 17190 4480
rect 1104 4378 21043 4400
rect 1104 4326 5894 4378
rect 5946 4326 5958 4378
rect 6010 4326 6022 4378
rect 6074 4326 6086 4378
rect 6138 4326 6150 4378
rect 6202 4326 10839 4378
rect 10891 4326 10903 4378
rect 10955 4326 10967 4378
rect 11019 4326 11031 4378
rect 11083 4326 11095 4378
rect 11147 4326 15784 4378
rect 15836 4326 15848 4378
rect 15900 4326 15912 4378
rect 15964 4326 15976 4378
rect 16028 4326 16040 4378
rect 16092 4326 20729 4378
rect 20781 4326 20793 4378
rect 20845 4326 20857 4378
rect 20909 4326 20921 4378
rect 20973 4326 20985 4378
rect 21037 4326 21043 4378
rect 1104 4304 21043 4326
rect 9858 4224 9864 4276
rect 9916 4264 9922 4276
rect 12986 4264 12992 4276
rect 9916 4236 12992 4264
rect 9916 4224 9922 4236
rect 12986 4224 12992 4236
rect 13044 4224 13050 4276
rect 16942 4224 16948 4276
rect 17000 4264 17006 4276
rect 17037 4267 17095 4273
rect 17037 4264 17049 4267
rect 17000 4236 17049 4264
rect 17000 4224 17006 4236
rect 17037 4233 17049 4236
rect 17083 4233 17095 4267
rect 17037 4227 17095 4233
rect 6638 4156 6644 4208
rect 6696 4196 6702 4208
rect 12894 4196 12900 4208
rect 6696 4168 12900 4196
rect 6696 4156 6702 4168
rect 12894 4156 12900 4168
rect 12952 4196 12958 4208
rect 13722 4196 13728 4208
rect 12952 4168 13728 4196
rect 12952 4156 12958 4168
rect 13722 4156 13728 4168
rect 13780 4196 13786 4208
rect 13780 4168 14504 4196
rect 13780 4156 13786 4168
rect 1578 4128 1584 4140
rect 1539 4100 1584 4128
rect 1578 4088 1584 4100
rect 1636 4088 1642 4140
rect 1854 4137 1860 4140
rect 1848 4091 1860 4137
rect 1912 4128 1918 4140
rect 4522 4128 4528 4140
rect 1912 4100 1948 4128
rect 4483 4100 4528 4128
rect 1854 4088 1860 4091
rect 1912 4088 1918 4100
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 4792 4131 4850 4137
rect 4792 4097 4804 4131
rect 4838 4128 4850 4131
rect 7098 4128 7104 4140
rect 4838 4100 6960 4128
rect 7059 4100 7104 4128
rect 4838 4097 4850 4100
rect 4792 4091 4850 4097
rect 6932 4060 6960 4100
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 7368 4131 7426 4137
rect 7368 4097 7380 4131
rect 7414 4128 7426 4131
rect 9674 4128 9680 4140
rect 7414 4100 9680 4128
rect 7414 4097 7426 4100
rect 7368 4091 7426 4097
rect 9674 4088 9680 4100
rect 9732 4088 9738 4140
rect 9852 4131 9910 4137
rect 9852 4097 9864 4131
rect 9898 4128 9910 4131
rect 11698 4128 11704 4140
rect 9898 4100 11704 4128
rect 9898 4097 9910 4100
rect 9852 4091 9910 4097
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 14185 4131 14243 4137
rect 14185 4097 14197 4131
rect 14231 4097 14243 4131
rect 14185 4091 14243 4097
rect 14369 4131 14427 4137
rect 14369 4097 14381 4131
rect 14415 4097 14427 4131
rect 14476 4128 14504 4168
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14476 4100 14657 4128
rect 14369 4091 14427 4097
rect 14645 4097 14657 4100
rect 14691 4097 14703 4131
rect 14826 4128 14832 4140
rect 14787 4100 14832 4128
rect 14645 4091 14703 4097
rect 7006 4060 7012 4072
rect 6932 4032 7012 4060
rect 7006 4020 7012 4032
rect 7064 4020 7070 4072
rect 9582 4060 9588 4072
rect 9543 4032 9588 4060
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 14200 3992 14228 4091
rect 14384 4060 14412 4091
rect 14826 4088 14832 4100
rect 14884 4088 14890 4140
rect 15010 4128 15016 4140
rect 14971 4100 15016 4128
rect 15010 4088 15016 4100
rect 15068 4088 15074 4140
rect 16850 4128 16856 4140
rect 16811 4100 16856 4128
rect 16850 4088 16856 4100
rect 16908 4088 16914 4140
rect 17126 4088 17132 4140
rect 17184 4128 17190 4140
rect 17221 4131 17279 4137
rect 17221 4128 17233 4131
rect 17184 4100 17233 4128
rect 17184 4088 17190 4100
rect 17221 4097 17233 4100
rect 17267 4097 17279 4131
rect 17221 4091 17279 4097
rect 17405 4131 17463 4137
rect 17405 4097 17417 4131
rect 17451 4097 17463 4131
rect 17405 4091 17463 4097
rect 14550 4060 14556 4072
rect 14384 4032 14556 4060
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 17310 4060 17316 4072
rect 16408 4032 17316 4060
rect 14918 3992 14924 4004
rect 10888 3964 12434 3992
rect 14200 3964 14924 3992
rect 1946 3884 1952 3936
rect 2004 3924 2010 3936
rect 2961 3927 3019 3933
rect 2961 3924 2973 3927
rect 2004 3896 2973 3924
rect 2004 3884 2010 3896
rect 2961 3893 2973 3896
rect 3007 3893 3019 3927
rect 2961 3887 3019 3893
rect 5905 3927 5963 3933
rect 5905 3893 5917 3927
rect 5951 3924 5963 3927
rect 8202 3924 8208 3936
rect 5951 3896 8208 3924
rect 5951 3893 5963 3896
rect 5905 3887 5963 3893
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8481 3927 8539 3933
rect 8481 3893 8493 3927
rect 8527 3924 8539 3927
rect 10888 3924 10916 3964
rect 8527 3896 10916 3924
rect 10965 3927 11023 3933
rect 8527 3893 8539 3896
rect 8481 3887 8539 3893
rect 10965 3893 10977 3927
rect 11011 3924 11023 3927
rect 11790 3924 11796 3936
rect 11011 3896 11796 3924
rect 11011 3893 11023 3896
rect 10965 3887 11023 3893
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 12406 3924 12434 3964
rect 14918 3952 14924 3964
rect 14976 3952 14982 4004
rect 16408 3924 16436 4032
rect 17310 4020 17316 4032
rect 17368 4060 17374 4072
rect 17420 4060 17448 4091
rect 17368 4032 17448 4060
rect 17368 4020 17374 4032
rect 12406 3896 16436 3924
rect 16482 3884 16488 3936
rect 16540 3924 16546 3936
rect 17034 3924 17040 3936
rect 16540 3896 17040 3924
rect 16540 3884 16546 3896
rect 17034 3884 17040 3896
rect 17092 3924 17098 3936
rect 17221 3927 17279 3933
rect 17221 3924 17233 3927
rect 17092 3896 17233 3924
rect 17092 3884 17098 3896
rect 17221 3893 17233 3896
rect 17267 3893 17279 3927
rect 17221 3887 17279 3893
rect 1104 3834 20884 3856
rect 1104 3782 3422 3834
rect 3474 3782 3486 3834
rect 3538 3782 3550 3834
rect 3602 3782 3614 3834
rect 3666 3782 3678 3834
rect 3730 3782 8367 3834
rect 8419 3782 8431 3834
rect 8483 3782 8495 3834
rect 8547 3782 8559 3834
rect 8611 3782 8623 3834
rect 8675 3782 13312 3834
rect 13364 3782 13376 3834
rect 13428 3782 13440 3834
rect 13492 3782 13504 3834
rect 13556 3782 13568 3834
rect 13620 3782 18257 3834
rect 18309 3782 18321 3834
rect 18373 3782 18385 3834
rect 18437 3782 18449 3834
rect 18501 3782 18513 3834
rect 18565 3782 20884 3834
rect 1104 3760 20884 3782
rect 3142 3680 3148 3732
rect 3200 3720 3206 3732
rect 5534 3720 5540 3732
rect 3200 3692 5540 3720
rect 3200 3680 3206 3692
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 12986 3720 12992 3732
rect 9732 3692 12434 3720
rect 12947 3692 12992 3720
rect 9732 3680 9738 3692
rect 11057 3655 11115 3661
rect 11057 3621 11069 3655
rect 11103 3621 11115 3655
rect 11057 3615 11115 3621
rect 11793 3655 11851 3661
rect 11793 3621 11805 3655
rect 11839 3652 11851 3655
rect 11882 3652 11888 3664
rect 11839 3624 11888 3652
rect 11839 3621 11851 3624
rect 11793 3615 11851 3621
rect 1578 3544 1584 3596
rect 1636 3584 1642 3596
rect 2041 3587 2099 3593
rect 2041 3584 2053 3587
rect 1636 3556 2053 3584
rect 1636 3544 1642 3556
rect 2041 3553 2053 3556
rect 2087 3553 2099 3587
rect 2041 3547 2099 3553
rect 8202 3544 8208 3596
rect 8260 3584 8266 3596
rect 11072 3584 11100 3615
rect 11882 3612 11888 3624
rect 11940 3612 11946 3664
rect 12406 3652 12434 3692
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 14277 3723 14335 3729
rect 14277 3689 14289 3723
rect 14323 3720 14335 3723
rect 14642 3720 14648 3732
rect 14323 3692 14648 3720
rect 14323 3689 14335 3692
rect 14277 3683 14335 3689
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 17218 3720 17224 3732
rect 17179 3692 17224 3720
rect 17218 3680 17224 3692
rect 17276 3720 17282 3732
rect 18233 3723 18291 3729
rect 18233 3720 18245 3723
rect 17276 3692 18245 3720
rect 17276 3680 17282 3692
rect 18233 3689 18245 3692
rect 18279 3689 18291 3723
rect 18233 3683 18291 3689
rect 16761 3655 16819 3661
rect 16761 3652 16773 3655
rect 12406 3624 16773 3652
rect 16761 3621 16773 3624
rect 16807 3621 16819 3655
rect 16761 3615 16819 3621
rect 12802 3584 12808 3596
rect 8260 3556 9812 3584
rect 11072 3556 12808 3584
rect 8260 3544 8266 3556
rect 7009 3519 7067 3525
rect 7009 3485 7021 3519
rect 7055 3516 7067 3519
rect 7098 3516 7104 3528
rect 7055 3488 7104 3516
rect 7055 3485 7067 3488
rect 7009 3479 7067 3485
rect 7098 3476 7104 3488
rect 7156 3516 7162 3528
rect 9582 3516 9588 3528
rect 7156 3488 9588 3516
rect 7156 3476 7162 3488
rect 9582 3476 9588 3488
rect 9640 3516 9646 3528
rect 9677 3519 9735 3525
rect 9677 3516 9689 3519
rect 9640 3488 9689 3516
rect 9640 3476 9646 3488
rect 9677 3485 9689 3488
rect 9723 3485 9735 3519
rect 9784 3516 9812 3556
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 13449 3587 13507 3593
rect 13449 3584 13461 3587
rect 13096 3556 13461 3584
rect 9944 3519 10002 3525
rect 9784 3488 9895 3516
rect 9677 3479 9735 3485
rect 2308 3451 2366 3457
rect 2308 3417 2320 3451
rect 2354 3448 2366 3451
rect 2958 3448 2964 3460
rect 2354 3420 2964 3448
rect 2354 3417 2366 3420
rect 2308 3411 2366 3417
rect 2958 3408 2964 3420
rect 3016 3408 3022 3460
rect 7276 3451 7334 3457
rect 7276 3417 7288 3451
rect 7322 3448 7334 3451
rect 9766 3448 9772 3460
rect 7322 3420 9772 3448
rect 7322 3417 7334 3420
rect 7276 3411 7334 3417
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 3326 3340 3332 3392
rect 3384 3380 3390 3392
rect 3421 3383 3479 3389
rect 3421 3380 3433 3383
rect 3384 3352 3433 3380
rect 3384 3340 3390 3352
rect 3421 3349 3433 3352
rect 3467 3349 3479 3383
rect 3421 3343 3479 3349
rect 4798 3340 4804 3392
rect 4856 3380 4862 3392
rect 6730 3380 6736 3392
rect 4856 3352 6736 3380
rect 4856 3340 4862 3352
rect 6730 3340 6736 3352
rect 6788 3340 6794 3392
rect 8389 3383 8447 3389
rect 8389 3349 8401 3383
rect 8435 3380 8447 3383
rect 8754 3380 8760 3392
rect 8435 3352 8760 3380
rect 8435 3349 8447 3352
rect 8389 3343 8447 3349
rect 8754 3340 8760 3352
rect 8812 3340 8818 3392
rect 9867 3380 9895 3488
rect 9944 3485 9956 3519
rect 9990 3516 10002 3519
rect 11238 3516 11244 3528
rect 9990 3488 11244 3516
rect 9990 3485 10002 3488
rect 9944 3479 10002 3485
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 11790 3516 11796 3528
rect 11751 3488 11796 3516
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 11974 3516 11980 3528
rect 11935 3488 11980 3516
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 12066 3476 12072 3528
rect 12124 3516 12130 3528
rect 13096 3516 13124 3556
rect 13449 3553 13461 3556
rect 13495 3584 13507 3587
rect 14553 3587 14611 3593
rect 14553 3584 14565 3587
rect 13495 3556 14565 3584
rect 13495 3553 13507 3556
rect 13449 3547 13507 3553
rect 14553 3553 14565 3556
rect 14599 3584 14611 3587
rect 15010 3584 15016 3596
rect 14599 3556 15016 3584
rect 14599 3553 14611 3556
rect 14553 3547 14611 3553
rect 15010 3544 15016 3556
rect 15068 3544 15074 3596
rect 16960 3556 18000 3584
rect 12124 3488 12169 3516
rect 13004 3488 13124 3516
rect 13173 3519 13231 3525
rect 12124 3476 12130 3488
rect 10410 3408 10416 3460
rect 10468 3448 10474 3460
rect 13004 3448 13032 3488
rect 13173 3485 13185 3519
rect 13219 3485 13231 3519
rect 13354 3516 13360 3528
rect 13315 3488 13360 3516
rect 13173 3479 13231 3485
rect 10468 3420 13032 3448
rect 13188 3448 13216 3479
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 13722 3476 13728 3528
rect 13780 3516 13786 3528
rect 14461 3519 14519 3525
rect 14461 3516 14473 3519
rect 13780 3488 14473 3516
rect 13780 3476 13786 3488
rect 14461 3485 14473 3488
rect 14507 3485 14519 3519
rect 14918 3516 14924 3528
rect 14831 3488 14924 3516
rect 14461 3479 14519 3485
rect 14918 3476 14924 3488
rect 14976 3516 14982 3528
rect 16298 3516 16304 3528
rect 14976 3488 16304 3516
rect 14976 3476 14982 3488
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 16960 3525 16988 3556
rect 17972 3528 18000 3556
rect 16945 3519 17003 3525
rect 16945 3485 16957 3519
rect 16991 3485 17003 3519
rect 16945 3479 17003 3485
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17310 3516 17316 3528
rect 17092 3488 17137 3516
rect 17271 3488 17316 3516
rect 17092 3476 17098 3488
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 17954 3516 17960 3528
rect 17915 3488 17960 3516
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 18046 3476 18052 3528
rect 18104 3516 18110 3528
rect 18325 3519 18383 3525
rect 18104 3488 18149 3516
rect 18104 3476 18110 3488
rect 18325 3485 18337 3519
rect 18371 3485 18383 3519
rect 18325 3479 18383 3485
rect 14182 3448 14188 3460
rect 13188 3420 14188 3448
rect 10468 3408 10474 3420
rect 14182 3408 14188 3420
rect 14240 3408 14246 3460
rect 14550 3408 14556 3460
rect 14608 3448 14614 3460
rect 14829 3451 14887 3457
rect 14829 3448 14841 3451
rect 14608 3420 14841 3448
rect 14608 3408 14614 3420
rect 14829 3417 14841 3420
rect 14875 3417 14887 3451
rect 14829 3411 14887 3417
rect 16850 3408 16856 3460
rect 16908 3448 16914 3460
rect 18340 3448 18368 3479
rect 16908 3420 18368 3448
rect 16908 3408 16914 3420
rect 14645 3383 14703 3389
rect 14645 3380 14657 3383
rect 9867 3352 14657 3380
rect 14645 3349 14657 3352
rect 14691 3380 14703 3383
rect 15378 3380 15384 3392
rect 14691 3352 15384 3380
rect 14691 3349 14703 3352
rect 14645 3343 14703 3349
rect 15378 3340 15384 3352
rect 15436 3340 15442 3392
rect 17770 3380 17776 3392
rect 17731 3352 17776 3380
rect 17770 3340 17776 3352
rect 17828 3340 17834 3392
rect 1104 3290 21043 3312
rect 1104 3238 5894 3290
rect 5946 3238 5958 3290
rect 6010 3238 6022 3290
rect 6074 3238 6086 3290
rect 6138 3238 6150 3290
rect 6202 3238 10839 3290
rect 10891 3238 10903 3290
rect 10955 3238 10967 3290
rect 11019 3238 11031 3290
rect 11083 3238 11095 3290
rect 11147 3238 15784 3290
rect 15836 3238 15848 3290
rect 15900 3238 15912 3290
rect 15964 3238 15976 3290
rect 16028 3238 16040 3290
rect 16092 3238 20729 3290
rect 20781 3238 20793 3290
rect 20845 3238 20857 3290
rect 20909 3238 20921 3290
rect 20973 3238 20985 3290
rect 21037 3238 21043 3290
rect 1104 3216 21043 3238
rect 1854 3176 1860 3188
rect 1815 3148 1860 3176
rect 1854 3136 1860 3148
rect 1912 3136 1918 3188
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 5537 3179 5595 3185
rect 3384 3148 5028 3176
rect 3384 3136 3390 3148
rect 2590 3108 2596 3120
rect 2551 3080 2596 3108
rect 2590 3068 2596 3080
rect 2648 3068 2654 3120
rect 4341 3111 4399 3117
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 4522 3108 4528 3120
rect 4387 3080 4528 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 4522 3068 4528 3080
rect 4580 3068 4586 3120
rect 4798 3108 4804 3120
rect 4759 3080 4804 3108
rect 4798 3068 4804 3080
rect 4856 3068 4862 3120
rect 5000 3108 5028 3148
rect 5537 3145 5549 3179
rect 5583 3176 5595 3179
rect 5626 3176 5632 3188
rect 5583 3148 5632 3176
rect 5583 3145 5595 3148
rect 5537 3139 5595 3145
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 7650 3176 7656 3188
rect 5736 3148 7656 3176
rect 5000 3080 5120 3108
rect 1765 3043 1823 3049
rect 1765 3009 1777 3043
rect 1811 3009 1823 3043
rect 1946 3040 1952 3052
rect 1907 3012 1952 3040
rect 1765 3003 1823 3009
rect 1780 2972 1808 3003
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 2314 2972 2320 2984
rect 1780 2944 2320 2972
rect 2314 2932 2320 2944
rect 2372 2932 2378 2984
rect 4816 2904 4844 3068
rect 5092 3049 5120 3080
rect 4985 3043 5043 3049
rect 4985 3009 4997 3043
rect 5031 3009 5043 3043
rect 4985 3003 5043 3009
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3040 5135 3043
rect 5626 3040 5632 3052
rect 5123 3012 5632 3040
rect 5123 3009 5135 3012
rect 5077 3003 5135 3009
rect 4890 2932 4896 2984
rect 4948 2972 4954 2984
rect 5000 2972 5028 3003
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 5736 3049 5764 3148
rect 7650 3136 7656 3148
rect 7708 3136 7714 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 10045 3179 10103 3185
rect 10045 3176 10057 3179
rect 9824 3148 10057 3176
rect 9824 3136 9830 3148
rect 10045 3145 10057 3148
rect 10091 3145 10103 3179
rect 10045 3139 10103 3145
rect 13354 3136 13360 3188
rect 13412 3176 13418 3188
rect 13630 3176 13636 3188
rect 13412 3148 13636 3176
rect 13412 3136 13418 3148
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 14182 3176 14188 3188
rect 14143 3148 14188 3176
rect 14182 3136 14188 3148
rect 14240 3136 14246 3188
rect 16209 3179 16267 3185
rect 16209 3176 16221 3179
rect 15212 3148 16221 3176
rect 6825 3111 6883 3117
rect 6825 3108 6837 3111
rect 6012 3080 6837 3108
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3009 5779 3043
rect 5721 3003 5779 3009
rect 5810 3000 5816 3052
rect 5868 3040 5874 3052
rect 6012 3049 6040 3080
rect 6825 3077 6837 3080
rect 6871 3077 6883 3111
rect 6825 3071 6883 3077
rect 6917 3111 6975 3117
rect 6917 3077 6929 3111
rect 6963 3077 6975 3111
rect 7834 3108 7840 3120
rect 7795 3080 7840 3108
rect 6917 3071 6975 3077
rect 5997 3043 6055 3049
rect 5997 3040 6009 3043
rect 5868 3012 6009 3040
rect 5868 3000 5874 3012
rect 5997 3009 6009 3012
rect 6043 3009 6055 3043
rect 6730 3040 6736 3052
rect 6691 3012 6736 3040
rect 5997 3003 6055 3009
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 6549 2975 6607 2981
rect 6549 2972 6561 2975
rect 4948 2944 6561 2972
rect 4948 2932 4954 2944
rect 6549 2941 6561 2944
rect 6595 2941 6607 2975
rect 6549 2935 6607 2941
rect 4816 2876 5672 2904
rect 5644 2848 5672 2876
rect 5718 2864 5724 2916
rect 5776 2904 5782 2916
rect 6932 2904 6960 3071
rect 7834 3068 7840 3080
rect 7892 3068 7898 3120
rect 9582 3108 9588 3120
rect 9543 3080 9588 3108
rect 9582 3068 9588 3080
rect 9640 3068 9646 3120
rect 12066 3068 12072 3120
rect 12124 3108 12130 3120
rect 15212 3108 15240 3148
rect 16209 3145 16221 3148
rect 16255 3145 16267 3179
rect 16209 3139 16267 3145
rect 12124 3080 12664 3108
rect 12124 3068 12130 3080
rect 10226 3040 10232 3052
rect 10187 3012 10232 3040
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 12529 3043 12587 3049
rect 12529 3040 12541 3043
rect 11848 3012 12541 3040
rect 11848 3000 11854 3012
rect 12529 3009 12541 3012
rect 12575 3009 12587 3043
rect 12529 3003 12587 3009
rect 7282 2972 7288 2984
rect 7243 2944 7288 2972
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 8754 2932 8760 2984
rect 8812 2972 8818 2984
rect 10505 2975 10563 2981
rect 10505 2972 10517 2975
rect 8812 2944 10517 2972
rect 8812 2932 8818 2944
rect 10505 2941 10517 2944
rect 10551 2972 10563 2975
rect 11974 2972 11980 2984
rect 10551 2944 11980 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 11974 2932 11980 2944
rect 12032 2972 12038 2984
rect 12345 2975 12403 2981
rect 12345 2972 12357 2975
rect 12032 2944 12357 2972
rect 12032 2932 12038 2944
rect 12345 2941 12357 2944
rect 12391 2941 12403 2975
rect 12636 2972 12664 3080
rect 14108 3080 15240 3108
rect 14108 3049 14136 3080
rect 12713 3043 12771 3049
rect 12713 3009 12725 3043
rect 12759 3040 12771 3043
rect 13449 3043 13507 3049
rect 13449 3040 13461 3043
rect 12759 3012 13461 3040
rect 12759 3009 12771 3012
rect 12713 3003 12771 3009
rect 13449 3009 13461 3012
rect 13495 3009 13507 3043
rect 13449 3003 13507 3009
rect 14093 3043 14151 3049
rect 14093 3009 14105 3043
rect 14139 3009 14151 3043
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 14093 3003 14151 3009
rect 13265 2975 13323 2981
rect 13265 2972 13277 2975
rect 12636 2944 13277 2972
rect 12345 2935 12403 2941
rect 13265 2941 13277 2944
rect 13311 2972 13323 2975
rect 13464 2972 13492 3003
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 14918 3040 14924 3052
rect 14879 3012 14924 3040
rect 14918 3000 14924 3012
rect 14976 3000 14982 3052
rect 15212 3049 15240 3080
rect 15841 3111 15899 3117
rect 15841 3077 15853 3111
rect 15887 3077 15899 3111
rect 15841 3071 15899 3077
rect 16057 3111 16115 3117
rect 16057 3077 16069 3111
rect 16103 3108 16115 3111
rect 16298 3108 16304 3120
rect 16103 3080 16304 3108
rect 16103 3077 16115 3080
rect 16057 3071 16115 3077
rect 15197 3043 15255 3049
rect 15197 3009 15209 3043
rect 15243 3040 15255 3043
rect 15286 3040 15292 3052
rect 15243 3012 15292 3040
rect 15243 3009 15255 3012
rect 15197 3003 15255 3009
rect 15286 3000 15292 3012
rect 15344 3000 15350 3052
rect 15378 3000 15384 3052
rect 15436 3040 15442 3052
rect 15436 3012 15481 3040
rect 15436 3000 15442 3012
rect 14826 2972 14832 2984
rect 13311 2944 13400 2972
rect 13464 2944 14832 2972
rect 13311 2941 13323 2944
rect 13265 2935 13323 2941
rect 5776 2876 6960 2904
rect 5776 2864 5782 2876
rect 7006 2864 7012 2916
rect 7064 2904 7070 2916
rect 13170 2904 13176 2916
rect 7064 2876 13176 2904
rect 7064 2864 7070 2876
rect 13170 2864 13176 2876
rect 13228 2864 13234 2916
rect 4798 2836 4804 2848
rect 4759 2808 4804 2836
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 5626 2796 5632 2848
rect 5684 2796 5690 2848
rect 5902 2836 5908 2848
rect 5863 2808 5908 2836
rect 5902 2796 5908 2808
rect 5960 2796 5966 2848
rect 8846 2796 8852 2848
rect 8904 2836 8910 2848
rect 10413 2839 10471 2845
rect 10413 2836 10425 2839
rect 8904 2808 10425 2836
rect 8904 2796 8910 2808
rect 10413 2805 10425 2808
rect 10459 2836 10471 2839
rect 12066 2836 12072 2848
rect 10459 2808 12072 2836
rect 10459 2805 10471 2808
rect 10413 2799 10471 2805
rect 12066 2796 12072 2808
rect 12124 2796 12130 2848
rect 13372 2836 13400 2944
rect 14826 2932 14832 2944
rect 14884 2932 14890 2984
rect 15010 2932 15016 2984
rect 15068 2972 15074 2984
rect 15856 2972 15884 3071
rect 16298 3068 16304 3080
rect 16356 3068 16362 3120
rect 17034 3040 17040 3052
rect 16995 3012 17040 3040
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 15068 2944 15884 2972
rect 17129 2975 17187 2981
rect 15068 2932 15074 2944
rect 17129 2941 17141 2975
rect 17175 2972 17187 2975
rect 17310 2972 17316 2984
rect 17175 2944 17316 2972
rect 17175 2941 17187 2944
rect 17129 2935 17187 2941
rect 17310 2932 17316 2944
rect 17368 2932 17374 2984
rect 17405 2975 17463 2981
rect 17405 2941 17417 2975
rect 17451 2972 17463 2975
rect 18046 2972 18052 2984
rect 17451 2944 18052 2972
rect 17451 2941 17463 2944
rect 17405 2935 17463 2941
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 13446 2864 13452 2916
rect 13504 2904 13510 2916
rect 14737 2907 14795 2913
rect 14737 2904 14749 2907
rect 13504 2876 14749 2904
rect 13504 2864 13510 2876
rect 14737 2873 14749 2876
rect 14783 2873 14795 2907
rect 14737 2867 14795 2873
rect 14550 2836 14556 2848
rect 13372 2808 14556 2836
rect 14550 2796 14556 2808
rect 14608 2836 14614 2848
rect 16025 2839 16083 2845
rect 16025 2836 16037 2839
rect 14608 2808 16037 2836
rect 14608 2796 14614 2808
rect 16025 2805 16037 2808
rect 16071 2805 16083 2839
rect 16025 2799 16083 2805
rect 1104 2746 20884 2768
rect 1104 2694 3422 2746
rect 3474 2694 3486 2746
rect 3538 2694 3550 2746
rect 3602 2694 3614 2746
rect 3666 2694 3678 2746
rect 3730 2694 8367 2746
rect 8419 2694 8431 2746
rect 8483 2694 8495 2746
rect 8547 2694 8559 2746
rect 8611 2694 8623 2746
rect 8675 2694 13312 2746
rect 13364 2694 13376 2746
rect 13428 2694 13440 2746
rect 13492 2694 13504 2746
rect 13556 2694 13568 2746
rect 13620 2694 18257 2746
rect 18309 2694 18321 2746
rect 18373 2694 18385 2746
rect 18437 2694 18449 2746
rect 18501 2694 18513 2746
rect 18565 2694 20884 2746
rect 1104 2672 20884 2694
rect 2958 2632 2964 2644
rect 2919 2604 2964 2632
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 3326 2632 3332 2644
rect 3287 2604 3332 2632
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 3970 2632 3976 2644
rect 3931 2604 3976 2632
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 5626 2632 5632 2644
rect 5587 2604 5632 2632
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 7650 2632 7656 2644
rect 7611 2604 7656 2632
rect 7650 2592 7656 2604
rect 7708 2592 7714 2644
rect 8297 2635 8355 2641
rect 8297 2601 8309 2635
rect 8343 2632 8355 2635
rect 10226 2632 10232 2644
rect 8343 2604 10232 2632
rect 8343 2601 8355 2604
rect 8297 2595 8355 2601
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 14829 2635 14887 2641
rect 10888 2604 13860 2632
rect 2225 2567 2283 2573
rect 2225 2533 2237 2567
rect 2271 2533 2283 2567
rect 2225 2527 2283 2533
rect 2240 2496 2268 2527
rect 2314 2524 2320 2576
rect 2372 2564 2378 2576
rect 4065 2567 4123 2573
rect 2372 2536 3556 2564
rect 2372 2524 2378 2536
rect 2240 2468 3188 2496
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2428 2283 2431
rect 2314 2428 2320 2440
rect 2271 2400 2320 2428
rect 2271 2397 2283 2400
rect 2225 2391 2283 2397
rect 2314 2388 2320 2400
rect 2372 2388 2378 2440
rect 3160 2437 3188 2468
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2397 3203 2431
rect 3145 2391 3203 2397
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2397 3479 2431
rect 3421 2391 3479 2397
rect 2516 2360 2544 2391
rect 3326 2360 3332 2372
rect 2516 2332 3332 2360
rect 3326 2320 3332 2332
rect 3384 2320 3390 2372
rect 1946 2252 1952 2304
rect 2004 2292 2010 2304
rect 2409 2295 2467 2301
rect 2409 2292 2421 2295
rect 2004 2264 2421 2292
rect 2004 2252 2010 2264
rect 2409 2261 2421 2264
rect 2455 2292 2467 2295
rect 3436 2292 3464 2391
rect 3528 2360 3556 2536
rect 4065 2533 4077 2567
rect 4111 2564 4123 2567
rect 5813 2567 5871 2573
rect 5813 2564 5825 2567
rect 4111 2536 5825 2564
rect 4111 2533 4123 2536
rect 4065 2527 4123 2533
rect 5813 2533 5825 2536
rect 5859 2564 5871 2567
rect 5902 2564 5908 2576
rect 5859 2536 5908 2564
rect 5859 2533 5871 2536
rect 5813 2527 5871 2533
rect 5902 2524 5908 2536
rect 5960 2524 5966 2576
rect 4798 2496 4804 2508
rect 3988 2468 4804 2496
rect 3988 2437 4016 2468
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 7282 2456 7288 2508
rect 7340 2496 7346 2508
rect 9582 2496 9588 2508
rect 7340 2468 8616 2496
rect 9543 2468 9588 2496
rect 7340 2456 7346 2468
rect 7668 2437 7696 2468
rect 8588 2437 8616 2468
rect 9582 2456 9588 2468
rect 9640 2456 9646 2508
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2428 4307 2431
rect 7653 2431 7711 2437
rect 4295 2400 6914 2428
rect 4295 2397 4307 2400
rect 4249 2391 4307 2397
rect 4264 2360 4292 2391
rect 3528 2332 4292 2360
rect 4982 2320 4988 2372
rect 5040 2360 5046 2372
rect 5718 2369 5724 2372
rect 5445 2363 5503 2369
rect 5445 2360 5457 2363
rect 5040 2332 5457 2360
rect 5040 2320 5046 2332
rect 5445 2329 5457 2332
rect 5491 2329 5503 2363
rect 5445 2323 5503 2329
rect 5661 2363 5724 2369
rect 5661 2329 5673 2363
rect 5707 2329 5724 2363
rect 5661 2323 5724 2329
rect 5718 2320 5724 2323
rect 5776 2320 5782 2372
rect 6886 2360 6914 2400
rect 7653 2397 7665 2431
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2428 7895 2431
rect 8297 2431 8355 2437
rect 8297 2428 8309 2431
rect 7883 2400 8309 2428
rect 7883 2397 7895 2400
rect 7837 2391 7895 2397
rect 8297 2397 8309 2400
rect 8343 2397 8355 2431
rect 8297 2391 8355 2397
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 8846 2428 8852 2440
rect 8619 2400 8852 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 7852 2360 7880 2391
rect 8846 2388 8852 2400
rect 8904 2388 8910 2440
rect 9852 2431 9910 2437
rect 9852 2397 9864 2431
rect 9898 2428 9910 2431
rect 10888 2428 10916 2604
rect 10965 2567 11023 2573
rect 10965 2533 10977 2567
rect 11011 2533 11023 2567
rect 10965 2527 11023 2533
rect 10980 2496 11008 2527
rect 11698 2524 11704 2576
rect 11756 2564 11762 2576
rect 11885 2567 11943 2573
rect 11885 2564 11897 2567
rect 11756 2536 11897 2564
rect 11756 2524 11762 2536
rect 11885 2533 11897 2536
rect 11931 2533 11943 2567
rect 11885 2527 11943 2533
rect 11977 2567 12035 2573
rect 11977 2533 11989 2567
rect 12023 2564 12035 2567
rect 13630 2564 13636 2576
rect 12023 2536 13636 2564
rect 12023 2533 12035 2536
rect 11977 2527 12035 2533
rect 13630 2524 13636 2536
rect 13688 2524 13694 2576
rect 13832 2496 13860 2604
rect 14829 2601 14841 2635
rect 14875 2632 14887 2635
rect 14918 2632 14924 2644
rect 14875 2604 14924 2632
rect 14875 2601 14887 2604
rect 14829 2595 14887 2601
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 17770 2496 17776 2508
rect 10980 2468 13768 2496
rect 13832 2468 17776 2496
rect 11882 2428 11888 2440
rect 9898 2400 10916 2428
rect 11843 2400 11888 2428
rect 9898 2397 9910 2400
rect 9852 2391 9910 2397
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 6886 2332 7880 2360
rect 8481 2363 8539 2369
rect 8481 2329 8493 2363
rect 8527 2360 8539 2363
rect 8754 2360 8760 2372
rect 8527 2332 8760 2360
rect 8527 2329 8539 2332
rect 8481 2323 8539 2329
rect 8754 2320 8760 2332
rect 8812 2320 8818 2372
rect 12161 2363 12219 2369
rect 12161 2329 12173 2363
rect 12207 2329 12219 2363
rect 13740 2360 13768 2468
rect 17770 2456 17776 2468
rect 17828 2456 17834 2508
rect 14274 2388 14280 2440
rect 14332 2428 14338 2440
rect 15013 2431 15071 2437
rect 15013 2428 15025 2431
rect 14332 2400 15025 2428
rect 14332 2388 14338 2400
rect 15013 2397 15025 2400
rect 15059 2397 15071 2431
rect 15286 2428 15292 2440
rect 15247 2400 15292 2428
rect 15013 2391 15071 2397
rect 15286 2388 15292 2400
rect 15344 2388 15350 2440
rect 16850 2360 16856 2372
rect 13740 2332 16856 2360
rect 12161 2323 12219 2329
rect 5000 2292 5028 2320
rect 2455 2264 5028 2292
rect 12176 2292 12204 2323
rect 16850 2320 16856 2332
rect 16908 2320 16914 2372
rect 14274 2292 14280 2304
rect 12176 2264 14280 2292
rect 2455 2261 2467 2264
rect 2409 2255 2467 2261
rect 14274 2252 14280 2264
rect 14332 2252 14338 2304
rect 15197 2295 15255 2301
rect 15197 2261 15209 2295
rect 15243 2292 15255 2295
rect 15378 2292 15384 2304
rect 15243 2264 15384 2292
rect 15243 2261 15255 2264
rect 15197 2255 15255 2261
rect 15378 2252 15384 2264
rect 15436 2252 15442 2304
rect 1104 2202 21043 2224
rect 1104 2150 5894 2202
rect 5946 2150 5958 2202
rect 6010 2150 6022 2202
rect 6074 2150 6086 2202
rect 6138 2150 6150 2202
rect 6202 2150 10839 2202
rect 10891 2150 10903 2202
rect 10955 2150 10967 2202
rect 11019 2150 11031 2202
rect 11083 2150 11095 2202
rect 11147 2150 15784 2202
rect 15836 2150 15848 2202
rect 15900 2150 15912 2202
rect 15964 2150 15976 2202
rect 16028 2150 16040 2202
rect 16092 2150 20729 2202
rect 20781 2150 20793 2202
rect 20845 2150 20857 2202
rect 20909 2150 20921 2202
rect 20973 2150 20985 2202
rect 21037 2150 21043 2202
rect 1104 2128 21043 2150
<< via1 >>
rect 5894 19558 5946 19610
rect 5958 19558 6010 19610
rect 6022 19558 6074 19610
rect 6086 19558 6138 19610
rect 6150 19558 6202 19610
rect 10839 19558 10891 19610
rect 10903 19558 10955 19610
rect 10967 19558 11019 19610
rect 11031 19558 11083 19610
rect 11095 19558 11147 19610
rect 15784 19558 15836 19610
rect 15848 19558 15900 19610
rect 15912 19558 15964 19610
rect 15976 19558 16028 19610
rect 16040 19558 16092 19610
rect 20729 19558 20781 19610
rect 20793 19558 20845 19610
rect 20857 19558 20909 19610
rect 20921 19558 20973 19610
rect 20985 19558 21037 19610
rect 3422 19014 3474 19066
rect 3486 19014 3538 19066
rect 3550 19014 3602 19066
rect 3614 19014 3666 19066
rect 3678 19014 3730 19066
rect 8367 19014 8419 19066
rect 8431 19014 8483 19066
rect 8495 19014 8547 19066
rect 8559 19014 8611 19066
rect 8623 19014 8675 19066
rect 13312 19014 13364 19066
rect 13376 19014 13428 19066
rect 13440 19014 13492 19066
rect 13504 19014 13556 19066
rect 13568 19014 13620 19066
rect 18257 19014 18309 19066
rect 18321 19014 18373 19066
rect 18385 19014 18437 19066
rect 18449 19014 18501 19066
rect 18513 19014 18565 19066
rect 2320 18708 2372 18760
rect 1860 18683 1912 18692
rect 1860 18649 1869 18683
rect 1869 18649 1903 18683
rect 1903 18649 1912 18683
rect 1860 18640 1912 18649
rect 5894 18470 5946 18522
rect 5958 18470 6010 18522
rect 6022 18470 6074 18522
rect 6086 18470 6138 18522
rect 6150 18470 6202 18522
rect 10839 18470 10891 18522
rect 10903 18470 10955 18522
rect 10967 18470 11019 18522
rect 11031 18470 11083 18522
rect 11095 18470 11147 18522
rect 15784 18470 15836 18522
rect 15848 18470 15900 18522
rect 15912 18470 15964 18522
rect 15976 18470 16028 18522
rect 16040 18470 16092 18522
rect 20729 18470 20781 18522
rect 20793 18470 20845 18522
rect 20857 18470 20909 18522
rect 20921 18470 20973 18522
rect 20985 18470 21037 18522
rect 3422 17926 3474 17978
rect 3486 17926 3538 17978
rect 3550 17926 3602 17978
rect 3614 17926 3666 17978
rect 3678 17926 3730 17978
rect 8367 17926 8419 17978
rect 8431 17926 8483 17978
rect 8495 17926 8547 17978
rect 8559 17926 8611 17978
rect 8623 17926 8675 17978
rect 13312 17926 13364 17978
rect 13376 17926 13428 17978
rect 13440 17926 13492 17978
rect 13504 17926 13556 17978
rect 13568 17926 13620 17978
rect 18257 17926 18309 17978
rect 18321 17926 18373 17978
rect 18385 17926 18437 17978
rect 18449 17926 18501 17978
rect 18513 17926 18565 17978
rect 5894 17382 5946 17434
rect 5958 17382 6010 17434
rect 6022 17382 6074 17434
rect 6086 17382 6138 17434
rect 6150 17382 6202 17434
rect 10839 17382 10891 17434
rect 10903 17382 10955 17434
rect 10967 17382 11019 17434
rect 11031 17382 11083 17434
rect 11095 17382 11147 17434
rect 15784 17382 15836 17434
rect 15848 17382 15900 17434
rect 15912 17382 15964 17434
rect 15976 17382 16028 17434
rect 16040 17382 16092 17434
rect 20729 17382 20781 17434
rect 20793 17382 20845 17434
rect 20857 17382 20909 17434
rect 20921 17382 20973 17434
rect 20985 17382 21037 17434
rect 5632 17212 5684 17264
rect 5540 17144 5592 17196
rect 7748 17187 7800 17196
rect 5632 17076 5684 17128
rect 7748 17153 7757 17187
rect 7757 17153 7791 17187
rect 7791 17153 7800 17187
rect 7748 17144 7800 17153
rect 7932 17187 7984 17196
rect 7932 17153 7941 17187
rect 7941 17153 7975 17187
rect 7975 17153 7984 17187
rect 7932 17144 7984 17153
rect 6828 17076 6880 17128
rect 4988 17008 5040 17060
rect 4528 16983 4580 16992
rect 4528 16949 4537 16983
rect 4537 16949 4571 16983
rect 4571 16949 4580 16983
rect 4528 16940 4580 16949
rect 6092 16940 6144 16992
rect 6552 16983 6604 16992
rect 6552 16949 6561 16983
rect 6561 16949 6595 16983
rect 6595 16949 6604 16983
rect 6552 16940 6604 16949
rect 7564 16940 7616 16992
rect 3422 16838 3474 16890
rect 3486 16838 3538 16890
rect 3550 16838 3602 16890
rect 3614 16838 3666 16890
rect 3678 16838 3730 16890
rect 8367 16838 8419 16890
rect 8431 16838 8483 16890
rect 8495 16838 8547 16890
rect 8559 16838 8611 16890
rect 8623 16838 8675 16890
rect 13312 16838 13364 16890
rect 13376 16838 13428 16890
rect 13440 16838 13492 16890
rect 13504 16838 13556 16890
rect 13568 16838 13620 16890
rect 18257 16838 18309 16890
rect 18321 16838 18373 16890
rect 18385 16838 18437 16890
rect 18449 16838 18501 16890
rect 18513 16838 18565 16890
rect 5632 16736 5684 16788
rect 4988 16668 5040 16720
rect 3332 16575 3384 16584
rect 3332 16541 3341 16575
rect 3341 16541 3375 16575
rect 3375 16541 3384 16575
rect 3332 16532 3384 16541
rect 4528 16532 4580 16584
rect 5540 16600 5592 16652
rect 6092 16643 6144 16652
rect 6092 16609 6101 16643
rect 6101 16609 6135 16643
rect 6135 16609 6144 16643
rect 6092 16600 6144 16609
rect 6920 16668 6972 16720
rect 5724 16532 5776 16584
rect 7564 16575 7616 16584
rect 7564 16541 7573 16575
rect 7573 16541 7607 16575
rect 7607 16541 7616 16575
rect 7564 16532 7616 16541
rect 7932 16532 7984 16584
rect 11520 16532 11572 16584
rect 15568 16600 15620 16652
rect 4712 16464 4764 16516
rect 3240 16439 3292 16448
rect 3240 16405 3249 16439
rect 3249 16405 3283 16439
rect 3283 16405 3292 16439
rect 3240 16396 3292 16405
rect 5172 16396 5224 16448
rect 5816 16396 5868 16448
rect 6828 16464 6880 16516
rect 7748 16464 7800 16516
rect 7472 16439 7524 16448
rect 7472 16405 7481 16439
rect 7481 16405 7515 16439
rect 7515 16405 7524 16439
rect 11704 16464 11756 16516
rect 14648 16464 14700 16516
rect 7472 16396 7524 16405
rect 15108 16396 15160 16448
rect 5894 16294 5946 16346
rect 5958 16294 6010 16346
rect 6022 16294 6074 16346
rect 6086 16294 6138 16346
rect 6150 16294 6202 16346
rect 10839 16294 10891 16346
rect 10903 16294 10955 16346
rect 10967 16294 11019 16346
rect 11031 16294 11083 16346
rect 11095 16294 11147 16346
rect 15784 16294 15836 16346
rect 15848 16294 15900 16346
rect 15912 16294 15964 16346
rect 15976 16294 16028 16346
rect 16040 16294 16092 16346
rect 20729 16294 20781 16346
rect 20793 16294 20845 16346
rect 20857 16294 20909 16346
rect 20921 16294 20973 16346
rect 20985 16294 21037 16346
rect 3332 16192 3384 16244
rect 4712 16099 4764 16108
rect 4712 16065 4721 16099
rect 4721 16065 4755 16099
rect 4755 16065 4764 16099
rect 4712 16056 4764 16065
rect 4988 16099 5040 16108
rect 4988 16065 4997 16099
rect 4997 16065 5031 16099
rect 5031 16065 5040 16099
rect 5724 16192 5776 16244
rect 11704 16192 11756 16244
rect 4988 16056 5040 16065
rect 5632 16099 5684 16108
rect 5632 16065 5641 16099
rect 5641 16065 5675 16099
rect 5675 16065 5684 16099
rect 5632 16056 5684 16065
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 5172 15988 5224 16040
rect 6920 15988 6972 16040
rect 7288 15988 7340 16040
rect 7564 16056 7616 16108
rect 9404 16099 9456 16108
rect 9404 16065 9413 16099
rect 9413 16065 9447 16099
rect 9447 16065 9456 16099
rect 9404 16056 9456 16065
rect 11244 16056 11296 16108
rect 13084 16099 13136 16108
rect 13084 16065 13093 16099
rect 13093 16065 13127 16099
rect 13127 16065 13136 16099
rect 13084 16056 13136 16065
rect 15200 16124 15252 16176
rect 14372 16056 14424 16108
rect 14556 16099 14608 16108
rect 14556 16065 14565 16099
rect 14565 16065 14599 16099
rect 14599 16065 14608 16099
rect 14556 16056 14608 16065
rect 14648 16099 14700 16108
rect 14648 16065 14658 16099
rect 14658 16065 14692 16099
rect 14692 16065 14700 16099
rect 14648 16056 14700 16065
rect 7840 16031 7892 16040
rect 7840 15997 7849 16031
rect 7849 15997 7883 16031
rect 7883 15997 7892 16031
rect 7840 15988 7892 15997
rect 9680 15988 9732 16040
rect 5080 15920 5132 15972
rect 7472 15920 7524 15972
rect 9220 15920 9272 15972
rect 11796 15988 11848 16040
rect 11336 15920 11388 15972
rect 14740 15988 14792 16040
rect 14924 16099 14976 16108
rect 14924 16065 14933 16099
rect 14933 16065 14967 16099
rect 14967 16065 14976 16099
rect 14924 16056 14976 16065
rect 15108 16056 15160 16108
rect 15660 16056 15712 16108
rect 3792 15895 3844 15904
rect 3792 15861 3801 15895
rect 3801 15861 3835 15895
rect 3835 15861 3844 15895
rect 3792 15852 3844 15861
rect 4712 15852 4764 15904
rect 6920 15852 6972 15904
rect 7656 15895 7708 15904
rect 7656 15861 7665 15895
rect 7665 15861 7699 15895
rect 7699 15861 7708 15895
rect 7656 15852 7708 15861
rect 8852 15852 8904 15904
rect 10416 15852 10468 15904
rect 10876 15852 10928 15904
rect 13176 15920 13228 15972
rect 14188 15920 14240 15972
rect 14556 15920 14608 15972
rect 15936 16031 15988 16040
rect 15936 15997 15945 16031
rect 15945 15997 15979 16031
rect 15979 15997 15988 16031
rect 15936 15988 15988 15997
rect 17040 15988 17092 16040
rect 14648 15852 14700 15904
rect 16120 15852 16172 15904
rect 3422 15750 3474 15802
rect 3486 15750 3538 15802
rect 3550 15750 3602 15802
rect 3614 15750 3666 15802
rect 3678 15750 3730 15802
rect 8367 15750 8419 15802
rect 8431 15750 8483 15802
rect 8495 15750 8547 15802
rect 8559 15750 8611 15802
rect 8623 15750 8675 15802
rect 13312 15750 13364 15802
rect 13376 15750 13428 15802
rect 13440 15750 13492 15802
rect 13504 15750 13556 15802
rect 13568 15750 13620 15802
rect 18257 15750 18309 15802
rect 18321 15750 18373 15802
rect 18385 15750 18437 15802
rect 18449 15750 18501 15802
rect 18513 15750 18565 15802
rect 9220 15691 9272 15700
rect 9220 15657 9229 15691
rect 9229 15657 9263 15691
rect 9263 15657 9272 15691
rect 9220 15648 9272 15657
rect 9404 15648 9456 15700
rect 10876 15691 10928 15700
rect 10876 15657 10885 15691
rect 10885 15657 10919 15691
rect 10919 15657 10928 15691
rect 10876 15648 10928 15657
rect 12532 15648 12584 15700
rect 6828 15580 6880 15632
rect 3148 15512 3200 15564
rect 3240 15444 3292 15496
rect 7748 15487 7800 15496
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 7748 15444 7800 15453
rect 9864 15580 9916 15632
rect 13084 15580 13136 15632
rect 13360 15623 13412 15632
rect 13360 15589 13369 15623
rect 13369 15589 13403 15623
rect 13403 15589 13412 15623
rect 13360 15580 13412 15589
rect 14740 15648 14792 15700
rect 15936 15648 15988 15700
rect 17040 15691 17092 15700
rect 17040 15657 17049 15691
rect 17049 15657 17083 15691
rect 17083 15657 17092 15691
rect 17040 15648 17092 15657
rect 14924 15580 14976 15632
rect 15292 15580 15344 15632
rect 8024 15376 8076 15428
rect 10416 15376 10468 15428
rect 10692 15487 10744 15496
rect 10692 15453 10701 15487
rect 10701 15453 10735 15487
rect 10735 15453 10744 15487
rect 10692 15444 10744 15453
rect 11060 15444 11112 15496
rect 11428 15487 11480 15496
rect 11428 15453 11437 15487
rect 11437 15453 11471 15487
rect 11471 15453 11480 15487
rect 11428 15444 11480 15453
rect 11520 15487 11572 15496
rect 11520 15453 11529 15487
rect 11529 15453 11563 15487
rect 11563 15453 11572 15487
rect 13820 15512 13872 15564
rect 11520 15444 11572 15453
rect 12532 15487 12584 15496
rect 12532 15453 12542 15487
rect 12542 15453 12576 15487
rect 12576 15453 12584 15487
rect 12532 15444 12584 15453
rect 13176 15444 13228 15496
rect 13636 15444 13688 15496
rect 14464 15487 14516 15496
rect 14464 15453 14473 15487
rect 14473 15453 14507 15487
rect 14507 15453 14516 15487
rect 14464 15444 14516 15453
rect 14648 15487 14700 15496
rect 14648 15453 14657 15487
rect 14657 15453 14691 15487
rect 14691 15453 14700 15487
rect 14648 15444 14700 15453
rect 16672 15512 16724 15564
rect 16488 15487 16540 15496
rect 16488 15453 16497 15487
rect 16497 15453 16531 15487
rect 16531 15453 16540 15487
rect 16488 15444 16540 15453
rect 16948 15376 17000 15428
rect 1952 15351 2004 15360
rect 1952 15317 1961 15351
rect 1961 15317 1995 15351
rect 1995 15317 2004 15351
rect 1952 15308 2004 15317
rect 2228 15308 2280 15360
rect 9772 15308 9824 15360
rect 11060 15308 11112 15360
rect 11704 15308 11756 15360
rect 15476 15308 15528 15360
rect 17500 15487 17552 15496
rect 17500 15453 17509 15487
rect 17509 15453 17543 15487
rect 17543 15453 17552 15487
rect 17500 15444 17552 15453
rect 18420 15376 18472 15428
rect 5894 15206 5946 15258
rect 5958 15206 6010 15258
rect 6022 15206 6074 15258
rect 6086 15206 6138 15258
rect 6150 15206 6202 15258
rect 10839 15206 10891 15258
rect 10903 15206 10955 15258
rect 10967 15206 11019 15258
rect 11031 15206 11083 15258
rect 11095 15206 11147 15258
rect 15784 15206 15836 15258
rect 15848 15206 15900 15258
rect 15912 15206 15964 15258
rect 15976 15206 16028 15258
rect 16040 15206 16092 15258
rect 20729 15206 20781 15258
rect 20793 15206 20845 15258
rect 20857 15206 20909 15258
rect 20921 15206 20973 15258
rect 20985 15206 21037 15258
rect 7840 15104 7892 15156
rect 9680 15104 9732 15156
rect 5724 15036 5776 15088
rect 7288 15079 7340 15088
rect 7288 15045 7297 15079
rect 7297 15045 7331 15079
rect 7331 15045 7340 15079
rect 7288 15036 7340 15045
rect 11428 15036 11480 15088
rect 2044 14968 2096 15020
rect 7932 15011 7984 15020
rect 2228 14900 2280 14952
rect 7932 14977 7941 15011
rect 7941 14977 7975 15011
rect 7975 14977 7984 15011
rect 7932 14968 7984 14977
rect 8024 14900 8076 14952
rect 3884 14832 3936 14884
rect 7104 14832 7156 14884
rect 7288 14832 7340 14884
rect 11980 15011 12032 15020
rect 11980 14977 11989 15011
rect 11989 14977 12023 15011
rect 12023 14977 12032 15011
rect 12164 15011 12216 15020
rect 11980 14968 12032 14977
rect 12164 14977 12173 15011
rect 12173 14977 12207 15011
rect 12207 14977 12216 15011
rect 12164 14968 12216 14977
rect 14280 15104 14332 15156
rect 14464 15104 14516 15156
rect 16212 15147 16264 15156
rect 16212 15113 16221 15147
rect 16221 15113 16255 15147
rect 16255 15113 16264 15147
rect 16212 15104 16264 15113
rect 16488 15104 16540 15156
rect 17500 15147 17552 15156
rect 17500 15113 17509 15147
rect 17509 15113 17543 15147
rect 17543 15113 17552 15147
rect 17500 15104 17552 15113
rect 19984 15104 20036 15156
rect 13728 14968 13780 15020
rect 13360 14943 13412 14952
rect 13360 14909 13369 14943
rect 13369 14909 13403 14943
rect 13403 14909 13412 14943
rect 13360 14900 13412 14909
rect 14556 15011 14608 15020
rect 14556 14977 14565 15011
rect 14565 14977 14599 15011
rect 14599 14977 14608 15011
rect 14556 14968 14608 14977
rect 15016 14968 15068 15020
rect 16672 15036 16724 15088
rect 17868 15036 17920 15088
rect 16396 14968 16448 15020
rect 18696 15011 18748 15020
rect 3148 14764 3200 14816
rect 6828 14764 6880 14816
rect 17132 14832 17184 14884
rect 18696 14977 18705 15011
rect 18705 14977 18739 15011
rect 18739 14977 18748 15011
rect 18696 14968 18748 14977
rect 18972 15011 19024 15020
rect 18972 14977 18981 15011
rect 18981 14977 19015 15011
rect 19015 14977 19024 15011
rect 18972 14968 19024 14977
rect 18420 14832 18472 14884
rect 8208 14764 8260 14816
rect 10600 14764 10652 14816
rect 11796 14764 11848 14816
rect 13084 14764 13136 14816
rect 14096 14764 14148 14816
rect 17868 14807 17920 14816
rect 17868 14773 17877 14807
rect 17877 14773 17911 14807
rect 17911 14773 17920 14807
rect 17868 14764 17920 14773
rect 17960 14807 18012 14816
rect 17960 14773 17969 14807
rect 17969 14773 18003 14807
rect 18003 14773 18012 14807
rect 17960 14764 18012 14773
rect 3422 14662 3474 14714
rect 3486 14662 3538 14714
rect 3550 14662 3602 14714
rect 3614 14662 3666 14714
rect 3678 14662 3730 14714
rect 8367 14662 8419 14714
rect 8431 14662 8483 14714
rect 8495 14662 8547 14714
rect 8559 14662 8611 14714
rect 8623 14662 8675 14714
rect 13312 14662 13364 14714
rect 13376 14662 13428 14714
rect 13440 14662 13492 14714
rect 13504 14662 13556 14714
rect 13568 14662 13620 14714
rect 18257 14662 18309 14714
rect 18321 14662 18373 14714
rect 18385 14662 18437 14714
rect 18449 14662 18501 14714
rect 18513 14662 18565 14714
rect 3056 14560 3108 14612
rect 3792 14560 3844 14612
rect 8208 14603 8260 14612
rect 8208 14569 8217 14603
rect 8217 14569 8251 14603
rect 8251 14569 8260 14603
rect 8208 14560 8260 14569
rect 10692 14560 10744 14612
rect 4160 14492 4212 14544
rect 4988 14492 5040 14544
rect 9496 14492 9548 14544
rect 3056 14399 3108 14408
rect 3056 14365 3065 14399
rect 3065 14365 3099 14399
rect 3099 14365 3108 14399
rect 3332 14399 3384 14408
rect 3056 14356 3108 14365
rect 3332 14365 3341 14399
rect 3341 14365 3375 14399
rect 3375 14365 3384 14399
rect 3332 14356 3384 14365
rect 3424 14399 3476 14408
rect 3424 14365 3433 14399
rect 3433 14365 3467 14399
rect 3467 14365 3476 14399
rect 3424 14356 3476 14365
rect 3884 14356 3936 14408
rect 4160 14399 4212 14408
rect 4160 14365 4169 14399
rect 4169 14365 4203 14399
rect 4203 14365 4212 14399
rect 4160 14356 4212 14365
rect 2044 14288 2096 14340
rect 2228 14288 2280 14340
rect 3240 14288 3292 14340
rect 2412 14220 2464 14272
rect 2780 14263 2832 14272
rect 2780 14229 2789 14263
rect 2789 14229 2823 14263
rect 2823 14229 2832 14263
rect 5080 14356 5132 14408
rect 5264 14424 5316 14476
rect 7564 14424 7616 14476
rect 7932 14424 7984 14476
rect 11244 14492 11296 14544
rect 11520 14492 11572 14544
rect 11612 14492 11664 14544
rect 5172 14331 5224 14340
rect 5172 14297 5181 14331
rect 5181 14297 5215 14331
rect 5215 14297 5224 14331
rect 5172 14288 5224 14297
rect 5724 14356 5776 14408
rect 5816 14356 5868 14408
rect 8024 14356 8076 14408
rect 9220 14399 9272 14408
rect 9220 14365 9262 14399
rect 9262 14365 9272 14399
rect 9680 14399 9732 14408
rect 9220 14356 9272 14365
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 9956 14356 10008 14408
rect 11796 14424 11848 14476
rect 12164 14560 12216 14612
rect 14280 14560 14332 14612
rect 14832 14560 14884 14612
rect 15476 14560 15528 14612
rect 7288 14288 7340 14340
rect 10784 14356 10836 14408
rect 11704 14399 11756 14408
rect 11704 14365 11713 14399
rect 11713 14365 11747 14399
rect 11747 14365 11756 14399
rect 11704 14356 11756 14365
rect 15568 14424 15620 14476
rect 19616 14560 19668 14612
rect 16304 14492 16356 14544
rect 11336 14288 11388 14340
rect 13176 14356 13228 14408
rect 13360 14399 13412 14408
rect 13360 14365 13369 14399
rect 13369 14365 13403 14399
rect 13403 14365 13412 14399
rect 13360 14356 13412 14365
rect 13636 14399 13688 14408
rect 13636 14365 13645 14399
rect 13645 14365 13679 14399
rect 13679 14365 13688 14399
rect 13636 14356 13688 14365
rect 14096 14356 14148 14408
rect 14556 14356 14608 14408
rect 16212 14356 16264 14408
rect 16488 14399 16540 14408
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 16672 14399 16724 14408
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 16672 14356 16724 14365
rect 18236 14399 18288 14408
rect 18236 14365 18245 14399
rect 18245 14365 18279 14399
rect 18279 14365 18288 14399
rect 18236 14356 18288 14365
rect 18420 14356 18472 14408
rect 14464 14288 14516 14340
rect 2780 14220 2832 14229
rect 5080 14220 5132 14272
rect 5540 14263 5592 14272
rect 5540 14229 5549 14263
rect 5549 14229 5583 14263
rect 5583 14229 5592 14263
rect 5540 14220 5592 14229
rect 7472 14220 7524 14272
rect 9312 14263 9364 14272
rect 9312 14229 9321 14263
rect 9321 14229 9355 14263
rect 9355 14229 9364 14263
rect 9312 14220 9364 14229
rect 13084 14220 13136 14272
rect 13728 14220 13780 14272
rect 14004 14220 14056 14272
rect 18880 14288 18932 14340
rect 14648 14220 14700 14272
rect 15292 14220 15344 14272
rect 15384 14220 15436 14272
rect 18052 14220 18104 14272
rect 5894 14118 5946 14170
rect 5958 14118 6010 14170
rect 6022 14118 6074 14170
rect 6086 14118 6138 14170
rect 6150 14118 6202 14170
rect 10839 14118 10891 14170
rect 10903 14118 10955 14170
rect 10967 14118 11019 14170
rect 11031 14118 11083 14170
rect 11095 14118 11147 14170
rect 15784 14118 15836 14170
rect 15848 14118 15900 14170
rect 15912 14118 15964 14170
rect 15976 14118 16028 14170
rect 16040 14118 16092 14170
rect 20729 14118 20781 14170
rect 20793 14118 20845 14170
rect 20857 14118 20909 14170
rect 20921 14118 20973 14170
rect 20985 14118 21037 14170
rect 1952 14016 2004 14068
rect 3332 14016 3384 14068
rect 5172 14016 5224 14068
rect 2412 13948 2464 14000
rect 7012 14016 7064 14068
rect 7104 14016 7156 14068
rect 6828 13948 6880 14000
rect 2044 13880 2096 13932
rect 2964 13812 3016 13864
rect 3148 13923 3200 13932
rect 3148 13889 3157 13923
rect 3157 13889 3191 13923
rect 3191 13889 3200 13923
rect 3148 13880 3200 13889
rect 3240 13812 3292 13864
rect 5632 13880 5684 13932
rect 6920 13957 6930 13966
rect 6930 13957 6964 13966
rect 6964 13957 6972 13966
rect 6920 13914 6972 13957
rect 7288 13948 7340 14000
rect 5724 13812 5776 13864
rect 6644 13855 6696 13864
rect 6644 13821 6653 13855
rect 6653 13821 6687 13855
rect 6687 13821 6696 13855
rect 6644 13812 6696 13821
rect 7196 13880 7248 13932
rect 7840 13923 7892 13932
rect 7840 13889 7849 13923
rect 7849 13889 7883 13923
rect 7883 13889 7892 13923
rect 7840 13880 7892 13889
rect 8024 13923 8076 13932
rect 8024 13889 8033 13923
rect 8033 13889 8067 13923
rect 8067 13889 8076 13923
rect 8024 13880 8076 13889
rect 9036 13880 9088 13932
rect 2872 13744 2924 13796
rect 10692 14016 10744 14068
rect 12072 14016 12124 14068
rect 13360 14016 13412 14068
rect 15476 14016 15528 14068
rect 16488 14016 16540 14068
rect 9220 13880 9272 13932
rect 11888 13880 11940 13932
rect 12900 13923 12952 13932
rect 7932 13744 7984 13796
rect 8944 13744 8996 13796
rect 11796 13812 11848 13864
rect 12348 13812 12400 13864
rect 12900 13889 12909 13923
rect 12909 13889 12943 13923
rect 12943 13889 12952 13923
rect 12900 13880 12952 13889
rect 14556 13880 14608 13932
rect 14740 13923 14792 13932
rect 14740 13889 14749 13923
rect 14749 13889 14783 13923
rect 14783 13889 14792 13923
rect 14740 13880 14792 13889
rect 15292 13948 15344 14000
rect 15660 13948 15712 14000
rect 16396 13948 16448 14000
rect 17960 14016 18012 14068
rect 18788 14016 18840 14068
rect 19616 14059 19668 14068
rect 17500 13880 17552 13932
rect 14004 13812 14056 13864
rect 17960 13880 18012 13932
rect 18236 13880 18288 13932
rect 18420 13923 18472 13932
rect 18420 13889 18429 13923
rect 18429 13889 18463 13923
rect 18463 13889 18472 13923
rect 18972 13948 19024 14000
rect 19616 14025 19625 14059
rect 19625 14025 19659 14059
rect 19659 14025 19668 14059
rect 19616 14016 19668 14025
rect 18420 13880 18472 13889
rect 18788 13880 18840 13932
rect 14464 13787 14516 13796
rect 1584 13719 1636 13728
rect 1584 13685 1593 13719
rect 1593 13685 1627 13719
rect 1627 13685 1636 13719
rect 1584 13676 1636 13685
rect 10416 13676 10468 13728
rect 13176 13676 13228 13728
rect 14464 13753 14473 13787
rect 14473 13753 14507 13787
rect 14507 13753 14516 13787
rect 14464 13744 14516 13753
rect 15200 13744 15252 13796
rect 16304 13744 16356 13796
rect 17132 13787 17184 13796
rect 17132 13753 17141 13787
rect 17141 13753 17175 13787
rect 17175 13753 17184 13787
rect 19800 13880 19852 13932
rect 20076 13855 20128 13864
rect 20076 13821 20085 13855
rect 20085 13821 20119 13855
rect 20119 13821 20128 13855
rect 20076 13812 20128 13821
rect 19984 13787 20036 13796
rect 17132 13744 17184 13753
rect 19984 13753 19993 13787
rect 19993 13753 20027 13787
rect 20027 13753 20036 13787
rect 19984 13744 20036 13753
rect 14188 13676 14240 13728
rect 14556 13719 14608 13728
rect 14556 13685 14565 13719
rect 14565 13685 14599 13719
rect 14599 13685 14608 13719
rect 14556 13676 14608 13685
rect 14648 13676 14700 13728
rect 15016 13676 15068 13728
rect 18144 13719 18196 13728
rect 18144 13685 18153 13719
rect 18153 13685 18187 13719
rect 18187 13685 18196 13719
rect 18144 13676 18196 13685
rect 3422 13574 3474 13626
rect 3486 13574 3538 13626
rect 3550 13574 3602 13626
rect 3614 13574 3666 13626
rect 3678 13574 3730 13626
rect 8367 13574 8419 13626
rect 8431 13574 8483 13626
rect 8495 13574 8547 13626
rect 8559 13574 8611 13626
rect 8623 13574 8675 13626
rect 13312 13574 13364 13626
rect 13376 13574 13428 13626
rect 13440 13574 13492 13626
rect 13504 13574 13556 13626
rect 13568 13574 13620 13626
rect 18257 13574 18309 13626
rect 18321 13574 18373 13626
rect 18385 13574 18437 13626
rect 18449 13574 18501 13626
rect 18513 13574 18565 13626
rect 7564 13515 7616 13524
rect 7564 13481 7573 13515
rect 7573 13481 7607 13515
rect 7607 13481 7616 13515
rect 7564 13472 7616 13481
rect 9312 13472 9364 13524
rect 12900 13472 12952 13524
rect 14464 13472 14516 13524
rect 17500 13515 17552 13524
rect 17500 13481 17509 13515
rect 17509 13481 17543 13515
rect 17543 13481 17552 13515
rect 17500 13472 17552 13481
rect 2964 13404 3016 13456
rect 3240 13404 3292 13456
rect 11612 13447 11664 13456
rect 11612 13413 11621 13447
rect 11621 13413 11655 13447
rect 11655 13413 11664 13447
rect 11612 13404 11664 13413
rect 4712 13379 4764 13388
rect 4712 13345 4721 13379
rect 4721 13345 4755 13379
rect 4755 13345 4764 13379
rect 4712 13336 4764 13345
rect 4896 13379 4948 13388
rect 4896 13345 4905 13379
rect 4905 13345 4939 13379
rect 4939 13345 4948 13379
rect 4896 13336 4948 13345
rect 8944 13336 8996 13388
rect 2044 13268 2096 13320
rect 5632 13268 5684 13320
rect 6828 13268 6880 13320
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 12348 13336 12400 13388
rect 2872 13200 2924 13252
rect 4068 13200 4120 13252
rect 8208 13200 8260 13252
rect 11796 13268 11848 13320
rect 12072 13268 12124 13320
rect 14924 13336 14976 13388
rect 15384 13336 15436 13388
rect 18144 13379 18196 13388
rect 18144 13345 18153 13379
rect 18153 13345 18187 13379
rect 18187 13345 18196 13379
rect 18144 13336 18196 13345
rect 10692 13200 10744 13252
rect 16856 13268 16908 13320
rect 17776 13311 17828 13320
rect 17776 13277 17785 13311
rect 17785 13277 17819 13311
rect 17819 13277 17828 13311
rect 18052 13311 18104 13320
rect 17776 13268 17828 13277
rect 18052 13277 18061 13311
rect 18061 13277 18095 13311
rect 18095 13277 18104 13311
rect 18052 13268 18104 13277
rect 19892 13311 19944 13320
rect 19892 13277 19901 13311
rect 19901 13277 19935 13311
rect 19935 13277 19944 13311
rect 19892 13268 19944 13277
rect 20076 13200 20128 13252
rect 4160 13132 4212 13184
rect 4620 13175 4672 13184
rect 4620 13141 4629 13175
rect 4629 13141 4663 13175
rect 4663 13141 4672 13175
rect 4620 13132 4672 13141
rect 5894 13030 5946 13082
rect 5958 13030 6010 13082
rect 6022 13030 6074 13082
rect 6086 13030 6138 13082
rect 6150 13030 6202 13082
rect 10839 13030 10891 13082
rect 10903 13030 10955 13082
rect 10967 13030 11019 13082
rect 11031 13030 11083 13082
rect 11095 13030 11147 13082
rect 15784 13030 15836 13082
rect 15848 13030 15900 13082
rect 15912 13030 15964 13082
rect 15976 13030 16028 13082
rect 16040 13030 16092 13082
rect 20729 13030 20781 13082
rect 20793 13030 20845 13082
rect 20857 13030 20909 13082
rect 20921 13030 20973 13082
rect 20985 13030 21037 13082
rect 4160 12971 4212 12980
rect 4160 12937 4169 12971
rect 4169 12937 4203 12971
rect 4203 12937 4212 12971
rect 4160 12928 4212 12937
rect 5540 12928 5592 12980
rect 7104 12928 7156 12980
rect 13176 12928 13228 12980
rect 15568 12928 15620 12980
rect 16856 12971 16908 12980
rect 16856 12937 16865 12971
rect 16865 12937 16899 12971
rect 16899 12937 16908 12971
rect 16856 12928 16908 12937
rect 4252 12860 4304 12912
rect 4344 12860 4396 12912
rect 9220 12860 9272 12912
rect 10692 12860 10744 12912
rect 3332 12792 3384 12844
rect 5356 12792 5408 12844
rect 5724 12792 5776 12844
rect 6920 12792 6972 12844
rect 7196 12835 7248 12844
rect 7196 12801 7205 12835
rect 7205 12801 7239 12835
rect 7239 12801 7248 12835
rect 7196 12792 7248 12801
rect 7380 12792 7432 12844
rect 9036 12835 9088 12844
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9036 12792 9088 12801
rect 9404 12792 9456 12844
rect 13176 12792 13228 12844
rect 14924 12792 14976 12844
rect 16028 12835 16080 12844
rect 16028 12801 16037 12835
rect 16037 12801 16071 12835
rect 16071 12801 16080 12835
rect 16028 12792 16080 12801
rect 16672 12792 16724 12844
rect 17224 12835 17276 12844
rect 17224 12801 17233 12835
rect 17233 12801 17267 12835
rect 17267 12801 17276 12835
rect 17224 12792 17276 12801
rect 17960 12792 18012 12844
rect 18604 12792 18656 12844
rect 19524 12792 19576 12844
rect 19892 12835 19944 12844
rect 19892 12801 19901 12835
rect 19901 12801 19935 12835
rect 19935 12801 19944 12835
rect 19892 12792 19944 12801
rect 2044 12724 2096 12776
rect 3056 12588 3108 12640
rect 4896 12724 4948 12776
rect 7288 12724 7340 12776
rect 8944 12767 8996 12776
rect 8944 12733 8953 12767
rect 8953 12733 8987 12767
rect 8987 12733 8996 12767
rect 8944 12724 8996 12733
rect 4068 12656 4120 12708
rect 4344 12588 4396 12640
rect 4896 12631 4948 12640
rect 4896 12597 4905 12631
rect 4905 12597 4939 12631
rect 4939 12597 4948 12631
rect 4896 12588 4948 12597
rect 7012 12631 7064 12640
rect 7012 12597 7021 12631
rect 7021 12597 7055 12631
rect 7055 12597 7064 12631
rect 7012 12588 7064 12597
rect 8760 12631 8812 12640
rect 8760 12597 8769 12631
rect 8769 12597 8803 12631
rect 8803 12597 8812 12631
rect 8760 12588 8812 12597
rect 9220 12767 9272 12776
rect 9220 12733 9229 12767
rect 9229 12733 9263 12767
rect 9263 12733 9272 12767
rect 9220 12724 9272 12733
rect 10508 12724 10560 12776
rect 12992 12724 13044 12776
rect 16580 12724 16632 12776
rect 12072 12656 12124 12708
rect 14556 12656 14608 12708
rect 17868 12724 17920 12776
rect 18696 12656 18748 12708
rect 9220 12588 9272 12640
rect 11704 12631 11756 12640
rect 11704 12597 11713 12631
rect 11713 12597 11747 12631
rect 11747 12597 11756 12631
rect 11704 12588 11756 12597
rect 14740 12588 14792 12640
rect 15292 12588 15344 12640
rect 19708 12631 19760 12640
rect 19708 12597 19717 12631
rect 19717 12597 19751 12631
rect 19751 12597 19760 12631
rect 19708 12588 19760 12597
rect 3422 12486 3474 12538
rect 3486 12486 3538 12538
rect 3550 12486 3602 12538
rect 3614 12486 3666 12538
rect 3678 12486 3730 12538
rect 8367 12486 8419 12538
rect 8431 12486 8483 12538
rect 8495 12486 8547 12538
rect 8559 12486 8611 12538
rect 8623 12486 8675 12538
rect 13312 12486 13364 12538
rect 13376 12486 13428 12538
rect 13440 12486 13492 12538
rect 13504 12486 13556 12538
rect 13568 12486 13620 12538
rect 18257 12486 18309 12538
rect 18321 12486 18373 12538
rect 18385 12486 18437 12538
rect 18449 12486 18501 12538
rect 18513 12486 18565 12538
rect 4068 12384 4120 12436
rect 5448 12384 5500 12436
rect 9128 12427 9180 12436
rect 9128 12393 9137 12427
rect 9137 12393 9171 12427
rect 9171 12393 9180 12427
rect 9128 12384 9180 12393
rect 9404 12384 9456 12436
rect 10508 12384 10560 12436
rect 10692 12384 10744 12436
rect 11796 12427 11848 12436
rect 11796 12393 11805 12427
rect 11805 12393 11839 12427
rect 11839 12393 11848 12427
rect 11796 12384 11848 12393
rect 6644 12316 6696 12368
rect 13268 12384 13320 12436
rect 15292 12384 15344 12436
rect 17776 12384 17828 12436
rect 19524 12384 19576 12436
rect 19800 12384 19852 12436
rect 20168 12384 20220 12436
rect 2964 12248 3016 12300
rect 2872 12180 2924 12232
rect 4068 12248 4120 12300
rect 4896 12248 4948 12300
rect 5448 12291 5500 12300
rect 5448 12257 5457 12291
rect 5457 12257 5491 12291
rect 5491 12257 5500 12291
rect 5448 12248 5500 12257
rect 5632 12248 5684 12300
rect 7288 12291 7340 12300
rect 4620 12180 4672 12232
rect 7288 12257 7297 12291
rect 7297 12257 7331 12291
rect 7331 12257 7340 12291
rect 7288 12248 7340 12257
rect 7104 12223 7156 12232
rect 7104 12189 7113 12223
rect 7113 12189 7147 12223
rect 7147 12189 7156 12223
rect 7104 12180 7156 12189
rect 7932 12180 7984 12232
rect 9036 12248 9088 12300
rect 8944 12180 8996 12232
rect 9128 12180 9180 12232
rect 9312 12223 9364 12232
rect 9312 12189 9321 12223
rect 9321 12189 9355 12223
rect 9355 12189 9364 12223
rect 9312 12180 9364 12189
rect 9864 12180 9916 12232
rect 10784 12180 10836 12232
rect 15108 12316 15160 12368
rect 17500 12316 17552 12368
rect 14372 12291 14424 12300
rect 11612 12180 11664 12232
rect 11980 12223 12032 12232
rect 11980 12189 11989 12223
rect 11989 12189 12023 12223
rect 12023 12189 12032 12223
rect 11980 12180 12032 12189
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 12072 12180 12124 12189
rect 12256 12223 12308 12232
rect 12256 12189 12265 12223
rect 12265 12189 12299 12223
rect 12299 12189 12308 12223
rect 12256 12180 12308 12189
rect 13268 12223 13320 12232
rect 4436 12112 4488 12164
rect 5264 12112 5316 12164
rect 9680 12155 9732 12164
rect 9680 12121 9689 12155
rect 9689 12121 9723 12155
rect 9723 12121 9732 12155
rect 9680 12112 9732 12121
rect 9772 12155 9824 12164
rect 9772 12121 9781 12155
rect 9781 12121 9815 12155
rect 9815 12121 9824 12155
rect 9772 12112 9824 12121
rect 10508 12112 10560 12164
rect 12440 12112 12492 12164
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 1860 12087 1912 12096
rect 1860 12053 1869 12087
rect 1869 12053 1903 12087
rect 1903 12053 1912 12087
rect 1860 12044 1912 12053
rect 2228 12087 2280 12096
rect 2228 12053 2237 12087
rect 2237 12053 2271 12087
rect 2271 12053 2280 12087
rect 2228 12044 2280 12053
rect 3332 12087 3384 12096
rect 3332 12053 3341 12087
rect 3341 12053 3375 12087
rect 3375 12053 3384 12087
rect 3332 12044 3384 12053
rect 4896 12044 4948 12096
rect 6920 12044 6972 12096
rect 8392 12087 8444 12096
rect 8392 12053 8407 12087
rect 8407 12053 8441 12087
rect 8441 12053 8444 12087
rect 8392 12044 8444 12053
rect 10692 12044 10744 12096
rect 10784 12044 10836 12096
rect 14372 12257 14381 12291
rect 14381 12257 14415 12291
rect 14415 12257 14424 12291
rect 14372 12248 14424 12257
rect 16580 12291 16632 12300
rect 13636 12180 13688 12232
rect 14280 12180 14332 12232
rect 14648 12223 14700 12232
rect 14648 12189 14657 12223
rect 14657 12189 14691 12223
rect 14691 12189 14700 12223
rect 14924 12223 14976 12232
rect 14648 12180 14700 12189
rect 14924 12189 14933 12223
rect 14933 12189 14967 12223
rect 14967 12189 14976 12223
rect 14924 12180 14976 12189
rect 15016 12180 15068 12232
rect 14464 12112 14516 12164
rect 15108 12112 15160 12164
rect 16212 12180 16264 12232
rect 16580 12257 16589 12291
rect 16589 12257 16623 12291
rect 16623 12257 16632 12291
rect 16580 12248 16632 12257
rect 17592 12180 17644 12232
rect 17868 12223 17920 12232
rect 17868 12189 17891 12223
rect 17891 12189 17920 12223
rect 17868 12180 17920 12189
rect 19616 12316 19668 12368
rect 18880 12248 18932 12300
rect 18052 12223 18104 12232
rect 18052 12189 18061 12223
rect 18061 12189 18095 12223
rect 18095 12189 18104 12223
rect 18052 12180 18104 12189
rect 16028 12112 16080 12164
rect 15200 12044 15252 12096
rect 18604 12180 18656 12232
rect 19248 12180 19300 12232
rect 19892 12180 19944 12232
rect 5894 11942 5946 11994
rect 5958 11942 6010 11994
rect 6022 11942 6074 11994
rect 6086 11942 6138 11994
rect 6150 11942 6202 11994
rect 10839 11942 10891 11994
rect 10903 11942 10955 11994
rect 10967 11942 11019 11994
rect 11031 11942 11083 11994
rect 11095 11942 11147 11994
rect 15784 11942 15836 11994
rect 15848 11942 15900 11994
rect 15912 11942 15964 11994
rect 15976 11942 16028 11994
rect 16040 11942 16092 11994
rect 20729 11942 20781 11994
rect 20793 11942 20845 11994
rect 20857 11942 20909 11994
rect 20921 11942 20973 11994
rect 20985 11942 21037 11994
rect 2320 11840 2372 11892
rect 2780 11840 2832 11892
rect 7656 11840 7708 11892
rect 9772 11840 9824 11892
rect 11244 11840 11296 11892
rect 11980 11840 12032 11892
rect 12348 11883 12400 11892
rect 4344 11772 4396 11824
rect 8760 11772 8812 11824
rect 9956 11772 10008 11824
rect 10600 11772 10652 11824
rect 12348 11849 12357 11883
rect 12357 11849 12391 11883
rect 12391 11849 12400 11883
rect 12348 11840 12400 11849
rect 13452 11840 13504 11892
rect 13636 11840 13688 11892
rect 2780 11704 2832 11756
rect 3240 11747 3292 11756
rect 3240 11713 3249 11747
rect 3249 11713 3283 11747
rect 3283 11713 3292 11747
rect 3240 11704 3292 11713
rect 3884 11704 3936 11756
rect 4436 11747 4488 11756
rect 2872 11636 2924 11688
rect 4436 11713 4445 11747
rect 4445 11713 4479 11747
rect 4479 11713 4488 11747
rect 4436 11704 4488 11713
rect 4620 11747 4672 11756
rect 4620 11713 4629 11747
rect 4629 11713 4663 11747
rect 4663 11713 4672 11747
rect 4620 11704 4672 11713
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 5816 11636 5868 11688
rect 5540 11568 5592 11620
rect 6920 11704 6972 11756
rect 8392 11704 8444 11756
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 10692 11747 10744 11756
rect 10692 11713 10701 11747
rect 10701 11713 10735 11747
rect 10735 11713 10744 11747
rect 10692 11704 10744 11713
rect 11612 11704 11664 11756
rect 12072 11747 12124 11756
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 7288 11636 7340 11688
rect 11704 11636 11756 11688
rect 7564 11568 7616 11620
rect 11520 11568 11572 11620
rect 13176 11772 13228 11824
rect 16672 11840 16724 11892
rect 19248 11883 19300 11892
rect 19248 11849 19257 11883
rect 19257 11849 19291 11883
rect 19291 11849 19300 11883
rect 19248 11840 19300 11849
rect 19984 11840 20036 11892
rect 12992 11704 13044 11756
rect 13544 11704 13596 11756
rect 14096 11747 14148 11756
rect 14096 11713 14105 11747
rect 14105 11713 14139 11747
rect 14139 11713 14148 11747
rect 14096 11704 14148 11713
rect 14280 11747 14332 11756
rect 14280 11713 14289 11747
rect 14289 11713 14323 11747
rect 14323 11713 14332 11747
rect 14280 11704 14332 11713
rect 15108 11704 15160 11756
rect 15292 11704 15344 11756
rect 15660 11747 15712 11756
rect 15660 11713 15669 11747
rect 15669 11713 15703 11747
rect 15703 11713 15712 11747
rect 15660 11704 15712 11713
rect 15752 11747 15804 11756
rect 15752 11713 15762 11747
rect 15762 11713 15796 11747
rect 15796 11713 15804 11747
rect 16212 11772 16264 11824
rect 17040 11772 17092 11824
rect 17868 11772 17920 11824
rect 15752 11704 15804 11713
rect 14188 11636 14240 11688
rect 3240 11500 3292 11552
rect 3792 11500 3844 11552
rect 7196 11500 7248 11552
rect 10324 11543 10376 11552
rect 10324 11509 10333 11543
rect 10333 11509 10367 11543
rect 10367 11509 10376 11543
rect 10324 11500 10376 11509
rect 12348 11568 12400 11620
rect 16396 11704 16448 11756
rect 17500 11747 17552 11756
rect 17500 11713 17509 11747
rect 17509 11713 17543 11747
rect 17543 11713 17552 11747
rect 17500 11704 17552 11713
rect 19156 11704 19208 11756
rect 19432 11772 19484 11824
rect 19708 11704 19760 11756
rect 17316 11679 17368 11688
rect 17316 11645 17325 11679
rect 17325 11645 17359 11679
rect 17359 11645 17368 11679
rect 17316 11636 17368 11645
rect 18880 11636 18932 11688
rect 19248 11568 19300 11620
rect 12256 11500 12308 11552
rect 13820 11500 13872 11552
rect 14096 11500 14148 11552
rect 14280 11500 14332 11552
rect 15568 11500 15620 11552
rect 16304 11543 16356 11552
rect 16304 11509 16313 11543
rect 16313 11509 16347 11543
rect 16347 11509 16356 11543
rect 16304 11500 16356 11509
rect 16396 11500 16448 11552
rect 19892 11500 19944 11552
rect 3422 11398 3474 11450
rect 3486 11398 3538 11450
rect 3550 11398 3602 11450
rect 3614 11398 3666 11450
rect 3678 11398 3730 11450
rect 8367 11398 8419 11450
rect 8431 11398 8483 11450
rect 8495 11398 8547 11450
rect 8559 11398 8611 11450
rect 8623 11398 8675 11450
rect 13312 11398 13364 11450
rect 13376 11398 13428 11450
rect 13440 11398 13492 11450
rect 13504 11398 13556 11450
rect 13568 11398 13620 11450
rect 18257 11398 18309 11450
rect 18321 11398 18373 11450
rect 18385 11398 18437 11450
rect 18449 11398 18501 11450
rect 18513 11398 18565 11450
rect 12440 11339 12492 11348
rect 12440 11305 12449 11339
rect 12449 11305 12483 11339
rect 12483 11305 12492 11339
rect 12440 11296 12492 11305
rect 15016 11296 15068 11348
rect 15752 11296 15804 11348
rect 1952 11228 2004 11280
rect 7104 11228 7156 11280
rect 13084 11228 13136 11280
rect 14464 11228 14516 11280
rect 3332 11160 3384 11212
rect 3884 11160 3936 11212
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 7196 11160 7248 11169
rect 7564 11160 7616 11212
rect 14188 11160 14240 11212
rect 18052 11228 18104 11280
rect 18880 11228 18932 11280
rect 17224 11160 17276 11212
rect 19248 11160 19300 11212
rect 2964 11092 3016 11144
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 14464 11092 14516 11144
rect 16396 11092 16448 11144
rect 17592 11135 17644 11144
rect 17592 11101 17601 11135
rect 17601 11101 17635 11135
rect 17635 11101 17644 11135
rect 17592 11092 17644 11101
rect 19156 11092 19208 11144
rect 20168 11203 20220 11212
rect 20168 11169 20177 11203
rect 20177 11169 20211 11203
rect 20211 11169 20220 11203
rect 20168 11160 20220 11169
rect 2872 11024 2924 11076
rect 7196 11024 7248 11076
rect 11336 11024 11388 11076
rect 19984 11024 20036 11076
rect 2780 10956 2832 11008
rect 2964 10956 3016 11008
rect 14004 10956 14056 11008
rect 16856 10956 16908 11008
rect 17776 10956 17828 11008
rect 5894 10854 5946 10906
rect 5958 10854 6010 10906
rect 6022 10854 6074 10906
rect 6086 10854 6138 10906
rect 6150 10854 6202 10906
rect 10839 10854 10891 10906
rect 10903 10854 10955 10906
rect 10967 10854 11019 10906
rect 11031 10854 11083 10906
rect 11095 10854 11147 10906
rect 15784 10854 15836 10906
rect 15848 10854 15900 10906
rect 15912 10854 15964 10906
rect 15976 10854 16028 10906
rect 16040 10854 16092 10906
rect 20729 10854 20781 10906
rect 20793 10854 20845 10906
rect 20857 10854 20909 10906
rect 20921 10854 20973 10906
rect 20985 10854 21037 10906
rect 6828 10752 6880 10804
rect 15476 10752 15528 10804
rect 1676 10727 1728 10736
rect 1676 10693 1685 10727
rect 1685 10693 1719 10727
rect 1719 10693 1728 10727
rect 1676 10684 1728 10693
rect 3976 10684 4028 10736
rect 10324 10684 10376 10736
rect 19156 10752 19208 10804
rect 13820 10659 13872 10668
rect 13820 10625 13829 10659
rect 13829 10625 13863 10659
rect 13863 10625 13872 10659
rect 13820 10616 13872 10625
rect 14924 10616 14976 10668
rect 16856 10659 16908 10668
rect 16856 10625 16865 10659
rect 16865 10625 16899 10659
rect 16899 10625 16908 10659
rect 16856 10616 16908 10625
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 19432 10684 19484 10736
rect 19800 10684 19852 10736
rect 17040 10616 17092 10625
rect 19248 10616 19300 10668
rect 19616 10659 19668 10668
rect 19616 10625 19625 10659
rect 19625 10625 19659 10659
rect 19659 10625 19668 10659
rect 19616 10616 19668 10625
rect 7012 10548 7064 10600
rect 9772 10591 9824 10600
rect 9772 10557 9781 10591
rect 9781 10557 9815 10591
rect 9815 10557 9824 10591
rect 9772 10548 9824 10557
rect 11244 10548 11296 10600
rect 13176 10548 13228 10600
rect 18052 10548 18104 10600
rect 9128 10523 9180 10532
rect 9128 10489 9137 10523
rect 9137 10489 9171 10523
rect 9171 10489 9180 10523
rect 9128 10480 9180 10489
rect 14280 10480 14332 10532
rect 15292 10480 15344 10532
rect 13728 10412 13780 10464
rect 14004 10455 14056 10464
rect 14004 10421 14013 10455
rect 14013 10421 14047 10455
rect 14047 10421 14056 10455
rect 14004 10412 14056 10421
rect 14556 10412 14608 10464
rect 17132 10412 17184 10464
rect 18696 10455 18748 10464
rect 18696 10421 18705 10455
rect 18705 10421 18739 10455
rect 18739 10421 18748 10455
rect 18696 10412 18748 10421
rect 3422 10310 3474 10362
rect 3486 10310 3538 10362
rect 3550 10310 3602 10362
rect 3614 10310 3666 10362
rect 3678 10310 3730 10362
rect 8367 10310 8419 10362
rect 8431 10310 8483 10362
rect 8495 10310 8547 10362
rect 8559 10310 8611 10362
rect 8623 10310 8675 10362
rect 13312 10310 13364 10362
rect 13376 10310 13428 10362
rect 13440 10310 13492 10362
rect 13504 10310 13556 10362
rect 13568 10310 13620 10362
rect 18257 10310 18309 10362
rect 18321 10310 18373 10362
rect 18385 10310 18437 10362
rect 18449 10310 18501 10362
rect 18513 10310 18565 10362
rect 2228 10208 2280 10260
rect 7196 10208 7248 10260
rect 11612 10251 11664 10260
rect 11612 10217 11621 10251
rect 11621 10217 11655 10251
rect 11655 10217 11664 10251
rect 11612 10208 11664 10217
rect 11336 10072 11388 10124
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 1860 10047 1912 10056
rect 1860 10013 1894 10047
rect 1894 10013 1912 10047
rect 1860 10004 1912 10013
rect 3884 10004 3936 10056
rect 6828 10004 6880 10056
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 7104 10004 7156 10056
rect 9772 10004 9824 10056
rect 11428 10004 11480 10056
rect 14924 10208 14976 10260
rect 15292 10208 15344 10260
rect 18696 10208 18748 10260
rect 18880 10208 18932 10260
rect 19616 10251 19668 10260
rect 19616 10217 19625 10251
rect 19625 10217 19659 10251
rect 19659 10217 19668 10251
rect 19616 10208 19668 10217
rect 12900 10140 12952 10192
rect 13084 10140 13136 10192
rect 13820 10140 13872 10192
rect 16856 10183 16908 10192
rect 16856 10149 16865 10183
rect 16865 10149 16899 10183
rect 16899 10149 16908 10183
rect 16856 10140 16908 10149
rect 19248 10140 19300 10192
rect 13176 10072 13228 10124
rect 14556 10115 14608 10124
rect 13084 10047 13136 10056
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 14556 10081 14565 10115
rect 14565 10081 14599 10115
rect 14599 10081 14608 10115
rect 14556 10072 14608 10081
rect 14832 10072 14884 10124
rect 13084 10004 13136 10013
rect 15568 10047 15620 10056
rect 15568 10013 15577 10047
rect 15577 10013 15611 10047
rect 15611 10013 15620 10047
rect 15568 10004 15620 10013
rect 14648 9936 14700 9988
rect 16304 10004 16356 10056
rect 17868 10047 17920 10056
rect 7840 9868 7892 9920
rect 14280 9911 14332 9920
rect 14280 9877 14289 9911
rect 14289 9877 14323 9911
rect 14323 9877 14332 9911
rect 14280 9868 14332 9877
rect 15384 9868 15436 9920
rect 16672 9979 16724 9988
rect 16672 9945 16697 9979
rect 16697 9945 16724 9979
rect 17868 10013 17877 10047
rect 17877 10013 17911 10047
rect 17911 10013 17920 10047
rect 17868 10004 17920 10013
rect 18052 10047 18104 10056
rect 18052 10013 18061 10047
rect 18061 10013 18095 10047
rect 18095 10013 18104 10047
rect 18052 10004 18104 10013
rect 16672 9936 16724 9945
rect 17960 9936 18012 9988
rect 19432 9979 19484 9988
rect 19432 9945 19441 9979
rect 19441 9945 19475 9979
rect 19475 9945 19484 9979
rect 19432 9936 19484 9945
rect 17592 9911 17644 9920
rect 17592 9877 17601 9911
rect 17601 9877 17635 9911
rect 17635 9877 17644 9911
rect 17592 9868 17644 9877
rect 5894 9766 5946 9818
rect 5958 9766 6010 9818
rect 6022 9766 6074 9818
rect 6086 9766 6138 9818
rect 6150 9766 6202 9818
rect 10839 9766 10891 9818
rect 10903 9766 10955 9818
rect 10967 9766 11019 9818
rect 11031 9766 11083 9818
rect 11095 9766 11147 9818
rect 15784 9766 15836 9818
rect 15848 9766 15900 9818
rect 15912 9766 15964 9818
rect 15976 9766 16028 9818
rect 16040 9766 16092 9818
rect 20729 9766 20781 9818
rect 20793 9766 20845 9818
rect 20857 9766 20909 9818
rect 20921 9766 20973 9818
rect 20985 9766 21037 9818
rect 13084 9707 13136 9716
rect 13084 9673 13093 9707
rect 13093 9673 13127 9707
rect 13127 9673 13136 9707
rect 13084 9664 13136 9673
rect 3792 9596 3844 9648
rect 8852 9528 8904 9580
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 14188 9596 14240 9648
rect 15384 9596 15436 9648
rect 17316 9664 17368 9716
rect 16856 9639 16908 9648
rect 13728 9528 13780 9580
rect 14464 9571 14516 9580
rect 14464 9537 14473 9571
rect 14473 9537 14507 9571
rect 14507 9537 14516 9571
rect 14464 9528 14516 9537
rect 15292 9571 15344 9580
rect 1584 9460 1636 9512
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 7012 9460 7064 9512
rect 12900 9460 12952 9512
rect 15292 9537 15301 9571
rect 15301 9537 15335 9571
rect 15335 9537 15344 9571
rect 16856 9605 16865 9639
rect 16865 9605 16899 9639
rect 16899 9605 16908 9639
rect 16856 9596 16908 9605
rect 15292 9528 15344 9537
rect 16212 9528 16264 9580
rect 17592 9596 17644 9648
rect 17132 9571 17184 9580
rect 17132 9537 17141 9571
rect 17141 9537 17175 9571
rect 17175 9537 17184 9571
rect 17132 9528 17184 9537
rect 18052 9528 18104 9580
rect 18880 9571 18932 9580
rect 18880 9537 18889 9571
rect 18889 9537 18923 9571
rect 18923 9537 18932 9571
rect 18880 9528 18932 9537
rect 4620 9392 4672 9444
rect 16948 9392 17000 9444
rect 19524 9392 19576 9444
rect 6736 9324 6788 9376
rect 14096 9324 14148 9376
rect 16672 9324 16724 9376
rect 3422 9222 3474 9274
rect 3486 9222 3538 9274
rect 3550 9222 3602 9274
rect 3614 9222 3666 9274
rect 3678 9222 3730 9274
rect 8367 9222 8419 9274
rect 8431 9222 8483 9274
rect 8495 9222 8547 9274
rect 8559 9222 8611 9274
rect 8623 9222 8675 9274
rect 13312 9222 13364 9274
rect 13376 9222 13428 9274
rect 13440 9222 13492 9274
rect 13504 9222 13556 9274
rect 13568 9222 13620 9274
rect 18257 9222 18309 9274
rect 18321 9222 18373 9274
rect 18385 9222 18437 9274
rect 18449 9222 18501 9274
rect 18513 9222 18565 9274
rect 2872 9120 2924 9172
rect 6920 9120 6972 9172
rect 11520 9120 11572 9172
rect 12348 9120 12400 9172
rect 15292 9120 15344 9172
rect 18052 9120 18104 9172
rect 19892 9163 19944 9172
rect 19892 9129 19901 9163
rect 19901 9129 19935 9163
rect 19935 9129 19944 9163
rect 19892 9120 19944 9129
rect 17960 9052 18012 9104
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 7012 8984 7064 9036
rect 11428 8984 11480 9036
rect 16212 8984 16264 9036
rect 1860 8959 1912 8968
rect 1860 8925 1894 8959
rect 1894 8925 1912 8959
rect 1860 8916 1912 8925
rect 3884 8916 3936 8968
rect 4896 8959 4948 8968
rect 4896 8925 4930 8959
rect 4930 8925 4948 8959
rect 4896 8916 4948 8925
rect 8208 8916 8260 8968
rect 9772 8916 9824 8968
rect 13728 8916 13780 8968
rect 16580 8959 16632 8968
rect 16580 8925 16589 8959
rect 16589 8925 16623 8959
rect 16623 8925 16632 8959
rect 16580 8916 16632 8925
rect 16948 8959 17000 8968
rect 16948 8925 16957 8959
rect 16957 8925 16991 8959
rect 16991 8925 17000 8959
rect 16948 8916 17000 8925
rect 17040 8959 17092 8968
rect 17040 8925 17049 8959
rect 17049 8925 17083 8959
rect 17083 8925 17092 8959
rect 18052 8984 18104 9036
rect 17040 8916 17092 8925
rect 14464 8848 14516 8900
rect 18604 8916 18656 8968
rect 18880 8848 18932 8900
rect 14004 8780 14056 8832
rect 5894 8678 5946 8730
rect 5958 8678 6010 8730
rect 6022 8678 6074 8730
rect 6086 8678 6138 8730
rect 6150 8678 6202 8730
rect 10839 8678 10891 8730
rect 10903 8678 10955 8730
rect 10967 8678 11019 8730
rect 11031 8678 11083 8730
rect 11095 8678 11147 8730
rect 15784 8678 15836 8730
rect 15848 8678 15900 8730
rect 15912 8678 15964 8730
rect 15976 8678 16028 8730
rect 16040 8678 16092 8730
rect 20729 8678 20781 8730
rect 20793 8678 20845 8730
rect 20857 8678 20909 8730
rect 20921 8678 20973 8730
rect 20985 8678 21037 8730
rect 5540 8576 5592 8628
rect 16580 8576 16632 8628
rect 3240 8551 3292 8560
rect 3240 8517 3274 8551
rect 3274 8517 3292 8551
rect 3240 8508 3292 8517
rect 12900 8508 12952 8560
rect 7932 8440 7984 8492
rect 13636 8508 13688 8560
rect 16948 8508 17000 8560
rect 17960 8576 18012 8628
rect 18696 8508 18748 8560
rect 2780 8372 2832 8424
rect 9772 8415 9824 8424
rect 9772 8381 9781 8415
rect 9781 8381 9815 8415
rect 9815 8381 9824 8415
rect 9772 8372 9824 8381
rect 13728 8440 13780 8492
rect 14004 8483 14056 8492
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14004 8440 14056 8449
rect 14096 8483 14148 8492
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 15200 8440 15252 8492
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 16672 8372 16724 8424
rect 17132 8372 17184 8424
rect 18604 8483 18656 8492
rect 18604 8449 18613 8483
rect 18613 8449 18647 8483
rect 18647 8449 18656 8483
rect 18604 8440 18656 8449
rect 13176 8304 13228 8356
rect 18604 8304 18656 8356
rect 13820 8279 13872 8288
rect 13820 8245 13829 8279
rect 13829 8245 13863 8279
rect 13863 8245 13872 8279
rect 13820 8236 13872 8245
rect 18880 8304 18932 8356
rect 19616 8236 19668 8288
rect 3422 8134 3474 8186
rect 3486 8134 3538 8186
rect 3550 8134 3602 8186
rect 3614 8134 3666 8186
rect 3678 8134 3730 8186
rect 8367 8134 8419 8186
rect 8431 8134 8483 8186
rect 8495 8134 8547 8186
rect 8559 8134 8611 8186
rect 8623 8134 8675 8186
rect 13312 8134 13364 8186
rect 13376 8134 13428 8186
rect 13440 8134 13492 8186
rect 13504 8134 13556 8186
rect 13568 8134 13620 8186
rect 18257 8134 18309 8186
rect 18321 8134 18373 8186
rect 18385 8134 18437 8186
rect 18449 8134 18501 8186
rect 18513 8134 18565 8186
rect 7380 8032 7432 8084
rect 8024 8032 8076 8084
rect 14464 8032 14516 8084
rect 15200 8032 15252 8084
rect 17040 8032 17092 8084
rect 7012 7939 7064 7948
rect 7012 7905 7021 7939
rect 7021 7905 7055 7939
rect 7055 7905 7064 7939
rect 7012 7896 7064 7905
rect 9772 7896 9824 7948
rect 3884 7828 3936 7880
rect 16120 7964 16172 8016
rect 13268 7939 13320 7948
rect 13268 7905 13277 7939
rect 13277 7905 13311 7939
rect 13311 7905 13320 7939
rect 18696 7964 18748 8016
rect 18880 7964 18932 8016
rect 13268 7896 13320 7905
rect 13820 7828 13872 7880
rect 15292 7828 15344 7880
rect 15568 7871 15620 7880
rect 15568 7837 15577 7871
rect 15577 7837 15611 7871
rect 15611 7837 15620 7871
rect 15568 7828 15620 7837
rect 16948 7828 17000 7880
rect 17132 7828 17184 7880
rect 18512 7871 18564 7880
rect 9496 7760 9548 7812
rect 14280 7760 14332 7812
rect 18512 7837 18521 7871
rect 18521 7837 18555 7871
rect 18555 7837 18564 7871
rect 18512 7828 18564 7837
rect 18880 7828 18932 7880
rect 12624 7735 12676 7744
rect 12624 7701 12633 7735
rect 12633 7701 12667 7735
rect 12667 7701 12676 7735
rect 12624 7692 12676 7701
rect 13728 7692 13780 7744
rect 16856 7692 16908 7744
rect 18604 7692 18656 7744
rect 18788 7692 18840 7744
rect 19616 7692 19668 7744
rect 5894 7590 5946 7642
rect 5958 7590 6010 7642
rect 6022 7590 6074 7642
rect 6086 7590 6138 7642
rect 6150 7590 6202 7642
rect 10839 7590 10891 7642
rect 10903 7590 10955 7642
rect 10967 7590 11019 7642
rect 11031 7590 11083 7642
rect 11095 7590 11147 7642
rect 15784 7590 15836 7642
rect 15848 7590 15900 7642
rect 15912 7590 15964 7642
rect 15976 7590 16028 7642
rect 16040 7590 16092 7642
rect 20729 7590 20781 7642
rect 20793 7590 20845 7642
rect 20857 7590 20909 7642
rect 20921 7590 20973 7642
rect 20985 7590 21037 7642
rect 7012 7488 7064 7540
rect 9772 7488 9824 7540
rect 18512 7488 18564 7540
rect 2596 7395 2648 7404
rect 2596 7361 2605 7395
rect 2605 7361 2639 7395
rect 2639 7361 2648 7395
rect 2596 7352 2648 7361
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 12900 7352 12952 7404
rect 15292 7420 15344 7472
rect 14280 7352 14332 7404
rect 15200 7395 15252 7404
rect 15200 7361 15209 7395
rect 15209 7361 15243 7395
rect 15243 7361 15252 7395
rect 15200 7352 15252 7361
rect 16948 7352 17000 7404
rect 13084 7216 13136 7268
rect 13268 7284 13320 7336
rect 15292 7327 15344 7336
rect 15292 7293 15301 7327
rect 15301 7293 15335 7327
rect 15335 7293 15344 7327
rect 15292 7284 15344 7293
rect 15476 7327 15528 7336
rect 15476 7293 15485 7327
rect 15485 7293 15519 7327
rect 15519 7293 15528 7327
rect 15476 7284 15528 7293
rect 2780 7148 2832 7200
rect 3884 7191 3936 7200
rect 3884 7157 3893 7191
rect 3893 7157 3927 7191
rect 3927 7157 3936 7191
rect 3884 7148 3936 7157
rect 11704 7148 11756 7200
rect 14832 7191 14884 7200
rect 14832 7157 14841 7191
rect 14841 7157 14875 7191
rect 14875 7157 14884 7191
rect 14832 7148 14884 7157
rect 3422 7046 3474 7098
rect 3486 7046 3538 7098
rect 3550 7046 3602 7098
rect 3614 7046 3666 7098
rect 3678 7046 3730 7098
rect 8367 7046 8419 7098
rect 8431 7046 8483 7098
rect 8495 7046 8547 7098
rect 8559 7046 8611 7098
rect 8623 7046 8675 7098
rect 13312 7046 13364 7098
rect 13376 7046 13428 7098
rect 13440 7046 13492 7098
rect 13504 7046 13556 7098
rect 13568 7046 13620 7098
rect 18257 7046 18309 7098
rect 18321 7046 18373 7098
rect 18385 7046 18437 7098
rect 18449 7046 18501 7098
rect 18513 7046 18565 7098
rect 14280 6987 14332 6996
rect 14280 6953 14289 6987
rect 14289 6953 14323 6987
rect 14323 6953 14332 6987
rect 14280 6944 14332 6953
rect 15292 6944 15344 6996
rect 17408 6987 17460 6996
rect 17408 6953 17417 6987
rect 17417 6953 17451 6987
rect 17451 6953 17460 6987
rect 17408 6944 17460 6953
rect 2596 6876 2648 6928
rect 7840 6876 7892 6928
rect 14464 6876 14516 6928
rect 9772 6851 9824 6860
rect 9772 6817 9781 6851
rect 9781 6817 9815 6851
rect 9815 6817 9824 6851
rect 9772 6808 9824 6817
rect 1584 6783 1636 6792
rect 1584 6749 1593 6783
rect 1593 6749 1627 6783
rect 1627 6749 1636 6783
rect 1584 6740 1636 6749
rect 1676 6740 1728 6792
rect 14832 6808 14884 6860
rect 15384 6876 15436 6928
rect 13176 6740 13228 6792
rect 13636 6783 13688 6792
rect 5540 6672 5592 6724
rect 13636 6749 13645 6783
rect 13645 6749 13679 6783
rect 13679 6749 13688 6783
rect 13636 6740 13688 6749
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 14464 6783 14516 6792
rect 13728 6740 13780 6749
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 15568 6740 15620 6792
rect 3148 6604 3200 6656
rect 9036 6604 9088 6656
rect 10324 6604 10376 6656
rect 12992 6604 13044 6656
rect 14924 6715 14976 6724
rect 14924 6681 14933 6715
rect 14933 6681 14967 6715
rect 14967 6681 14976 6715
rect 16120 6740 16172 6792
rect 17040 6740 17092 6792
rect 18788 6808 18840 6860
rect 14924 6672 14976 6681
rect 15200 6604 15252 6656
rect 17224 6604 17276 6656
rect 17868 6740 17920 6792
rect 18604 6783 18656 6792
rect 18604 6749 18613 6783
rect 18613 6749 18647 6783
rect 18647 6749 18656 6783
rect 18604 6740 18656 6749
rect 18696 6783 18748 6792
rect 18696 6749 18705 6783
rect 18705 6749 18739 6783
rect 18739 6749 18748 6783
rect 18696 6740 18748 6749
rect 18052 6604 18104 6656
rect 18328 6647 18380 6656
rect 18328 6613 18337 6647
rect 18337 6613 18371 6647
rect 18371 6613 18380 6647
rect 18328 6604 18380 6613
rect 5894 6502 5946 6554
rect 5958 6502 6010 6554
rect 6022 6502 6074 6554
rect 6086 6502 6138 6554
rect 6150 6502 6202 6554
rect 10839 6502 10891 6554
rect 10903 6502 10955 6554
rect 10967 6502 11019 6554
rect 11031 6502 11083 6554
rect 11095 6502 11147 6554
rect 15784 6502 15836 6554
rect 15848 6502 15900 6554
rect 15912 6502 15964 6554
rect 15976 6502 16028 6554
rect 16040 6502 16092 6554
rect 20729 6502 20781 6554
rect 20793 6502 20845 6554
rect 20857 6502 20909 6554
rect 20921 6502 20973 6554
rect 20985 6502 21037 6554
rect 4252 6400 4304 6452
rect 12992 6443 13044 6452
rect 3056 6375 3108 6384
rect 3056 6341 3090 6375
rect 3090 6341 3108 6375
rect 3056 6332 3108 6341
rect 2780 6307 2832 6316
rect 2780 6273 2789 6307
rect 2789 6273 2823 6307
rect 2823 6273 2832 6307
rect 9772 6332 9824 6384
rect 12992 6409 13001 6443
rect 13001 6409 13035 6443
rect 13035 6409 13044 6443
rect 12992 6400 13044 6409
rect 15568 6400 15620 6452
rect 14464 6375 14516 6384
rect 14464 6341 14473 6375
rect 14473 6341 14507 6375
rect 14507 6341 14516 6375
rect 14464 6332 14516 6341
rect 2780 6264 2832 6273
rect 7104 6239 7156 6248
rect 7104 6205 7113 6239
rect 7113 6205 7147 6239
rect 7147 6205 7156 6239
rect 7104 6196 7156 6205
rect 10508 6264 10560 6316
rect 13728 6264 13780 6316
rect 15476 6264 15528 6316
rect 18696 6400 18748 6452
rect 17408 6332 17460 6384
rect 17224 6307 17276 6316
rect 17224 6273 17233 6307
rect 17233 6273 17267 6307
rect 17267 6273 17276 6307
rect 17224 6264 17276 6273
rect 17960 6264 18012 6316
rect 18788 6307 18840 6316
rect 18788 6273 18797 6307
rect 18797 6273 18831 6307
rect 18831 6273 18840 6307
rect 18788 6264 18840 6273
rect 18972 6307 19024 6316
rect 18972 6273 18981 6307
rect 18981 6273 19015 6307
rect 19015 6273 19024 6307
rect 18972 6264 19024 6273
rect 13084 6196 13136 6248
rect 13636 6128 13688 6180
rect 10324 6103 10376 6112
rect 10324 6069 10333 6103
rect 10333 6069 10367 6103
rect 10367 6069 10376 6103
rect 10324 6060 10376 6069
rect 11428 6060 11480 6112
rect 18328 6128 18380 6180
rect 16672 6060 16724 6112
rect 3422 5958 3474 6010
rect 3486 5958 3538 6010
rect 3550 5958 3602 6010
rect 3614 5958 3666 6010
rect 3678 5958 3730 6010
rect 8367 5958 8419 6010
rect 8431 5958 8483 6010
rect 8495 5958 8547 6010
rect 8559 5958 8611 6010
rect 8623 5958 8675 6010
rect 13312 5958 13364 6010
rect 13376 5958 13428 6010
rect 13440 5958 13492 6010
rect 13504 5958 13556 6010
rect 13568 5958 13620 6010
rect 18257 5958 18309 6010
rect 18321 5958 18373 6010
rect 18385 5958 18437 6010
rect 18449 5958 18501 6010
rect 18513 5958 18565 6010
rect 12900 5856 12952 5908
rect 14924 5856 14976 5908
rect 13728 5788 13780 5840
rect 15016 5788 15068 5840
rect 17224 5788 17276 5840
rect 18972 5788 19024 5840
rect 1584 5763 1636 5772
rect 1584 5729 1593 5763
rect 1593 5729 1627 5763
rect 1627 5729 1636 5763
rect 1584 5720 1636 5729
rect 16672 5763 16724 5772
rect 16672 5729 16681 5763
rect 16681 5729 16715 5763
rect 16715 5729 16724 5763
rect 16672 5720 16724 5729
rect 1952 5652 2004 5704
rect 2320 5652 2372 5704
rect 4528 5652 4580 5704
rect 9588 5652 9640 5704
rect 11704 5584 11756 5636
rect 14464 5652 14516 5704
rect 16120 5652 16172 5704
rect 17500 5695 17552 5704
rect 12624 5584 12676 5636
rect 5816 5516 5868 5568
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 17500 5652 17552 5661
rect 19616 5695 19668 5704
rect 18880 5584 18932 5636
rect 19616 5661 19625 5695
rect 19625 5661 19659 5695
rect 19659 5661 19668 5695
rect 19616 5652 19668 5661
rect 13728 5516 13780 5568
rect 15476 5516 15528 5568
rect 16488 5559 16540 5568
rect 16488 5525 16497 5559
rect 16497 5525 16531 5559
rect 16531 5525 16540 5559
rect 16488 5516 16540 5525
rect 5894 5414 5946 5466
rect 5958 5414 6010 5466
rect 6022 5414 6074 5466
rect 6086 5414 6138 5466
rect 6150 5414 6202 5466
rect 10839 5414 10891 5466
rect 10903 5414 10955 5466
rect 10967 5414 11019 5466
rect 11031 5414 11083 5466
rect 11095 5414 11147 5466
rect 15784 5414 15836 5466
rect 15848 5414 15900 5466
rect 15912 5414 15964 5466
rect 15976 5414 16028 5466
rect 16040 5414 16092 5466
rect 20729 5414 20781 5466
rect 20793 5414 20845 5466
rect 20857 5414 20909 5466
rect 20921 5414 20973 5466
rect 20985 5414 21037 5466
rect 7564 5312 7616 5364
rect 1584 5244 1636 5296
rect 4528 5176 4580 5228
rect 5632 5176 5684 5228
rect 15476 5244 15528 5296
rect 11428 5176 11480 5228
rect 12900 5219 12952 5228
rect 12900 5185 12909 5219
rect 12909 5185 12943 5219
rect 12943 5185 12952 5219
rect 12900 5176 12952 5185
rect 13912 5176 13964 5228
rect 9588 5108 9640 5160
rect 12808 5108 12860 5160
rect 14280 5108 14332 5160
rect 15016 5176 15068 5228
rect 15200 5219 15252 5228
rect 15200 5185 15209 5219
rect 15209 5185 15243 5219
rect 15243 5185 15252 5219
rect 15200 5176 15252 5185
rect 14832 5108 14884 5160
rect 15384 5219 15436 5228
rect 15384 5185 15393 5219
rect 15393 5185 15427 5219
rect 15427 5185 15436 5219
rect 17500 5312 17552 5364
rect 15384 5176 15436 5185
rect 17040 5176 17092 5228
rect 2780 5083 2832 5092
rect 2780 5049 2789 5083
rect 2789 5049 2823 5083
rect 2823 5049 2832 5083
rect 11152 5083 11204 5092
rect 2780 5040 2832 5049
rect 11152 5049 11161 5083
rect 11161 5049 11195 5083
rect 11195 5049 11204 5083
rect 11152 5040 11204 5049
rect 11244 5040 11296 5092
rect 5816 4972 5868 5024
rect 12624 4972 12676 5024
rect 3422 4870 3474 4922
rect 3486 4870 3538 4922
rect 3550 4870 3602 4922
rect 3614 4870 3666 4922
rect 3678 4870 3730 4922
rect 8367 4870 8419 4922
rect 8431 4870 8483 4922
rect 8495 4870 8547 4922
rect 8559 4870 8611 4922
rect 8623 4870 8675 4922
rect 13312 4870 13364 4922
rect 13376 4870 13428 4922
rect 13440 4870 13492 4922
rect 13504 4870 13556 4922
rect 13568 4870 13620 4922
rect 18257 4870 18309 4922
rect 18321 4870 18373 4922
rect 18385 4870 18437 4922
rect 18449 4870 18501 4922
rect 18513 4870 18565 4922
rect 1584 4632 1636 4684
rect 4528 4632 4580 4684
rect 7104 4675 7156 4684
rect 7104 4641 7113 4675
rect 7113 4641 7147 4675
rect 7147 4641 7156 4675
rect 7104 4632 7156 4641
rect 12624 4768 12676 4820
rect 14648 4768 14700 4820
rect 15384 4768 15436 4820
rect 9588 4564 9640 4616
rect 14924 4700 14976 4752
rect 15108 4700 15160 4752
rect 15200 4632 15252 4684
rect 19616 4700 19668 4752
rect 12808 4564 12860 4616
rect 14648 4607 14700 4616
rect 14648 4573 14657 4607
rect 14657 4573 14691 4607
rect 14691 4573 14700 4607
rect 14648 4564 14700 4573
rect 15384 4564 15436 4616
rect 3976 4496 4028 4548
rect 9864 4496 9916 4548
rect 14740 4496 14792 4548
rect 17500 4632 17552 4684
rect 16672 4564 16724 4616
rect 17224 4607 17276 4616
rect 17224 4573 17233 4607
rect 17233 4573 17267 4607
rect 17267 4573 17276 4607
rect 17224 4564 17276 4573
rect 18052 4607 18104 4616
rect 18052 4573 18061 4607
rect 18061 4573 18095 4607
rect 18095 4573 18104 4607
rect 18052 4564 18104 4573
rect 16856 4496 16908 4548
rect 4804 4428 4856 4480
rect 6644 4471 6696 4480
rect 6644 4437 6653 4471
rect 6653 4437 6687 4471
rect 6687 4437 6696 4471
rect 6644 4428 6696 4437
rect 10416 4428 10468 4480
rect 17132 4428 17184 4480
rect 5894 4326 5946 4378
rect 5958 4326 6010 4378
rect 6022 4326 6074 4378
rect 6086 4326 6138 4378
rect 6150 4326 6202 4378
rect 10839 4326 10891 4378
rect 10903 4326 10955 4378
rect 10967 4326 11019 4378
rect 11031 4326 11083 4378
rect 11095 4326 11147 4378
rect 15784 4326 15836 4378
rect 15848 4326 15900 4378
rect 15912 4326 15964 4378
rect 15976 4326 16028 4378
rect 16040 4326 16092 4378
rect 20729 4326 20781 4378
rect 20793 4326 20845 4378
rect 20857 4326 20909 4378
rect 20921 4326 20973 4378
rect 20985 4326 21037 4378
rect 9864 4224 9916 4276
rect 12992 4224 13044 4276
rect 16948 4224 17000 4276
rect 6644 4156 6696 4208
rect 12900 4156 12952 4208
rect 13728 4156 13780 4208
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 1860 4131 1912 4140
rect 1860 4097 1894 4131
rect 1894 4097 1912 4131
rect 4528 4131 4580 4140
rect 1860 4088 1912 4097
rect 4528 4097 4537 4131
rect 4537 4097 4571 4131
rect 4571 4097 4580 4131
rect 4528 4088 4580 4097
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 9680 4088 9732 4140
rect 11704 4088 11756 4140
rect 14832 4131 14884 4140
rect 7012 4020 7064 4072
rect 9588 4063 9640 4072
rect 9588 4029 9597 4063
rect 9597 4029 9631 4063
rect 9631 4029 9640 4063
rect 9588 4020 9640 4029
rect 14832 4097 14841 4131
rect 14841 4097 14875 4131
rect 14875 4097 14884 4131
rect 14832 4088 14884 4097
rect 15016 4131 15068 4140
rect 15016 4097 15025 4131
rect 15025 4097 15059 4131
rect 15059 4097 15068 4131
rect 15016 4088 15068 4097
rect 16856 4131 16908 4140
rect 16856 4097 16865 4131
rect 16865 4097 16899 4131
rect 16899 4097 16908 4131
rect 16856 4088 16908 4097
rect 17132 4088 17184 4140
rect 14556 4020 14608 4072
rect 1952 3884 2004 3936
rect 8208 3884 8260 3936
rect 11796 3884 11848 3936
rect 14924 3952 14976 4004
rect 17316 4020 17368 4072
rect 16488 3884 16540 3936
rect 17040 3884 17092 3936
rect 3422 3782 3474 3834
rect 3486 3782 3538 3834
rect 3550 3782 3602 3834
rect 3614 3782 3666 3834
rect 3678 3782 3730 3834
rect 8367 3782 8419 3834
rect 8431 3782 8483 3834
rect 8495 3782 8547 3834
rect 8559 3782 8611 3834
rect 8623 3782 8675 3834
rect 13312 3782 13364 3834
rect 13376 3782 13428 3834
rect 13440 3782 13492 3834
rect 13504 3782 13556 3834
rect 13568 3782 13620 3834
rect 18257 3782 18309 3834
rect 18321 3782 18373 3834
rect 18385 3782 18437 3834
rect 18449 3782 18501 3834
rect 18513 3782 18565 3834
rect 3148 3680 3200 3732
rect 5540 3680 5592 3732
rect 9680 3680 9732 3732
rect 12992 3723 13044 3732
rect 1584 3544 1636 3596
rect 8208 3544 8260 3596
rect 11888 3612 11940 3664
rect 12992 3689 13001 3723
rect 13001 3689 13035 3723
rect 13035 3689 13044 3723
rect 12992 3680 13044 3689
rect 14648 3680 14700 3732
rect 17224 3723 17276 3732
rect 17224 3689 17233 3723
rect 17233 3689 17267 3723
rect 17267 3689 17276 3723
rect 17224 3680 17276 3689
rect 7104 3476 7156 3528
rect 9588 3476 9640 3528
rect 12808 3544 12860 3596
rect 2964 3408 3016 3460
rect 9772 3408 9824 3460
rect 3332 3340 3384 3392
rect 4804 3340 4856 3392
rect 6736 3340 6788 3392
rect 8760 3340 8812 3392
rect 11244 3476 11296 3528
rect 11796 3519 11848 3528
rect 11796 3485 11805 3519
rect 11805 3485 11839 3519
rect 11839 3485 11848 3519
rect 11796 3476 11848 3485
rect 11980 3519 12032 3528
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 12072 3519 12124 3528
rect 12072 3485 12081 3519
rect 12081 3485 12115 3519
rect 12115 3485 12124 3519
rect 15016 3544 15068 3596
rect 12072 3476 12124 3485
rect 10416 3408 10468 3460
rect 13360 3519 13412 3528
rect 13360 3485 13369 3519
rect 13369 3485 13403 3519
rect 13403 3485 13412 3519
rect 13360 3476 13412 3485
rect 13728 3476 13780 3528
rect 14924 3519 14976 3528
rect 14924 3485 14933 3519
rect 14933 3485 14967 3519
rect 14967 3485 14976 3519
rect 14924 3476 14976 3485
rect 16304 3476 16356 3528
rect 17040 3519 17092 3528
rect 17040 3485 17049 3519
rect 17049 3485 17083 3519
rect 17083 3485 17092 3519
rect 17316 3519 17368 3528
rect 17040 3476 17092 3485
rect 17316 3485 17325 3519
rect 17325 3485 17359 3519
rect 17359 3485 17368 3519
rect 17316 3476 17368 3485
rect 17960 3519 18012 3528
rect 17960 3485 17969 3519
rect 17969 3485 18003 3519
rect 18003 3485 18012 3519
rect 17960 3476 18012 3485
rect 18052 3519 18104 3528
rect 18052 3485 18061 3519
rect 18061 3485 18095 3519
rect 18095 3485 18104 3519
rect 18052 3476 18104 3485
rect 14188 3408 14240 3460
rect 14556 3408 14608 3460
rect 16856 3408 16908 3460
rect 15384 3340 15436 3392
rect 17776 3383 17828 3392
rect 17776 3349 17785 3383
rect 17785 3349 17819 3383
rect 17819 3349 17828 3383
rect 17776 3340 17828 3349
rect 5894 3238 5946 3290
rect 5958 3238 6010 3290
rect 6022 3238 6074 3290
rect 6086 3238 6138 3290
rect 6150 3238 6202 3290
rect 10839 3238 10891 3290
rect 10903 3238 10955 3290
rect 10967 3238 11019 3290
rect 11031 3238 11083 3290
rect 11095 3238 11147 3290
rect 15784 3238 15836 3290
rect 15848 3238 15900 3290
rect 15912 3238 15964 3290
rect 15976 3238 16028 3290
rect 16040 3238 16092 3290
rect 20729 3238 20781 3290
rect 20793 3238 20845 3290
rect 20857 3238 20909 3290
rect 20921 3238 20973 3290
rect 20985 3238 21037 3290
rect 1860 3179 1912 3188
rect 1860 3145 1869 3179
rect 1869 3145 1903 3179
rect 1903 3145 1912 3179
rect 1860 3136 1912 3145
rect 3332 3136 3384 3188
rect 2596 3111 2648 3120
rect 2596 3077 2605 3111
rect 2605 3077 2639 3111
rect 2639 3077 2648 3111
rect 2596 3068 2648 3077
rect 4528 3068 4580 3120
rect 4804 3111 4856 3120
rect 4804 3077 4813 3111
rect 4813 3077 4847 3111
rect 4847 3077 4856 3111
rect 4804 3068 4856 3077
rect 5632 3136 5684 3188
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 2320 2932 2372 2984
rect 4896 2932 4948 2984
rect 5632 3000 5684 3052
rect 7656 3136 7708 3188
rect 9772 3136 9824 3188
rect 13360 3136 13412 3188
rect 13636 3179 13688 3188
rect 13636 3145 13645 3179
rect 13645 3145 13679 3179
rect 13679 3145 13688 3179
rect 13636 3136 13688 3145
rect 14188 3179 14240 3188
rect 14188 3145 14197 3179
rect 14197 3145 14231 3179
rect 14231 3145 14240 3179
rect 14188 3136 14240 3145
rect 5816 3000 5868 3052
rect 7840 3111 7892 3120
rect 6736 3043 6788 3052
rect 6736 3009 6745 3043
rect 6745 3009 6779 3043
rect 6779 3009 6788 3043
rect 6736 3000 6788 3009
rect 5724 2864 5776 2916
rect 7840 3077 7849 3111
rect 7849 3077 7883 3111
rect 7883 3077 7892 3111
rect 7840 3068 7892 3077
rect 9588 3111 9640 3120
rect 9588 3077 9597 3111
rect 9597 3077 9631 3111
rect 9631 3077 9640 3111
rect 9588 3068 9640 3077
rect 12072 3068 12124 3120
rect 10232 3043 10284 3052
rect 10232 3009 10241 3043
rect 10241 3009 10275 3043
rect 10275 3009 10284 3043
rect 10232 3000 10284 3009
rect 11796 3000 11848 3052
rect 7288 2975 7340 2984
rect 7288 2941 7297 2975
rect 7297 2941 7331 2975
rect 7331 2941 7340 2975
rect 7288 2932 7340 2941
rect 8760 2932 8812 2984
rect 11980 2932 12032 2984
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 14924 3043 14976 3052
rect 14924 3009 14933 3043
rect 14933 3009 14967 3043
rect 14967 3009 14976 3043
rect 14924 3000 14976 3009
rect 15292 3000 15344 3052
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 7012 2864 7064 2916
rect 13176 2864 13228 2916
rect 4804 2839 4856 2848
rect 4804 2805 4813 2839
rect 4813 2805 4847 2839
rect 4847 2805 4856 2839
rect 4804 2796 4856 2805
rect 5632 2796 5684 2848
rect 5908 2839 5960 2848
rect 5908 2805 5917 2839
rect 5917 2805 5951 2839
rect 5951 2805 5960 2839
rect 5908 2796 5960 2805
rect 8852 2796 8904 2848
rect 12072 2796 12124 2848
rect 14832 2932 14884 2984
rect 15016 2932 15068 2984
rect 16304 3068 16356 3120
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 17316 2932 17368 2984
rect 18052 2932 18104 2984
rect 13452 2864 13504 2916
rect 14556 2796 14608 2848
rect 3422 2694 3474 2746
rect 3486 2694 3538 2746
rect 3550 2694 3602 2746
rect 3614 2694 3666 2746
rect 3678 2694 3730 2746
rect 8367 2694 8419 2746
rect 8431 2694 8483 2746
rect 8495 2694 8547 2746
rect 8559 2694 8611 2746
rect 8623 2694 8675 2746
rect 13312 2694 13364 2746
rect 13376 2694 13428 2746
rect 13440 2694 13492 2746
rect 13504 2694 13556 2746
rect 13568 2694 13620 2746
rect 18257 2694 18309 2746
rect 18321 2694 18373 2746
rect 18385 2694 18437 2746
rect 18449 2694 18501 2746
rect 18513 2694 18565 2746
rect 2964 2635 3016 2644
rect 2964 2601 2973 2635
rect 2973 2601 3007 2635
rect 3007 2601 3016 2635
rect 2964 2592 3016 2601
rect 3332 2635 3384 2644
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 3976 2635 4028 2644
rect 3976 2601 3985 2635
rect 3985 2601 4019 2635
rect 4019 2601 4028 2635
rect 3976 2592 4028 2601
rect 5632 2635 5684 2644
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 7656 2635 7708 2644
rect 7656 2601 7665 2635
rect 7665 2601 7699 2635
rect 7699 2601 7708 2635
rect 7656 2592 7708 2601
rect 10232 2592 10284 2644
rect 2320 2524 2372 2576
rect 2320 2388 2372 2440
rect 3332 2320 3384 2372
rect 1952 2252 2004 2304
rect 5908 2524 5960 2576
rect 4804 2456 4856 2508
rect 7288 2456 7340 2508
rect 9588 2499 9640 2508
rect 9588 2465 9597 2499
rect 9597 2465 9631 2499
rect 9631 2465 9640 2499
rect 9588 2456 9640 2465
rect 4988 2320 5040 2372
rect 5724 2320 5776 2372
rect 8852 2388 8904 2440
rect 11704 2524 11756 2576
rect 13636 2524 13688 2576
rect 14924 2592 14976 2644
rect 11888 2431 11940 2440
rect 11888 2397 11897 2431
rect 11897 2397 11931 2431
rect 11931 2397 11940 2431
rect 11888 2388 11940 2397
rect 8760 2320 8812 2372
rect 17776 2456 17828 2508
rect 14280 2388 14332 2440
rect 15292 2431 15344 2440
rect 15292 2397 15301 2431
rect 15301 2397 15335 2431
rect 15335 2397 15344 2431
rect 15292 2388 15344 2397
rect 16856 2320 16908 2372
rect 14280 2252 14332 2304
rect 15384 2252 15436 2304
rect 5894 2150 5946 2202
rect 5958 2150 6010 2202
rect 6022 2150 6074 2202
rect 6086 2150 6138 2202
rect 6150 2150 6202 2202
rect 10839 2150 10891 2202
rect 10903 2150 10955 2202
rect 10967 2150 11019 2202
rect 11031 2150 11083 2202
rect 11095 2150 11147 2202
rect 15784 2150 15836 2202
rect 15848 2150 15900 2202
rect 15912 2150 15964 2202
rect 15976 2150 16028 2202
rect 16040 2150 16092 2202
rect 20729 2150 20781 2202
rect 20793 2150 20845 2202
rect 20857 2150 20909 2202
rect 20921 2150 20973 2202
rect 20985 2150 21037 2202
<< metal2 >>
rect 5894 19612 6202 19621
rect 5894 19610 5900 19612
rect 5956 19610 5980 19612
rect 6036 19610 6060 19612
rect 6116 19610 6140 19612
rect 6196 19610 6202 19612
rect 5956 19558 5958 19610
rect 6138 19558 6140 19610
rect 5894 19556 5900 19558
rect 5956 19556 5980 19558
rect 6036 19556 6060 19558
rect 6116 19556 6140 19558
rect 6196 19556 6202 19558
rect 5894 19547 6202 19556
rect 10839 19612 11147 19621
rect 10839 19610 10845 19612
rect 10901 19610 10925 19612
rect 10981 19610 11005 19612
rect 11061 19610 11085 19612
rect 11141 19610 11147 19612
rect 10901 19558 10903 19610
rect 11083 19558 11085 19610
rect 10839 19556 10845 19558
rect 10901 19556 10925 19558
rect 10981 19556 11005 19558
rect 11061 19556 11085 19558
rect 11141 19556 11147 19558
rect 10839 19547 11147 19556
rect 15784 19612 16092 19621
rect 15784 19610 15790 19612
rect 15846 19610 15870 19612
rect 15926 19610 15950 19612
rect 16006 19610 16030 19612
rect 16086 19610 16092 19612
rect 15846 19558 15848 19610
rect 16028 19558 16030 19610
rect 15784 19556 15790 19558
rect 15846 19556 15870 19558
rect 15926 19556 15950 19558
rect 16006 19556 16030 19558
rect 16086 19556 16092 19558
rect 15784 19547 16092 19556
rect 20729 19612 21037 19621
rect 20729 19610 20735 19612
rect 20791 19610 20815 19612
rect 20871 19610 20895 19612
rect 20951 19610 20975 19612
rect 21031 19610 21037 19612
rect 20791 19558 20793 19610
rect 20973 19558 20975 19610
rect 20729 19556 20735 19558
rect 20791 19556 20815 19558
rect 20871 19556 20895 19558
rect 20951 19556 20975 19558
rect 21031 19556 21037 19558
rect 20729 19547 21037 19556
rect 3422 19068 3730 19077
rect 3422 19066 3428 19068
rect 3484 19066 3508 19068
rect 3564 19066 3588 19068
rect 3644 19066 3668 19068
rect 3724 19066 3730 19068
rect 3484 19014 3486 19066
rect 3666 19014 3668 19066
rect 3422 19012 3428 19014
rect 3484 19012 3508 19014
rect 3564 19012 3588 19014
rect 3644 19012 3668 19014
rect 3724 19012 3730 19014
rect 3422 19003 3730 19012
rect 8367 19068 8675 19077
rect 8367 19066 8373 19068
rect 8429 19066 8453 19068
rect 8509 19066 8533 19068
rect 8589 19066 8613 19068
rect 8669 19066 8675 19068
rect 8429 19014 8431 19066
rect 8611 19014 8613 19066
rect 8367 19012 8373 19014
rect 8429 19012 8453 19014
rect 8509 19012 8533 19014
rect 8589 19012 8613 19014
rect 8669 19012 8675 19014
rect 8367 19003 8675 19012
rect 13312 19068 13620 19077
rect 13312 19066 13318 19068
rect 13374 19066 13398 19068
rect 13454 19066 13478 19068
rect 13534 19066 13558 19068
rect 13614 19066 13620 19068
rect 13374 19014 13376 19066
rect 13556 19014 13558 19066
rect 13312 19012 13318 19014
rect 13374 19012 13398 19014
rect 13454 19012 13478 19014
rect 13534 19012 13558 19014
rect 13614 19012 13620 19014
rect 13312 19003 13620 19012
rect 18257 19068 18565 19077
rect 18257 19066 18263 19068
rect 18319 19066 18343 19068
rect 18399 19066 18423 19068
rect 18479 19066 18503 19068
rect 18559 19066 18565 19068
rect 18319 19014 18321 19066
rect 18501 19014 18503 19066
rect 18257 19012 18263 19014
rect 18319 19012 18343 19014
rect 18399 19012 18423 19014
rect 18479 19012 18503 19014
rect 18559 19012 18565 19014
rect 18257 19003 18565 19012
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 1860 18692 1912 18698
rect 1860 18634 1912 18640
rect 1872 18329 1900 18634
rect 1858 18320 1914 18329
rect 1858 18255 1914 18264
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 2228 15360 2280 15366
rect 2228 15302 2280 15308
rect 1964 14074 1992 15302
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2056 14346 2084 14962
rect 2240 14958 2268 15302
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2240 14346 2268 14894
rect 2044 14340 2096 14346
rect 2044 14282 2096 14288
rect 2228 14340 2280 14346
rect 2228 14282 2280 14288
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2056 13938 2084 14282
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1596 10282 1624 13670
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2056 12782 2084 13262
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1674 10976 1730 10985
rect 1674 10911 1730 10920
rect 1688 10742 1716 10911
rect 1676 10736 1728 10742
rect 1676 10678 1728 10684
rect 1596 10254 1716 10282
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1596 9518 1624 9998
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1596 9042 1624 9454
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1688 6798 1716 10254
rect 1872 10062 1900 12038
rect 1952 11280 2004 11286
rect 1952 11222 2004 11228
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1860 8968 1912 8974
rect 1964 8956 1992 11222
rect 1912 8928 1992 8956
rect 1860 8910 1912 8916
rect 2056 6914 2084 12718
rect 2240 12102 2268 14282
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2240 10266 2268 12038
rect 2332 11898 2360 18702
rect 5894 18524 6202 18533
rect 5894 18522 5900 18524
rect 5956 18522 5980 18524
rect 6036 18522 6060 18524
rect 6116 18522 6140 18524
rect 6196 18522 6202 18524
rect 5956 18470 5958 18522
rect 6138 18470 6140 18522
rect 5894 18468 5900 18470
rect 5956 18468 5980 18470
rect 6036 18468 6060 18470
rect 6116 18468 6140 18470
rect 6196 18468 6202 18470
rect 5894 18459 6202 18468
rect 10839 18524 11147 18533
rect 10839 18522 10845 18524
rect 10901 18522 10925 18524
rect 10981 18522 11005 18524
rect 11061 18522 11085 18524
rect 11141 18522 11147 18524
rect 10901 18470 10903 18522
rect 11083 18470 11085 18522
rect 10839 18468 10845 18470
rect 10901 18468 10925 18470
rect 10981 18468 11005 18470
rect 11061 18468 11085 18470
rect 11141 18468 11147 18470
rect 10839 18459 11147 18468
rect 15784 18524 16092 18533
rect 15784 18522 15790 18524
rect 15846 18522 15870 18524
rect 15926 18522 15950 18524
rect 16006 18522 16030 18524
rect 16086 18522 16092 18524
rect 15846 18470 15848 18522
rect 16028 18470 16030 18522
rect 15784 18468 15790 18470
rect 15846 18468 15870 18470
rect 15926 18468 15950 18470
rect 16006 18468 16030 18470
rect 16086 18468 16092 18470
rect 15784 18459 16092 18468
rect 20729 18524 21037 18533
rect 20729 18522 20735 18524
rect 20791 18522 20815 18524
rect 20871 18522 20895 18524
rect 20951 18522 20975 18524
rect 21031 18522 21037 18524
rect 20791 18470 20793 18522
rect 20973 18470 20975 18522
rect 20729 18468 20735 18470
rect 20791 18468 20815 18470
rect 20871 18468 20895 18470
rect 20951 18468 20975 18470
rect 21031 18468 21037 18470
rect 20729 18459 21037 18468
rect 3422 17980 3730 17989
rect 3422 17978 3428 17980
rect 3484 17978 3508 17980
rect 3564 17978 3588 17980
rect 3644 17978 3668 17980
rect 3724 17978 3730 17980
rect 3484 17926 3486 17978
rect 3666 17926 3668 17978
rect 3422 17924 3428 17926
rect 3484 17924 3508 17926
rect 3564 17924 3588 17926
rect 3644 17924 3668 17926
rect 3724 17924 3730 17926
rect 3422 17915 3730 17924
rect 8367 17980 8675 17989
rect 8367 17978 8373 17980
rect 8429 17978 8453 17980
rect 8509 17978 8533 17980
rect 8589 17978 8613 17980
rect 8669 17978 8675 17980
rect 8429 17926 8431 17978
rect 8611 17926 8613 17978
rect 8367 17924 8373 17926
rect 8429 17924 8453 17926
rect 8509 17924 8533 17926
rect 8589 17924 8613 17926
rect 8669 17924 8675 17926
rect 8367 17915 8675 17924
rect 13312 17980 13620 17989
rect 13312 17978 13318 17980
rect 13374 17978 13398 17980
rect 13454 17978 13478 17980
rect 13534 17978 13558 17980
rect 13614 17978 13620 17980
rect 13374 17926 13376 17978
rect 13556 17926 13558 17978
rect 13312 17924 13318 17926
rect 13374 17924 13398 17926
rect 13454 17924 13478 17926
rect 13534 17924 13558 17926
rect 13614 17924 13620 17926
rect 13312 17915 13620 17924
rect 18257 17980 18565 17989
rect 18257 17978 18263 17980
rect 18319 17978 18343 17980
rect 18399 17978 18423 17980
rect 18479 17978 18503 17980
rect 18559 17978 18565 17980
rect 18319 17926 18321 17978
rect 18501 17926 18503 17978
rect 18257 17924 18263 17926
rect 18319 17924 18343 17926
rect 18399 17924 18423 17926
rect 18479 17924 18503 17926
rect 18559 17924 18565 17926
rect 18257 17915 18565 17924
rect 5894 17436 6202 17445
rect 5894 17434 5900 17436
rect 5956 17434 5980 17436
rect 6036 17434 6060 17436
rect 6116 17434 6140 17436
rect 6196 17434 6202 17436
rect 5956 17382 5958 17434
rect 6138 17382 6140 17434
rect 5894 17380 5900 17382
rect 5956 17380 5980 17382
rect 6036 17380 6060 17382
rect 6116 17380 6140 17382
rect 6196 17380 6202 17382
rect 5894 17371 6202 17380
rect 10839 17436 11147 17445
rect 10839 17434 10845 17436
rect 10901 17434 10925 17436
rect 10981 17434 11005 17436
rect 11061 17434 11085 17436
rect 11141 17434 11147 17436
rect 10901 17382 10903 17434
rect 11083 17382 11085 17434
rect 10839 17380 10845 17382
rect 10901 17380 10925 17382
rect 10981 17380 11005 17382
rect 11061 17380 11085 17382
rect 11141 17380 11147 17382
rect 10839 17371 11147 17380
rect 15784 17436 16092 17445
rect 15784 17434 15790 17436
rect 15846 17434 15870 17436
rect 15926 17434 15950 17436
rect 16006 17434 16030 17436
rect 16086 17434 16092 17436
rect 15846 17382 15848 17434
rect 16028 17382 16030 17434
rect 15784 17380 15790 17382
rect 15846 17380 15870 17382
rect 15926 17380 15950 17382
rect 16006 17380 16030 17382
rect 16086 17380 16092 17382
rect 15784 17371 16092 17380
rect 20729 17436 21037 17445
rect 20729 17434 20735 17436
rect 20791 17434 20815 17436
rect 20871 17434 20895 17436
rect 20951 17434 20975 17436
rect 21031 17434 21037 17436
rect 20791 17382 20793 17434
rect 20973 17382 20975 17434
rect 20729 17380 20735 17382
rect 20791 17380 20815 17382
rect 20871 17380 20895 17382
rect 20951 17380 20975 17382
rect 21031 17380 21037 17382
rect 20729 17371 21037 17380
rect 5632 17264 5684 17270
rect 5632 17206 5684 17212
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 4988 17060 5040 17066
rect 4988 17002 5040 17008
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 3422 16892 3730 16901
rect 3422 16890 3428 16892
rect 3484 16890 3508 16892
rect 3564 16890 3588 16892
rect 3644 16890 3668 16892
rect 3724 16890 3730 16892
rect 3484 16838 3486 16890
rect 3666 16838 3668 16890
rect 3422 16836 3428 16838
rect 3484 16836 3508 16838
rect 3564 16836 3588 16838
rect 3644 16836 3668 16838
rect 3724 16836 3730 16838
rect 3422 16827 3730 16836
rect 4540 16590 4568 16934
rect 5000 16726 5028 17002
rect 4988 16720 5040 16726
rect 4988 16662 5040 16668
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 3240 16448 3292 16454
rect 3240 16390 3292 16396
rect 3148 15564 3200 15570
rect 3148 15506 3200 15512
rect 3160 15314 3188 15506
rect 3252 15502 3280 16390
rect 3344 16250 3372 16526
rect 4712 16516 4764 16522
rect 4712 16458 4764 16464
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 4724 16114 4752 16458
rect 5000 16114 5028 16662
rect 5552 16658 5580 17138
rect 5644 17134 5672 17206
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 5644 16794 5672 17070
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 3792 15904 3844 15910
rect 3792 15846 3844 15852
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 3422 15804 3730 15813
rect 3422 15802 3428 15804
rect 3484 15802 3508 15804
rect 3564 15802 3588 15804
rect 3644 15802 3668 15804
rect 3724 15802 3730 15804
rect 3484 15750 3486 15802
rect 3666 15750 3668 15802
rect 3422 15748 3428 15750
rect 3484 15748 3508 15750
rect 3564 15748 3588 15750
rect 3644 15748 3668 15750
rect 3724 15748 3730 15750
rect 3422 15739 3730 15748
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3160 15286 3280 15314
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 3068 14414 3096 14554
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2424 14006 2452 14214
rect 2412 14000 2464 14006
rect 2412 13942 2464 13948
rect 2792 11898 2820 14214
rect 3160 13938 3188 14758
rect 3252 14346 3280 15286
rect 3422 14716 3730 14725
rect 3422 14714 3428 14716
rect 3484 14714 3508 14716
rect 3564 14714 3588 14716
rect 3644 14714 3668 14716
rect 3724 14714 3730 14716
rect 3484 14662 3486 14714
rect 3666 14662 3668 14714
rect 3422 14660 3428 14662
rect 3484 14660 3508 14662
rect 3564 14660 3588 14662
rect 3644 14660 3668 14662
rect 3724 14660 3730 14662
rect 3422 14651 3730 14660
rect 3804 14618 3832 15846
rect 3884 14884 3936 14890
rect 3884 14826 3936 14832
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 3896 14414 3924 14826
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 4172 14414 4200 14486
rect 3332 14408 3384 14414
rect 3332 14350 3384 14356
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 3240 14340 3292 14346
rect 3240 14282 3292 14288
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 3252 13870 3280 14282
rect 3344 14074 3372 14350
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 2964 13864 3016 13870
rect 3240 13864 3292 13870
rect 3016 13812 3188 13818
rect 2964 13806 3188 13812
rect 3436 13818 3464 14350
rect 3240 13806 3292 13812
rect 2872 13796 2924 13802
rect 2976 13790 3188 13806
rect 2872 13738 2924 13744
rect 2884 13258 2912 13738
rect 2964 13456 3016 13462
rect 2964 13398 3016 13404
rect 2872 13252 2924 13258
rect 2872 13194 2924 13200
rect 2976 12306 3004 13398
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2792 11014 2820 11698
rect 2884 11694 2912 12174
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2884 11082 2912 11630
rect 2976 11150 3004 12242
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2792 8430 2820 9454
rect 2884 9178 2912 11018
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2608 6934 2636 7346
rect 2792 7206 2820 8366
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 1964 6886 2084 6914
rect 2596 6928 2648 6934
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1596 5778 1624 6734
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1596 5302 1624 5714
rect 1964 5710 1992 6886
rect 2596 6870 2648 6876
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 1584 5296 1636 5302
rect 1584 5238 1636 5244
rect 1596 4690 1624 5238
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 1596 4146 1624 4626
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1596 3602 1624 4082
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1872 3194 1900 4082
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 1964 3058 1992 3878
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 1964 2310 1992 2994
rect 2332 2990 2360 5646
rect 2608 3126 2636 6870
rect 2792 6322 2820 7142
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2976 5137 3004 10950
rect 3068 6390 3096 12582
rect 3160 6662 3188 13790
rect 3252 13462 3280 13806
rect 3344 13790 3464 13818
rect 3240 13456 3292 13462
rect 3240 13398 3292 13404
rect 3344 12850 3372 13790
rect 3422 13628 3730 13637
rect 3422 13626 3428 13628
rect 3484 13626 3508 13628
rect 3564 13626 3588 13628
rect 3644 13626 3668 13628
rect 3724 13626 3730 13628
rect 3484 13574 3486 13626
rect 3666 13574 3668 13626
rect 3422 13572 3428 13574
rect 3484 13572 3508 13574
rect 3564 13572 3588 13574
rect 3644 13572 3668 13574
rect 3724 13572 3730 13574
rect 3422 13563 3730 13572
rect 4724 13394 4752 15846
rect 5000 14550 5028 16050
rect 5184 16046 5212 16390
rect 5644 16114 5672 16730
rect 6104 16658 6132 16934
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 5736 16250 5764 16526
rect 5816 16448 5868 16454
rect 5816 16390 5868 16396
rect 5724 16244 5776 16250
rect 5724 16186 5776 16192
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 5080 15972 5132 15978
rect 5080 15914 5132 15920
rect 4988 14544 5040 14550
rect 4988 14486 5040 14492
rect 5092 14414 5120 15914
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5080 14408 5132 14414
rect 5080 14350 5132 14356
rect 5092 14278 5120 14350
rect 5172 14340 5224 14346
rect 5172 14282 5224 14288
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 5184 14074 5212 14282
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3344 12434 3372 12786
rect 4080 12714 4108 13194
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4172 12986 4200 13126
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4252 12912 4304 12918
rect 4252 12854 4304 12860
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 3422 12540 3730 12549
rect 3422 12538 3428 12540
rect 3484 12538 3508 12540
rect 3564 12538 3588 12540
rect 3644 12538 3668 12540
rect 3724 12538 3730 12540
rect 3484 12486 3486 12538
rect 3666 12486 3668 12538
rect 3422 12484 3428 12486
rect 3484 12484 3508 12486
rect 3564 12484 3588 12486
rect 3644 12484 3668 12486
rect 3724 12484 3730 12486
rect 3422 12475 3730 12484
rect 4080 12442 4108 12650
rect 3252 12406 3372 12434
rect 4068 12436 4120 12442
rect 3252 11762 3280 12406
rect 4068 12378 4120 12384
rect 4080 12306 4108 12378
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3252 8566 3280 11494
rect 3344 11218 3372 12038
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3422 11452 3730 11461
rect 3422 11450 3428 11452
rect 3484 11450 3508 11452
rect 3564 11450 3588 11452
rect 3644 11450 3668 11452
rect 3724 11450 3730 11452
rect 3484 11398 3486 11450
rect 3666 11398 3668 11450
rect 3422 11396 3428 11398
rect 3484 11396 3508 11398
rect 3564 11396 3588 11398
rect 3644 11396 3668 11398
rect 3724 11396 3730 11398
rect 3422 11387 3730 11396
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3422 10364 3730 10373
rect 3422 10362 3428 10364
rect 3484 10362 3508 10364
rect 3564 10362 3588 10364
rect 3644 10362 3668 10364
rect 3724 10362 3730 10364
rect 3484 10310 3486 10362
rect 3666 10310 3668 10362
rect 3422 10308 3428 10310
rect 3484 10308 3508 10310
rect 3564 10308 3588 10310
rect 3644 10308 3668 10310
rect 3724 10308 3730 10310
rect 3422 10299 3730 10308
rect 3804 9654 3832 11494
rect 3896 11218 3924 11698
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3988 10742 4016 11086
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3422 9276 3730 9285
rect 3422 9274 3428 9276
rect 3484 9274 3508 9276
rect 3564 9274 3588 9276
rect 3644 9274 3668 9276
rect 3724 9274 3730 9276
rect 3484 9222 3486 9274
rect 3666 9222 3668 9274
rect 3422 9220 3428 9222
rect 3484 9220 3508 9222
rect 3564 9220 3588 9222
rect 3644 9220 3668 9222
rect 3724 9220 3730 9222
rect 3422 9211 3730 9220
rect 3896 8974 3924 9998
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 3422 8188 3730 8197
rect 3422 8186 3428 8188
rect 3484 8186 3508 8188
rect 3564 8186 3588 8188
rect 3644 8186 3668 8188
rect 3724 8186 3730 8188
rect 3484 8134 3486 8186
rect 3666 8134 3668 8186
rect 3422 8132 3428 8134
rect 3484 8132 3508 8134
rect 3564 8132 3588 8134
rect 3644 8132 3668 8134
rect 3724 8132 3730 8134
rect 3422 8123 3730 8132
rect 3896 7886 3924 8910
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3896 7206 3924 7822
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3422 7100 3730 7109
rect 3422 7098 3428 7100
rect 3484 7098 3508 7100
rect 3564 7098 3588 7100
rect 3644 7098 3668 7100
rect 3724 7098 3730 7100
rect 3484 7046 3486 7098
rect 3666 7046 3668 7098
rect 3422 7044 3428 7046
rect 3484 7044 3508 7046
rect 3564 7044 3588 7046
rect 3644 7044 3668 7046
rect 3724 7044 3730 7046
rect 3422 7035 3730 7044
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 4264 6458 4292 12854
rect 4356 12646 4384 12854
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4356 11830 4384 12582
rect 4632 12238 4660 13126
rect 4908 12782 4936 13330
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4908 12306 4936 12582
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4436 12164 4488 12170
rect 4436 12106 4488 12112
rect 4344 11824 4396 11830
rect 4344 11766 4396 11772
rect 4448 11762 4476 12106
rect 4632 11762 4660 12174
rect 5276 12170 5304 14418
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 12986 5580 14214
rect 5644 13938 5672 16050
rect 5736 15094 5764 16186
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 5736 14414 5764 15030
rect 5828 14414 5856 16390
rect 5894 16348 6202 16357
rect 5894 16346 5900 16348
rect 5956 16346 5980 16348
rect 6036 16346 6060 16348
rect 6116 16346 6140 16348
rect 6196 16346 6202 16348
rect 5956 16294 5958 16346
rect 6138 16294 6140 16346
rect 5894 16292 5900 16294
rect 5956 16292 5980 16294
rect 6036 16292 6060 16294
rect 6116 16292 6140 16294
rect 6196 16292 6202 16294
rect 5894 16283 6202 16292
rect 6564 16114 6592 16934
rect 6840 16522 6868 17070
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 6828 16516 6880 16522
rect 6828 16458 6880 16464
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6840 15638 6868 16458
rect 6932 16046 6960 16662
rect 7576 16590 7604 16934
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 5894 15260 6202 15269
rect 5894 15258 5900 15260
rect 5956 15258 5980 15260
rect 6036 15258 6060 15260
rect 6116 15258 6140 15260
rect 6196 15258 6202 15260
rect 5956 15206 5958 15258
rect 6138 15206 6140 15258
rect 5894 15204 5900 15206
rect 5956 15204 5980 15206
rect 6036 15204 6060 15206
rect 6116 15204 6140 15206
rect 6196 15204 6202 15206
rect 5894 15195 6202 15204
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5644 13326 5672 13874
rect 5736 13870 5764 14350
rect 5894 14172 6202 14181
rect 5894 14170 5900 14172
rect 5956 14170 5980 14172
rect 6036 14170 6060 14172
rect 6116 14170 6140 14172
rect 6196 14170 6202 14172
rect 5956 14118 5958 14170
rect 6138 14118 6140 14170
rect 5894 14116 5900 14118
rect 5956 14116 5980 14118
rect 6036 14116 6060 14118
rect 6116 14116 6140 14118
rect 6196 14116 6202 14118
rect 5894 14107 6202 14116
rect 6840 14006 6868 14758
rect 6828 14000 6880 14006
rect 6932 13972 6960 15846
rect 7300 15094 7328 15982
rect 7484 15978 7512 16390
rect 7576 16114 7604 16526
rect 7760 16522 7788 17138
rect 7944 16590 7972 17138
rect 8367 16892 8675 16901
rect 8367 16890 8373 16892
rect 8429 16890 8453 16892
rect 8509 16890 8533 16892
rect 8589 16890 8613 16892
rect 8669 16890 8675 16892
rect 8429 16838 8431 16890
rect 8611 16838 8613 16890
rect 8367 16836 8373 16838
rect 8429 16836 8453 16838
rect 8509 16836 8533 16838
rect 8589 16836 8613 16838
rect 8669 16836 8675 16838
rect 8367 16827 8675 16836
rect 13312 16892 13620 16901
rect 13312 16890 13318 16892
rect 13374 16890 13398 16892
rect 13454 16890 13478 16892
rect 13534 16890 13558 16892
rect 13614 16890 13620 16892
rect 13374 16838 13376 16890
rect 13556 16838 13558 16890
rect 13312 16836 13318 16838
rect 13374 16836 13398 16838
rect 13454 16836 13478 16838
rect 13534 16836 13558 16838
rect 13614 16836 13620 16838
rect 13312 16827 13620 16836
rect 18257 16892 18565 16901
rect 18257 16890 18263 16892
rect 18319 16890 18343 16892
rect 18399 16890 18423 16892
rect 18479 16890 18503 16892
rect 18559 16890 18565 16892
rect 18319 16838 18321 16890
rect 18501 16838 18503 16890
rect 18257 16836 18263 16838
rect 18319 16836 18343 16838
rect 18399 16836 18423 16838
rect 18479 16836 18503 16838
rect 18559 16836 18565 16838
rect 18257 16827 18565 16836
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7288 15088 7340 15094
rect 7288 15030 7340 15036
rect 7300 14890 7328 15030
rect 7104 14884 7156 14890
rect 7104 14826 7156 14832
rect 7288 14884 7340 14890
rect 7288 14826 7340 14832
rect 7116 14074 7144 14826
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7288 14340 7340 14346
rect 7288 14282 7340 14288
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 6828 13942 6880 13948
rect 6920 13966 6972 13972
rect 6920 13908 6972 13914
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5894 13084 6202 13093
rect 5894 13082 5900 13084
rect 5956 13082 5980 13084
rect 6036 13082 6060 13084
rect 6116 13082 6140 13084
rect 6196 13082 6202 13084
rect 5956 13030 5958 13082
rect 6138 13030 6140 13082
rect 5894 13028 5900 13030
rect 5956 13028 5980 13030
rect 6036 13028 6060 13030
rect 6116 13028 6140 13030
rect 6196 13028 6202 13030
rect 5894 13019 6202 13028
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5368 12594 5396 12786
rect 5368 12566 5672 12594
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5460 12306 5488 12378
rect 5644 12306 5672 12566
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5264 12164 5316 12170
rect 5264 12106 5316 12112
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4632 9450 4660 11698
rect 4620 9444 4672 9450
rect 4620 9386 4672 9392
rect 4908 8974 4936 12038
rect 5460 11762 5488 12242
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5736 11642 5764 12786
rect 6656 12374 6684 13806
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6840 12434 6868 13262
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6748 12406 6868 12434
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 5894 11996 6202 12005
rect 5894 11994 5900 11996
rect 5956 11994 5980 11996
rect 6036 11994 6060 11996
rect 6116 11994 6140 11996
rect 6196 11994 6202 11996
rect 5956 11942 5958 11994
rect 6138 11942 6140 11994
rect 5894 11940 5900 11942
rect 5956 11940 5980 11942
rect 6036 11940 6060 11942
rect 6116 11940 6140 11942
rect 6196 11940 6202 11942
rect 5894 11931 6202 11940
rect 5552 11626 5764 11642
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 5540 11620 5764 11626
rect 5592 11614 5764 11620
rect 5540 11562 5592 11568
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 5552 8634 5580 11562
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 3422 6012 3730 6021
rect 3422 6010 3428 6012
rect 3484 6010 3508 6012
rect 3564 6010 3588 6012
rect 3644 6010 3668 6012
rect 3724 6010 3730 6012
rect 3484 5958 3486 6010
rect 3666 5958 3668 6010
rect 3422 5956 3428 5958
rect 3484 5956 3508 5958
rect 3564 5956 3588 5958
rect 3644 5956 3668 5958
rect 3724 5956 3730 5958
rect 3422 5947 3730 5956
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4540 5234 4568 5646
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 2778 5128 2834 5137
rect 2778 5063 2780 5072
rect 2832 5063 2834 5072
rect 2962 5128 3018 5137
rect 2962 5063 3018 5072
rect 2780 5034 2832 5040
rect 3422 4924 3730 4933
rect 3422 4922 3428 4924
rect 3484 4922 3508 4924
rect 3564 4922 3588 4924
rect 3644 4922 3668 4924
rect 3724 4922 3730 4924
rect 3484 4870 3486 4922
rect 3666 4870 3668 4922
rect 3422 4868 3428 4870
rect 3484 4868 3508 4870
rect 3564 4868 3588 4870
rect 3644 4868 3668 4870
rect 3724 4868 3730 4870
rect 3422 4859 3730 4868
rect 4540 4690 4568 5170
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 3422 3836 3730 3845
rect 3422 3834 3428 3836
rect 3484 3834 3508 3836
rect 3564 3834 3588 3836
rect 3644 3834 3668 3836
rect 3724 3834 3730 3836
rect 3484 3782 3486 3834
rect 3666 3782 3668 3834
rect 3422 3780 3428 3782
rect 3484 3780 3508 3782
rect 3564 3780 3588 3782
rect 3644 3780 3668 3782
rect 3724 3780 3730 3782
rect 3422 3771 3730 3780
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3160 3641 3188 3674
rect 3146 3632 3202 3641
rect 3146 3567 3202 3576
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 2332 2582 2360 2926
rect 2976 2650 3004 3402
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3344 3194 3372 3334
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3344 2650 3372 3130
rect 3422 2748 3730 2757
rect 3422 2746 3428 2748
rect 3484 2746 3508 2748
rect 3564 2746 3588 2748
rect 3644 2746 3668 2748
rect 3724 2746 3730 2748
rect 3484 2694 3486 2746
rect 3666 2694 3668 2746
rect 3422 2692 3428 2694
rect 3484 2692 3508 2694
rect 3564 2692 3588 2694
rect 3644 2692 3668 2694
rect 3724 2692 3730 2694
rect 3422 2683 3730 2692
rect 3988 2650 4016 4490
rect 4540 4146 4568 4626
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4540 3126 4568 4082
rect 4816 3398 4844 4422
rect 5552 3738 5580 6666
rect 5828 5574 5856 11630
rect 5894 10908 6202 10917
rect 5894 10906 5900 10908
rect 5956 10906 5980 10908
rect 6036 10906 6060 10908
rect 6116 10906 6140 10908
rect 6196 10906 6202 10908
rect 5956 10854 5958 10906
rect 6138 10854 6140 10906
rect 5894 10852 5900 10854
rect 5956 10852 5980 10854
rect 6036 10852 6060 10854
rect 6116 10852 6140 10854
rect 6196 10852 6202 10854
rect 5894 10843 6202 10852
rect 5894 9820 6202 9829
rect 5894 9818 5900 9820
rect 5956 9818 5980 9820
rect 6036 9818 6060 9820
rect 6116 9818 6140 9820
rect 6196 9818 6202 9820
rect 5956 9766 5958 9818
rect 6138 9766 6140 9818
rect 5894 9764 5900 9766
rect 5956 9764 5980 9766
rect 6036 9764 6060 9766
rect 6116 9764 6140 9766
rect 6196 9764 6202 9766
rect 5894 9755 6202 9764
rect 6748 9382 6776 12406
rect 6932 12102 6960 12786
rect 7024 12646 7052 14010
rect 7300 14006 7328 14282
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7288 14000 7340 14006
rect 7288 13942 7340 13948
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 7116 12238 7144 12922
rect 7208 12850 7236 13874
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7300 12782 7328 13942
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7300 12306 7328 12718
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6932 11762 6960 12038
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6840 10062 6868 10746
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6932 9178 6960 11698
rect 7300 11694 7328 12242
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 7024 10062 7052 10542
rect 7116 10062 7144 11222
rect 7208 11218 7236 11494
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7392 11098 7420 12786
rect 7208 11082 7420 11098
rect 7196 11076 7420 11082
rect 7248 11070 7420 11076
rect 7196 11018 7248 11024
rect 7208 10266 7236 11018
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7024 9518 7052 9998
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7024 9042 7052 9454
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 5894 8732 6202 8741
rect 5894 8730 5900 8732
rect 5956 8730 5980 8732
rect 6036 8730 6060 8732
rect 6116 8730 6140 8732
rect 6196 8730 6202 8732
rect 5956 8678 5958 8730
rect 6138 8678 6140 8730
rect 5894 8676 5900 8678
rect 5956 8676 5980 8678
rect 6036 8676 6060 8678
rect 6116 8676 6140 8678
rect 6196 8676 6202 8678
rect 5894 8667 6202 8676
rect 7024 7954 7052 8978
rect 7484 8242 7512 14214
rect 7576 13530 7604 14418
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7668 11898 7696 15846
rect 7760 15502 7788 16458
rect 10839 16348 11147 16357
rect 10839 16346 10845 16348
rect 10901 16346 10925 16348
rect 10981 16346 11005 16348
rect 11061 16346 11085 16348
rect 11141 16346 11147 16348
rect 10901 16294 10903 16346
rect 11083 16294 11085 16346
rect 10839 16292 10845 16294
rect 10901 16292 10925 16294
rect 10981 16292 11005 16294
rect 11061 16292 11085 16294
rect 11141 16292 11147 16294
rect 10839 16283 11147 16292
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7760 15042 7788 15438
rect 7852 15162 7880 15982
rect 9220 15972 9272 15978
rect 9220 15914 9272 15920
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8367 15804 8675 15813
rect 8367 15802 8373 15804
rect 8429 15802 8453 15804
rect 8509 15802 8533 15804
rect 8589 15802 8613 15804
rect 8669 15802 8675 15804
rect 8429 15750 8431 15802
rect 8611 15750 8613 15802
rect 8367 15748 8373 15750
rect 8429 15748 8453 15750
rect 8509 15748 8533 15750
rect 8589 15748 8613 15750
rect 8669 15748 8675 15750
rect 8367 15739 8675 15748
rect 8024 15428 8076 15434
rect 8024 15370 8076 15376
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7760 15014 7880 15042
rect 7852 13938 7880 15014
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 7944 14482 7972 14962
rect 8036 14958 8064 15370
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 8036 14414 8064 14894
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8220 14618 8248 14758
rect 8367 14716 8675 14725
rect 8367 14714 8373 14716
rect 8429 14714 8453 14716
rect 8509 14714 8533 14716
rect 8589 14714 8613 14716
rect 8669 14714 8675 14716
rect 8429 14662 8431 14714
rect 8611 14662 8613 14714
rect 8367 14660 8373 14662
rect 8429 14660 8453 14662
rect 8509 14660 8533 14662
rect 8589 14660 8613 14662
rect 8669 14660 8675 14662
rect 8367 14651 8675 14660
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 8036 13938 8064 14350
rect 7840 13932 7892 13938
rect 7840 13874 7892 13880
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7564 11620 7616 11626
rect 7564 11562 7616 11568
rect 7576 11218 7604 11562
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7392 8214 7512 8242
rect 7392 8090 7420 8214
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7012 7948 7064 7954
rect 7012 7890 7064 7896
rect 5894 7644 6202 7653
rect 5894 7642 5900 7644
rect 5956 7642 5980 7644
rect 6036 7642 6060 7644
rect 6116 7642 6140 7644
rect 6196 7642 6202 7644
rect 5956 7590 5958 7642
rect 6138 7590 6140 7642
rect 5894 7588 5900 7590
rect 5956 7588 5980 7590
rect 6036 7588 6060 7590
rect 6116 7588 6140 7590
rect 6196 7588 6202 7590
rect 5894 7579 6202 7588
rect 7024 7546 7052 7890
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 5894 6556 6202 6565
rect 5894 6554 5900 6556
rect 5956 6554 5980 6556
rect 6036 6554 6060 6556
rect 6116 6554 6140 6556
rect 6196 6554 6202 6556
rect 5956 6502 5958 6554
rect 6138 6502 6140 6554
rect 5894 6500 5900 6502
rect 5956 6500 5980 6502
rect 6036 6500 6060 6502
rect 6116 6500 6140 6502
rect 6196 6500 6202 6502
rect 5894 6491 6202 6500
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5894 5468 6202 5477
rect 5894 5466 5900 5468
rect 5956 5466 5980 5468
rect 6036 5466 6060 5468
rect 6116 5466 6140 5468
rect 6196 5466 6202 5468
rect 5956 5414 5958 5466
rect 6138 5414 6140 5466
rect 5894 5412 5900 5414
rect 5956 5412 5980 5414
rect 6036 5412 6060 5414
rect 6116 5412 6140 5414
rect 6196 5412 6202 5414
rect 5894 5403 6202 5412
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 4816 3126 4844 3334
rect 5644 3194 5672 5170
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 5828 3058 5856 4966
rect 7116 4690 7144 6190
rect 7576 5370 7604 11154
rect 7852 9926 7880 13874
rect 7932 13796 7984 13802
rect 7932 13738 7984 13744
rect 7944 12238 7972 13738
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7944 8498 7972 12174
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 8036 8090 8064 13874
rect 8367 13628 8675 13637
rect 8367 13626 8373 13628
rect 8429 13626 8453 13628
rect 8509 13626 8533 13628
rect 8589 13626 8613 13628
rect 8669 13626 8675 13628
rect 8429 13574 8431 13626
rect 8611 13574 8613 13626
rect 8367 13572 8373 13574
rect 8429 13572 8453 13574
rect 8509 13572 8533 13574
rect 8589 13572 8613 13574
rect 8669 13572 8675 13574
rect 8367 13563 8675 13572
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 8220 8974 8248 13194
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8367 12540 8675 12549
rect 8367 12538 8373 12540
rect 8429 12538 8453 12540
rect 8509 12538 8533 12540
rect 8589 12538 8613 12540
rect 8669 12538 8675 12540
rect 8429 12486 8431 12538
rect 8611 12486 8613 12538
rect 8367 12484 8373 12486
rect 8429 12484 8453 12486
rect 8509 12484 8533 12486
rect 8589 12484 8613 12486
rect 8669 12484 8675 12486
rect 8367 12475 8675 12484
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8404 11762 8432 12038
rect 8772 11830 8800 12582
rect 8760 11824 8812 11830
rect 8760 11766 8812 11772
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8367 11452 8675 11461
rect 8367 11450 8373 11452
rect 8429 11450 8453 11452
rect 8509 11450 8533 11452
rect 8589 11450 8613 11452
rect 8669 11450 8675 11452
rect 8429 11398 8431 11450
rect 8611 11398 8613 11450
rect 8367 11396 8373 11398
rect 8429 11396 8453 11398
rect 8509 11396 8533 11398
rect 8589 11396 8613 11398
rect 8669 11396 8675 11398
rect 8367 11387 8675 11396
rect 8367 10364 8675 10373
rect 8367 10362 8373 10364
rect 8429 10362 8453 10364
rect 8509 10362 8533 10364
rect 8589 10362 8613 10364
rect 8669 10362 8675 10364
rect 8429 10310 8431 10362
rect 8611 10310 8613 10362
rect 8367 10308 8373 10310
rect 8429 10308 8453 10310
rect 8509 10308 8533 10310
rect 8589 10308 8613 10310
rect 8669 10308 8675 10310
rect 8367 10299 8675 10308
rect 8864 9586 8892 15846
rect 9232 15706 9260 15914
rect 9416 15706 9444 16050
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9232 14414 9260 15642
rect 9692 15162 9720 15982
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9496 14544 9548 14550
rect 9496 14486 9548 14492
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 8944 13796 8996 13802
rect 8944 13738 8996 13744
rect 8956 13394 8984 13738
rect 8944 13388 8996 13394
rect 8944 13330 8996 13336
rect 8956 12782 8984 13330
rect 9048 12850 9076 13874
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8956 12238 8984 12718
rect 9140 12442 9168 13262
rect 9232 12918 9260 13874
rect 9324 13530 9352 14214
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 9232 12782 9260 12854
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 9232 12322 9260 12582
rect 9416 12442 9444 12786
rect 9404 12436 9456 12442
rect 9048 12306 9260 12322
rect 9036 12300 9260 12306
rect 9088 12294 9260 12300
rect 9324 12406 9404 12434
rect 9036 12242 9088 12248
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8367 9276 8675 9285
rect 8367 9274 8373 9276
rect 8429 9274 8453 9276
rect 8509 9274 8533 9276
rect 8589 9274 8613 9276
rect 8669 9274 8675 9276
rect 8429 9222 8431 9274
rect 8611 9222 8613 9274
rect 8367 9220 8373 9222
rect 8429 9220 8453 9222
rect 8509 9220 8533 9222
rect 8589 9220 8613 9222
rect 8669 9220 8675 9222
rect 8367 9211 8675 9220
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8367 8188 8675 8197
rect 8367 8186 8373 8188
rect 8429 8186 8453 8188
rect 8509 8186 8533 8188
rect 8589 8186 8613 8188
rect 8669 8186 8675 8188
rect 8429 8134 8431 8186
rect 8611 8134 8613 8186
rect 8367 8132 8373 8134
rect 8429 8132 8453 8134
rect 8509 8132 8533 8134
rect 8589 8132 8613 8134
rect 8669 8132 8675 8134
rect 8367 8123 8675 8132
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7852 6934 7880 7346
rect 8367 7100 8675 7109
rect 8367 7098 8373 7100
rect 8429 7098 8453 7100
rect 8509 7098 8533 7100
rect 8589 7098 8613 7100
rect 8669 7098 8675 7100
rect 8429 7046 8431 7098
rect 8611 7046 8613 7098
rect 8367 7044 8373 7046
rect 8429 7044 8453 7046
rect 8509 7044 8533 7046
rect 8589 7044 8613 7046
rect 8669 7044 8675 7046
rect 8367 7035 8675 7044
rect 7840 6928 7892 6934
rect 7840 6870 7892 6876
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 5894 4380 6202 4389
rect 5894 4378 5900 4380
rect 5956 4378 5980 4380
rect 6036 4378 6060 4380
rect 6116 4378 6140 4380
rect 6196 4378 6202 4380
rect 5956 4326 5958 4378
rect 6138 4326 6140 4378
rect 5894 4324 5900 4326
rect 5956 4324 5980 4326
rect 6036 4324 6060 4326
rect 6116 4324 6140 4326
rect 6196 4324 6202 4326
rect 5894 4315 6202 4324
rect 6656 4214 6684 4422
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 7116 4146 7144 4626
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 5894 3292 6202 3301
rect 5894 3290 5900 3292
rect 5956 3290 5980 3292
rect 6036 3290 6060 3292
rect 6116 3290 6140 3292
rect 6196 3290 6202 3292
rect 5956 3238 5958 3290
rect 6138 3238 6140 3290
rect 5894 3236 5900 3238
rect 5956 3236 5980 3238
rect 6036 3236 6060 3238
rect 6116 3236 6140 3238
rect 6196 3236 6202 3238
rect 5894 3227 6202 3236
rect 6748 3058 6776 3334
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 5644 2938 5672 2994
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 2320 2576 2372 2582
rect 2320 2518 2372 2524
rect 2332 2446 2360 2518
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 3344 2378 3372 2586
rect 4816 2514 4844 2790
rect 4908 2774 4936 2926
rect 5644 2922 5764 2938
rect 7024 2922 7052 4014
rect 7116 3534 7144 4082
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 5644 2916 5776 2922
rect 5644 2910 5724 2916
rect 5724 2858 5776 2864
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 4908 2746 5028 2774
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 5000 2378 5028 2746
rect 5644 2650 5672 2790
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5736 2378 5764 2858
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 5920 2582 5948 2790
rect 5908 2576 5960 2582
rect 5908 2518 5960 2524
rect 7300 2514 7328 2926
rect 7668 2650 7696 3130
rect 7852 3126 7880 6870
rect 9048 6662 9076 12242
rect 9324 12238 9352 12406
rect 9404 12378 9456 12384
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9140 10538 9168 12174
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 9508 7818 9536 14486
rect 9692 14414 9720 15098
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9678 12200 9734 12209
rect 9784 12170 9812 15302
rect 9876 12238 9904 15574
rect 10428 15434 10456 15846
rect 10888 15706 10916 15846
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 10416 15428 10468 15434
rect 10416 15370 10468 15376
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9678 12135 9680 12144
rect 9732 12135 9734 12144
rect 9772 12164 9824 12170
rect 9680 12106 9732 12112
rect 9772 12106 9824 12112
rect 9784 11898 9812 12106
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9968 11830 9996 14350
rect 10428 13734 10456 15370
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 10428 11744 10456 13670
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10520 12442 10548 12718
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 10520 12170 10548 12378
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10612 11830 10640 14758
rect 10704 14618 10732 15438
rect 11072 15366 11100 15438
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10839 15260 11147 15269
rect 10839 15258 10845 15260
rect 10901 15258 10925 15260
rect 10981 15258 11005 15260
rect 11061 15258 11085 15260
rect 11141 15258 11147 15260
rect 10901 15206 10903 15258
rect 11083 15206 11085 15258
rect 10839 15204 10845 15206
rect 10901 15204 10925 15206
rect 10981 15204 11005 15206
rect 11061 15204 11085 15206
rect 11141 15204 11147 15206
rect 10839 15195 11147 15204
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 11256 14550 11284 16050
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 11244 14544 11296 14550
rect 11244 14486 11296 14492
rect 10784 14408 10836 14414
rect 10704 14368 10784 14396
rect 10704 14074 10732 14368
rect 10784 14350 10836 14356
rect 11348 14346 11376 15914
rect 11532 15502 11560 16526
rect 11704 16516 11756 16522
rect 11704 16458 11756 16464
rect 14648 16516 14700 16522
rect 14648 16458 14700 16464
rect 11716 16250 11744 16458
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11440 15094 11468 15438
rect 11716 15366 11744 16186
rect 14660 16114 14688 16458
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15120 16114 15148 16390
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11428 15088 11480 15094
rect 11428 15030 11480 15036
rect 11520 14544 11572 14550
rect 11520 14486 11572 14492
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11336 14340 11388 14346
rect 11336 14282 11388 14288
rect 10839 14172 11147 14181
rect 10839 14170 10845 14172
rect 10901 14170 10925 14172
rect 10981 14170 11005 14172
rect 11061 14170 11085 14172
rect 11141 14170 11147 14172
rect 10901 14118 10903 14170
rect 11083 14118 11085 14170
rect 10839 14116 10845 14118
rect 10901 14116 10925 14118
rect 10981 14116 11005 14118
rect 11061 14116 11085 14118
rect 11141 14116 11147 14118
rect 10839 14107 11147 14116
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10704 12918 10732 13194
rect 10839 13084 11147 13093
rect 10839 13082 10845 13084
rect 10901 13082 10925 13084
rect 10981 13082 11005 13084
rect 11061 13082 11085 13084
rect 11141 13082 11147 13084
rect 10901 13030 10903 13082
rect 11083 13030 11085 13082
rect 10839 13028 10845 13030
rect 10901 13028 10925 13030
rect 10981 13028 11005 13030
rect 11061 13028 11085 13030
rect 11141 13028 11147 13030
rect 10839 13019 11147 13028
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10704 12442 10732 12854
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10796 12102 10824 12174
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10704 11762 10732 12038
rect 10839 11996 11147 12005
rect 10839 11994 10845 11996
rect 10901 11994 10925 11996
rect 10981 11994 11005 11996
rect 11061 11994 11085 11996
rect 11141 11994 11147 11996
rect 10901 11942 10903 11994
rect 11083 11942 11085 11994
rect 10839 11940 10845 11942
rect 10901 11940 10925 11942
rect 10981 11940 11005 11942
rect 11061 11940 11085 11942
rect 11141 11940 11147 11942
rect 10839 11931 11147 11940
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 10508 11756 10560 11762
rect 10428 11716 10508 11744
rect 10508 11698 10560 11704
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10336 10742 10364 11494
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9784 10062 9812 10542
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9784 8974 9812 9998
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9784 8430 9812 8910
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9784 7954 9812 8366
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9784 7546 9812 7890
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9784 6866 9812 7482
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9784 6390 9812 6802
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 10336 6118 10364 6598
rect 10520 6322 10548 11698
rect 10839 10908 11147 10917
rect 10839 10906 10845 10908
rect 10901 10906 10925 10908
rect 10981 10906 11005 10908
rect 11061 10906 11085 10908
rect 11141 10906 11147 10908
rect 10901 10854 10903 10906
rect 11083 10854 11085 10906
rect 10839 10852 10845 10854
rect 10901 10852 10925 10854
rect 10981 10852 11005 10854
rect 11061 10852 11085 10854
rect 11141 10852 11147 10854
rect 10839 10843 11147 10852
rect 11256 10606 11284 11834
rect 11532 11626 11560 14486
rect 11624 13462 11652 14486
rect 11716 14414 11744 15302
rect 11808 14822 11836 15982
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12544 15502 12572 15642
rect 13096 15638 13124 16050
rect 13176 15972 13228 15978
rect 13176 15914 13228 15920
rect 14188 15972 14240 15978
rect 14188 15914 14240 15920
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 13188 15502 13216 15914
rect 13312 15804 13620 15813
rect 13312 15802 13318 15804
rect 13374 15802 13398 15804
rect 13454 15802 13478 15804
rect 13534 15802 13558 15804
rect 13614 15802 13620 15804
rect 13374 15750 13376 15802
rect 13556 15750 13558 15802
rect 13312 15748 13318 15750
rect 13374 15748 13398 15750
rect 13454 15748 13478 15750
rect 13534 15748 13558 15750
rect 13614 15748 13620 15750
rect 13312 15739 13620 15748
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13188 15314 13216 15438
rect 13004 15286 13216 15314
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11808 14482 11836 14758
rect 11992 14498 12020 14962
rect 12176 14618 12204 14962
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 11796 14476 11848 14482
rect 11796 14418 11848 14424
rect 11900 14470 12020 14498
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11900 13938 11928 14470
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11808 13326 11836 13806
rect 12084 13326 12112 14010
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12360 13394 12388 13806
rect 12912 13530 12940 13874
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11624 11762 11652 12174
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11348 10130 11376 11018
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 10839 9820 11147 9829
rect 10839 9818 10845 9820
rect 10901 9818 10925 9820
rect 10981 9818 11005 9820
rect 11061 9818 11085 9820
rect 11141 9818 11147 9820
rect 10901 9766 10903 9818
rect 11083 9766 11085 9818
rect 10839 9764 10845 9766
rect 10901 9764 10925 9766
rect 10981 9764 11005 9766
rect 11061 9764 11085 9766
rect 11141 9764 11147 9766
rect 10839 9755 11147 9764
rect 11440 9042 11468 9998
rect 11532 9178 11560 11562
rect 11624 10266 11652 11698
rect 11716 11694 11744 12582
rect 11808 12442 11836 13262
rect 12084 12714 12112 13262
rect 12072 12708 12124 12714
rect 12072 12650 12124 12656
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 11992 11898 12020 12174
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12084 11762 12112 12174
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 12268 11558 12296 12174
rect 12360 11898 12388 13330
rect 13004 12782 13032 15286
rect 13372 14958 13400 15574
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13096 14278 13124 14758
rect 13312 14716 13620 14725
rect 13312 14714 13318 14716
rect 13374 14714 13398 14716
rect 13454 14714 13478 14716
rect 13534 14714 13558 14716
rect 13614 14714 13620 14716
rect 13374 14662 13376 14714
rect 13556 14662 13558 14714
rect 13312 14660 13318 14662
rect 13374 14660 13398 14662
rect 13454 14660 13478 14662
rect 13534 14660 13558 14662
rect 13614 14660 13620 14662
rect 13312 14651 13620 14660
rect 13648 14414 13676 15438
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13176 14408 13228 14414
rect 13360 14408 13412 14414
rect 13176 14350 13228 14356
rect 13358 14376 13360 14385
rect 13636 14408 13688 14414
rect 13412 14376 13414 14385
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12348 11620 12400 11626
rect 12348 11562 12400 11568
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12360 11150 12388 11562
rect 12452 11354 12480 12106
rect 13004 11762 13032 12718
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 12360 9178 12388 11086
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 12912 9518 12940 10134
rect 13004 9586 13032 11698
rect 13096 11286 13124 14214
rect 13188 13734 13216 14350
rect 13636 14350 13688 14356
rect 13358 14311 13414 14320
rect 13372 14074 13400 14311
rect 13740 14278 13768 14962
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 13188 12986 13216 13670
rect 13312 13628 13620 13637
rect 13312 13626 13318 13628
rect 13374 13626 13398 13628
rect 13454 13626 13478 13628
rect 13534 13626 13558 13628
rect 13614 13626 13620 13628
rect 13374 13574 13376 13626
rect 13556 13574 13558 13626
rect 13312 13572 13318 13574
rect 13374 13572 13398 13574
rect 13454 13572 13478 13574
rect 13534 13572 13558 13574
rect 13614 13572 13620 13574
rect 13312 13563 13620 13572
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13188 11830 13216 12786
rect 13740 12594 13768 14214
rect 13648 12566 13768 12594
rect 13312 12540 13620 12549
rect 13312 12538 13318 12540
rect 13374 12538 13398 12540
rect 13454 12538 13478 12540
rect 13534 12538 13558 12540
rect 13614 12538 13620 12540
rect 13374 12486 13376 12538
rect 13556 12486 13558 12538
rect 13312 12484 13318 12486
rect 13374 12484 13398 12486
rect 13454 12484 13478 12486
rect 13534 12484 13558 12486
rect 13614 12484 13620 12486
rect 13312 12475 13620 12484
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13280 12238 13308 12378
rect 13450 12336 13506 12345
rect 13450 12271 13506 12280
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 13280 11540 13308 12174
rect 13464 11898 13492 12271
rect 13648 12238 13676 12566
rect 13832 12458 13860 15506
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14108 14414 14136 14758
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 14016 13870 14044 14214
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 13740 12430 13860 12458
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13452 11892 13504 11898
rect 13636 11892 13688 11898
rect 13452 11834 13504 11840
rect 13556 11852 13636 11880
rect 13556 11762 13584 11852
rect 13636 11834 13688 11840
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13188 11512 13308 11540
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 13188 10690 13216 11512
rect 13312 11452 13620 11461
rect 13312 11450 13318 11452
rect 13374 11450 13398 11452
rect 13454 11450 13478 11452
rect 13534 11450 13558 11452
rect 13614 11450 13620 11452
rect 13374 11398 13376 11450
rect 13556 11398 13558 11450
rect 13312 11396 13318 11398
rect 13374 11396 13398 11398
rect 13454 11396 13478 11398
rect 13534 11396 13558 11398
rect 13614 11396 13620 11398
rect 13312 11387 13620 11396
rect 13096 10662 13216 10690
rect 13096 10198 13124 10662
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 13740 10554 13768 12430
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13832 10674 13860 11494
rect 14016 11098 14044 13806
rect 14108 11762 14136 14350
rect 14200 13734 14228 15914
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14292 14618 14320 15098
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14384 12306 14412 16050
rect 14568 15978 14596 16050
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14660 15502 14688 15846
rect 14752 15706 14780 15982
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 14936 15638 14964 16050
rect 14924 15632 14976 15638
rect 14924 15574 14976 15580
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14476 15162 14504 15438
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14568 14414 14596 14962
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14556 14408 14608 14414
rect 14556 14350 14608 14356
rect 14464 14340 14516 14346
rect 14464 14282 14516 14288
rect 14476 13802 14504 14282
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14660 14090 14688 14214
rect 14568 14062 14688 14090
rect 14568 13938 14596 14062
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14464 13796 14516 13802
rect 14464 13738 14516 13744
rect 14476 13530 14504 13738
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14568 12714 14596 13670
rect 14556 12708 14608 12714
rect 14556 12650 14608 12656
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14292 11762 14320 12174
rect 14464 12164 14516 12170
rect 14464 12106 14516 12112
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 14108 11558 14136 11698
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14200 11218 14228 11630
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 13924 11070 14044 11098
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 13188 10130 13216 10542
rect 13740 10526 13860 10554
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13312 10364 13620 10373
rect 13312 10362 13318 10364
rect 13374 10362 13398 10364
rect 13454 10362 13478 10364
rect 13534 10362 13558 10364
rect 13614 10362 13620 10364
rect 13374 10310 13376 10362
rect 13556 10310 13558 10362
rect 13312 10308 13318 10310
rect 13374 10308 13398 10310
rect 13454 10308 13478 10310
rect 13534 10308 13558 10310
rect 13614 10308 13620 10310
rect 13312 10299 13620 10308
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 13096 9722 13124 9998
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13740 9586 13768 10406
rect 13832 10198 13860 10526
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 10839 8732 11147 8741
rect 10839 8730 10845 8732
rect 10901 8730 10925 8732
rect 10981 8730 11005 8732
rect 11061 8730 11085 8732
rect 11141 8730 11147 8732
rect 10901 8678 10903 8730
rect 11083 8678 11085 8730
rect 10839 8676 10845 8678
rect 10901 8676 10925 8678
rect 10981 8676 11005 8678
rect 11061 8676 11085 8678
rect 11141 8676 11147 8678
rect 10839 8667 11147 8676
rect 12912 8566 12940 9454
rect 13312 9276 13620 9285
rect 13312 9274 13318 9276
rect 13374 9274 13398 9276
rect 13454 9274 13478 9276
rect 13534 9274 13558 9276
rect 13614 9274 13620 9276
rect 13374 9222 13376 9274
rect 13556 9222 13558 9274
rect 13312 9220 13318 9222
rect 13374 9220 13398 9222
rect 13454 9220 13478 9222
rect 13534 9220 13558 9222
rect 13614 9220 13620 9222
rect 13312 9211 13620 9220
rect 13740 8974 13768 9522
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 10839 7644 11147 7653
rect 10839 7642 10845 7644
rect 10901 7642 10925 7644
rect 10981 7642 11005 7644
rect 11061 7642 11085 7644
rect 11141 7642 11147 7644
rect 10901 7590 10903 7642
rect 11083 7590 11085 7642
rect 10839 7588 10845 7590
rect 10901 7588 10925 7590
rect 10981 7588 11005 7590
rect 11061 7588 11085 7590
rect 11141 7588 11147 7590
rect 10839 7579 11147 7588
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 10839 6556 11147 6565
rect 10839 6554 10845 6556
rect 10901 6554 10925 6556
rect 10981 6554 11005 6556
rect 11061 6554 11085 6556
rect 11141 6554 11147 6556
rect 10901 6502 10903 6554
rect 11083 6502 11085 6554
rect 10839 6500 10845 6502
rect 10901 6500 10925 6502
rect 10981 6500 11005 6502
rect 11061 6500 11085 6502
rect 11141 6500 11147 6502
rect 10839 6491 11147 6500
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 8367 6012 8675 6021
rect 8367 6010 8373 6012
rect 8429 6010 8453 6012
rect 8509 6010 8533 6012
rect 8589 6010 8613 6012
rect 8669 6010 8675 6012
rect 8429 5958 8431 6010
rect 8611 5958 8613 6010
rect 8367 5956 8373 5958
rect 8429 5956 8453 5958
rect 8509 5956 8533 5958
rect 8589 5956 8613 5958
rect 8669 5956 8675 5958
rect 8367 5947 8675 5956
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9600 5166 9628 5646
rect 10839 5468 11147 5477
rect 10839 5466 10845 5468
rect 10901 5466 10925 5468
rect 10981 5466 11005 5468
rect 11061 5466 11085 5468
rect 11141 5466 11147 5468
rect 10901 5414 10903 5466
rect 11083 5414 11085 5466
rect 10839 5412 10845 5414
rect 10901 5412 10925 5414
rect 10981 5412 11005 5414
rect 11061 5412 11085 5414
rect 11141 5412 11147 5414
rect 10839 5403 11147 5412
rect 11150 5264 11206 5273
rect 11440 5234 11468 6054
rect 11716 5642 11744 7142
rect 12636 5642 12664 7686
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12912 5914 12940 7346
rect 13084 7268 13136 7274
rect 13084 7210 13136 7216
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 13004 6458 13032 6598
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 13096 6254 13124 7210
rect 13188 6798 13216 8298
rect 13312 8188 13620 8197
rect 13312 8186 13318 8188
rect 13374 8186 13398 8188
rect 13454 8186 13478 8188
rect 13534 8186 13558 8188
rect 13614 8186 13620 8188
rect 13374 8134 13376 8186
rect 13556 8134 13558 8186
rect 13312 8132 13318 8134
rect 13374 8132 13398 8134
rect 13454 8132 13478 8134
rect 13534 8132 13558 8134
rect 13614 8132 13620 8134
rect 13312 8123 13620 8132
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13280 7342 13308 7890
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13312 7100 13620 7109
rect 13312 7098 13318 7100
rect 13374 7098 13398 7100
rect 13454 7098 13478 7100
rect 13534 7098 13558 7100
rect 13614 7098 13620 7100
rect 13374 7046 13376 7098
rect 13556 7046 13558 7098
rect 13312 7044 13318 7046
rect 13374 7044 13398 7046
rect 13454 7044 13478 7046
rect 13534 7044 13558 7046
rect 13614 7044 13620 7046
rect 13312 7035 13620 7044
rect 13648 6798 13676 8502
rect 13740 8498 13768 8910
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13832 7886 13860 8230
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13740 6798 13768 7686
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 13648 6186 13676 6734
rect 13740 6322 13768 6734
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13312 6012 13620 6021
rect 13312 6010 13318 6012
rect 13374 6010 13398 6012
rect 13454 6010 13478 6012
rect 13534 6010 13558 6012
rect 13614 6010 13620 6012
rect 13374 5958 13376 6010
rect 13556 5958 13558 6010
rect 13312 5956 13318 5958
rect 13374 5956 13398 5958
rect 13454 5956 13478 5958
rect 13534 5956 13558 5958
rect 13614 5956 13620 5958
rect 13312 5947 13620 5956
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 13740 5846 13768 6258
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 12624 5636 12676 5642
rect 12624 5578 12676 5584
rect 13740 5574 13768 5782
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13924 5234 13952 11070
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 14016 10470 14044 10950
rect 14292 10538 14320 11494
rect 14476 11286 14504 12106
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 14476 11150 14504 11222
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14568 10554 14596 12650
rect 14660 12238 14688 13670
rect 14752 12646 14780 13874
rect 14740 12640 14792 12646
rect 14740 12582 14792 12588
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14280 10532 14332 10538
rect 14568 10526 14688 10554
rect 14280 10474 14332 10480
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 14292 10010 14320 10474
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14568 10130 14596 10406
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14200 9982 14320 10010
rect 14660 9994 14688 10526
rect 14844 10130 14872 14554
rect 14936 13394 14964 15574
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 15028 13734 15056 14962
rect 15212 13802 15240 16118
rect 15292 15632 15344 15638
rect 15292 15574 15344 15580
rect 15304 14278 15332 15574
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15488 14618 15516 15302
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15580 14482 15608 16594
rect 15784 16348 16092 16357
rect 15784 16346 15790 16348
rect 15846 16346 15870 16348
rect 15926 16346 15950 16348
rect 16006 16346 16030 16348
rect 16086 16346 16092 16348
rect 15846 16294 15848 16346
rect 16028 16294 16030 16346
rect 15784 16292 15790 16294
rect 15846 16292 15870 16294
rect 15926 16292 15950 16294
rect 16006 16292 16030 16294
rect 16086 16292 16092 16294
rect 15784 16283 16092 16292
rect 20729 16348 21037 16357
rect 20729 16346 20735 16348
rect 20791 16346 20815 16348
rect 20871 16346 20895 16348
rect 20951 16346 20975 16348
rect 21031 16346 21037 16348
rect 20791 16294 20793 16346
rect 20973 16294 20975 16346
rect 20729 16292 20735 16294
rect 20791 16292 20815 16294
rect 20871 16292 20895 16294
rect 20951 16292 20975 16294
rect 21031 16292 21037 16294
rect 20729 16283 21037 16292
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15304 14113 15332 14214
rect 15290 14104 15346 14113
rect 15290 14039 15346 14048
rect 15292 14000 15344 14006
rect 15396 13988 15424 14214
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15344 13960 15424 13988
rect 15292 13942 15344 13948
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14936 12238 14964 12786
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15304 12442 15332 12582
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 14936 10674 14964 12174
rect 15028 11354 15056 12174
rect 15120 12170 15148 12310
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15212 11778 15240 12038
rect 15120 11762 15240 11778
rect 15304 11762 15332 12378
rect 15108 11756 15240 11762
rect 15160 11750 15240 11756
rect 15292 11756 15344 11762
rect 15108 11698 15160 11704
rect 15292 11698 15344 11704
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14936 10266 14964 10610
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 15304 10266 15332 10474
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 14832 10124 14884 10130
rect 14832 10066 14884 10072
rect 14648 9988 14700 9994
rect 14200 9654 14228 9982
rect 14648 9930 14700 9936
rect 15396 9926 15424 13330
rect 15488 10810 15516 14010
rect 15580 12986 15608 14418
rect 15672 14006 15700 16050
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 15948 15706 15976 15982
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 15784 15260 16092 15269
rect 15784 15258 15790 15260
rect 15846 15258 15870 15260
rect 15926 15258 15950 15260
rect 16006 15258 16030 15260
rect 16086 15258 16092 15260
rect 15846 15206 15848 15258
rect 16028 15206 16030 15258
rect 15784 15204 15790 15206
rect 15846 15204 15870 15206
rect 15926 15204 15950 15206
rect 16006 15204 16030 15206
rect 16086 15204 16092 15206
rect 15784 15195 16092 15204
rect 15784 14172 16092 14181
rect 15784 14170 15790 14172
rect 15846 14170 15870 14172
rect 15926 14170 15950 14172
rect 16006 14170 16030 14172
rect 16086 14170 16092 14172
rect 15846 14118 15848 14170
rect 16028 14118 16030 14170
rect 15784 14116 15790 14118
rect 15846 14116 15870 14118
rect 15926 14116 15950 14118
rect 16006 14116 16030 14118
rect 16086 14116 16092 14118
rect 15784 14107 16092 14116
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15658 13832 15714 13841
rect 15658 13767 15714 13776
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15672 11762 15700 13767
rect 15784 13084 16092 13093
rect 15784 13082 15790 13084
rect 15846 13082 15870 13084
rect 15926 13082 15950 13084
rect 16006 13082 16030 13084
rect 16086 13082 16092 13084
rect 15846 13030 15848 13082
rect 16028 13030 16030 13082
rect 15784 13028 15790 13030
rect 15846 13028 15870 13030
rect 15926 13028 15950 13030
rect 16006 13028 16030 13030
rect 16086 13028 16092 13030
rect 15784 13019 16092 13028
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 16040 12170 16068 12786
rect 16028 12164 16080 12170
rect 16028 12106 16080 12112
rect 15784 11996 16092 12005
rect 15784 11994 15790 11996
rect 15846 11994 15870 11996
rect 15926 11994 15950 11996
rect 16006 11994 16030 11996
rect 16086 11994 16092 11996
rect 15846 11942 15848 11994
rect 16028 11942 16030 11994
rect 15784 11940 15790 11942
rect 15846 11940 15870 11942
rect 15926 11940 15950 11942
rect 16006 11940 16030 11942
rect 16086 11940 16092 11942
rect 15784 11931 16092 11940
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15580 10062 15608 11494
rect 15764 11354 15792 11698
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15784 10908 16092 10917
rect 15784 10906 15790 10908
rect 15846 10906 15870 10908
rect 15926 10906 15950 10908
rect 16006 10906 16030 10908
rect 16086 10906 16092 10908
rect 15846 10854 15848 10906
rect 16028 10854 16030 10906
rect 15784 10852 15790 10854
rect 15846 10852 15870 10854
rect 15926 10852 15950 10854
rect 16006 10852 16030 10854
rect 16086 10852 16092 10854
rect 15784 10843 16092 10852
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 14016 8498 14044 8774
rect 14108 8498 14136 9318
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14292 7818 14320 9862
rect 15396 9654 15424 9862
rect 15784 9820 16092 9829
rect 15784 9818 15790 9820
rect 15846 9818 15870 9820
rect 15926 9818 15950 9820
rect 16006 9818 16030 9820
rect 16086 9818 16092 9820
rect 15846 9766 15848 9818
rect 16028 9766 16030 9818
rect 15784 9764 15790 9766
rect 15846 9764 15870 9766
rect 15926 9764 15950 9766
rect 16006 9764 16030 9766
rect 16086 9764 16092 9766
rect 15784 9755 16092 9764
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 14476 8906 14504 9522
rect 15304 9178 15332 9522
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 14476 8090 14504 8842
rect 15784 8732 16092 8741
rect 15784 8730 15790 8732
rect 15846 8730 15870 8732
rect 15926 8730 15950 8732
rect 16006 8730 16030 8732
rect 16086 8730 16092 8732
rect 15846 8678 15848 8730
rect 16028 8678 16030 8730
rect 15784 8676 15790 8678
rect 15846 8676 15870 8678
rect 15926 8676 15950 8678
rect 16006 8676 16030 8678
rect 16086 8676 16092 8678
rect 15784 8667 16092 8676
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15212 8090 15240 8434
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14292 7002 14320 7346
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14476 6934 14504 8026
rect 15212 7410 15240 8026
rect 16132 8022 16160 15846
rect 17052 15706 17080 15982
rect 18257 15804 18565 15813
rect 18257 15802 18263 15804
rect 18319 15802 18343 15804
rect 18399 15802 18423 15804
rect 18479 15802 18503 15804
rect 18559 15802 18565 15804
rect 18319 15750 18321 15802
rect 18501 15750 18503 15802
rect 18257 15748 18263 15750
rect 18319 15748 18343 15750
rect 18399 15748 18423 15750
rect 18479 15748 18503 15750
rect 18559 15748 18565 15750
rect 18257 15739 18565 15748
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 16672 15564 16724 15570
rect 16592 15524 16672 15552
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16500 15162 16528 15438
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16224 14414 16252 15098
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16304 14544 16356 14550
rect 16304 14486 16356 14492
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16316 13802 16344 14486
rect 16408 14006 16436 14962
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16500 14074 16528 14350
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16304 13796 16356 13802
rect 16304 13738 16356 13744
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16224 11830 16252 12174
rect 16212 11824 16264 11830
rect 16212 11766 16264 11772
rect 16408 11762 16436 13942
rect 16592 12782 16620 15524
rect 16672 15506 16724 15512
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 16948 15428 17000 15434
rect 16948 15370 17000 15376
rect 16672 15088 16724 15094
rect 16672 15030 16724 15036
rect 16684 14414 16712 15030
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16684 12850 16712 14350
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16868 12986 16896 13262
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16684 12730 16712 12786
rect 16592 12345 16620 12718
rect 16684 12702 16804 12730
rect 16776 12434 16804 12702
rect 16684 12406 16804 12434
rect 16578 12336 16634 12345
rect 16578 12271 16580 12280
rect 16632 12271 16634 12280
rect 16580 12242 16632 12248
rect 16592 12211 16620 12242
rect 16684 11898 16712 12406
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16316 10062 16344 11494
rect 16408 11150 16436 11494
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16684 9994 16712 11834
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16868 10674 16896 10950
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16868 9654 16896 10134
rect 16856 9648 16908 9654
rect 16856 9590 16908 9596
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16224 9042 16252 9522
rect 16960 9450 16988 15370
rect 17512 15162 17540 15438
rect 18420 15428 18472 15434
rect 18420 15370 18472 15376
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17868 15088 17920 15094
rect 17868 15030 17920 15036
rect 17132 14884 17184 14890
rect 17132 14826 17184 14832
rect 17144 13802 17172 14826
rect 17880 14822 17908 15030
rect 18432 14890 18460 15370
rect 20729 15260 21037 15269
rect 20729 15258 20735 15260
rect 20791 15258 20815 15260
rect 20871 15258 20895 15260
rect 20951 15258 20975 15260
rect 21031 15258 21037 15260
rect 20791 15206 20793 15258
rect 20973 15206 20975 15258
rect 20729 15204 20735 15206
rect 20791 15204 20815 15206
rect 20871 15204 20895 15206
rect 20951 15204 20975 15206
rect 21031 15204 21037 15206
rect 20729 15195 21037 15204
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 18696 15020 18748 15026
rect 18696 14962 18748 14968
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 18420 14884 18472 14890
rect 18420 14826 18472 14832
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17880 14385 17908 14758
rect 17866 14376 17922 14385
rect 17866 14311 17922 14320
rect 17972 14074 18000 14758
rect 18257 14716 18565 14725
rect 18257 14714 18263 14716
rect 18319 14714 18343 14716
rect 18399 14714 18423 14716
rect 18479 14714 18503 14716
rect 18559 14714 18565 14716
rect 18319 14662 18321 14714
rect 18501 14662 18503 14714
rect 18257 14660 18263 14662
rect 18319 14660 18343 14662
rect 18399 14660 18423 14662
rect 18479 14660 18503 14662
rect 18559 14660 18565 14662
rect 18257 14651 18565 14660
rect 18236 14408 18288 14414
rect 18234 14376 18236 14385
rect 18420 14408 18472 14414
rect 18288 14376 18290 14385
rect 18420 14350 18472 14356
rect 18234 14311 18290 14320
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 17960 14068 18012 14074
rect 17880 14028 17960 14056
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17132 13796 17184 13802
rect 17132 13738 17184 13744
rect 17512 13530 17540 13874
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17040 11824 17092 11830
rect 17040 11766 17092 11772
rect 17052 10674 17080 11766
rect 17236 11218 17264 12786
rect 17788 12442 17816 13262
rect 17880 12782 17908 14028
rect 17960 14010 18012 14016
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 17972 12850 18000 13874
rect 18064 13326 18092 14214
rect 18248 13938 18276 14311
rect 18432 13938 18460 14350
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18156 13394 18184 13670
rect 18257 13628 18565 13637
rect 18257 13626 18263 13628
rect 18319 13626 18343 13628
rect 18399 13626 18423 13628
rect 18479 13626 18503 13628
rect 18559 13626 18565 13628
rect 18319 13574 18321 13626
rect 18501 13574 18503 13626
rect 18257 13572 18263 13574
rect 18319 13572 18343 13574
rect 18399 13572 18423 13574
rect 18479 13572 18503 13574
rect 18559 13572 18565 13574
rect 18257 13563 18565 13572
rect 18144 13388 18196 13394
rect 18144 13330 18196 13336
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 17960 12844 18012 12850
rect 18604 12844 18656 12850
rect 18012 12804 18092 12832
rect 17960 12786 18012 12792
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17500 12368 17552 12374
rect 17500 12310 17552 12316
rect 17512 11762 17540 12310
rect 18064 12238 18092 12804
rect 18604 12786 18656 12792
rect 18257 12540 18565 12549
rect 18257 12538 18263 12540
rect 18319 12538 18343 12540
rect 18399 12538 18423 12540
rect 18479 12538 18503 12540
rect 18559 12538 18565 12540
rect 18319 12486 18321 12538
rect 18501 12486 18503 12538
rect 18257 12484 18263 12486
rect 18319 12484 18343 12486
rect 18399 12484 18423 12486
rect 18479 12484 18503 12486
rect 18559 12484 18565 12486
rect 18257 12475 18565 12484
rect 18616 12238 18644 12786
rect 18708 12714 18736 14962
rect 18880 14340 18932 14346
rect 18880 14282 18932 14288
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18800 13938 18828 14010
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18892 12306 18920 14282
rect 18984 14006 19012 14962
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19628 14074 19656 14554
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19536 12442 19564 12786
rect 19524 12436 19576 12442
rect 19444 12406 19524 12434
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 17592 12232 17644 12238
rect 17868 12232 17920 12238
rect 17592 12174 17644 12180
rect 17788 12192 17868 12220
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17224 11212 17276 11218
rect 17224 11154 17276 11160
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17144 9586 17172 10406
rect 17328 9722 17356 11630
rect 17512 9908 17540 11698
rect 17604 11150 17632 12174
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17788 11014 17816 12192
rect 17868 12174 17920 12180
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 17868 11824 17920 11830
rect 17868 11766 17920 11772
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17880 10062 17908 11766
rect 18892 11694 18920 12242
rect 19248 12232 19300 12238
rect 19444 12209 19472 12406
rect 19524 12378 19576 12384
rect 19628 12374 19656 14010
rect 19800 13932 19852 13938
rect 19800 13874 19852 13880
rect 19708 12640 19760 12646
rect 19708 12582 19760 12588
rect 19616 12368 19668 12374
rect 19616 12310 19668 12316
rect 19248 12174 19300 12180
rect 19430 12200 19486 12209
rect 19260 11898 19288 12174
rect 19430 12135 19486 12144
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19444 11830 19472 12135
rect 19432 11824 19484 11830
rect 19432 11766 19484 11772
rect 19156 11756 19208 11762
rect 19156 11698 19208 11704
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18257 11452 18565 11461
rect 18257 11450 18263 11452
rect 18319 11450 18343 11452
rect 18399 11450 18423 11452
rect 18479 11450 18503 11452
rect 18559 11450 18565 11452
rect 18319 11398 18321 11450
rect 18501 11398 18503 11450
rect 18257 11396 18263 11398
rect 18319 11396 18343 11398
rect 18399 11396 18423 11398
rect 18479 11396 18503 11398
rect 18559 11396 18565 11398
rect 18257 11387 18565 11396
rect 18892 11286 18920 11630
rect 18052 11280 18104 11286
rect 18052 11222 18104 11228
rect 18880 11280 18932 11286
rect 18880 11222 18932 11228
rect 18064 10606 18092 11222
rect 19168 11150 19196 11698
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19260 11218 19288 11562
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19168 10810 19196 11086
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 19260 10674 19288 11154
rect 19444 10826 19472 11766
rect 19720 11762 19748 12582
rect 19812 12442 19840 13874
rect 19996 13802 20024 15098
rect 20729 14172 21037 14181
rect 20729 14170 20735 14172
rect 20791 14170 20815 14172
rect 20871 14170 20895 14172
rect 20951 14170 20975 14172
rect 21031 14170 21037 14172
rect 20791 14118 20793 14170
rect 20973 14118 20975 14170
rect 20729 14116 20735 14118
rect 20791 14116 20815 14118
rect 20871 14116 20895 14118
rect 20951 14116 20975 14118
rect 21031 14116 21037 14118
rect 20729 14107 21037 14116
rect 20076 13864 20128 13870
rect 20076 13806 20128 13812
rect 19984 13796 20036 13802
rect 19984 13738 20036 13744
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19904 12850 19932 13262
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19800 12436 19852 12442
rect 19800 12378 19852 12384
rect 19904 12322 19932 12786
rect 19812 12294 19932 12322
rect 19708 11756 19760 11762
rect 19708 11698 19760 11704
rect 19444 10798 19564 10826
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 18064 10062 18092 10542
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18257 10364 18565 10373
rect 18257 10362 18263 10364
rect 18319 10362 18343 10364
rect 18399 10362 18423 10364
rect 18479 10362 18503 10364
rect 18559 10362 18565 10364
rect 18319 10310 18321 10362
rect 18501 10310 18503 10362
rect 18257 10308 18263 10310
rect 18319 10308 18343 10310
rect 18399 10308 18423 10310
rect 18479 10308 18503 10310
rect 18559 10308 18565 10310
rect 18257 10299 18565 10308
rect 18708 10266 18736 10406
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 17592 9920 17644 9926
rect 17512 9880 17592 9908
rect 17592 9862 17644 9868
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17604 9654 17632 9862
rect 17592 9648 17644 9654
rect 17592 9590 17644 9596
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16592 8634 16620 8910
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16684 8430 16712 9318
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 16960 8566 16988 8910
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16120 8016 16172 8022
rect 16120 7958 16172 7964
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15304 7478 15332 7822
rect 15292 7472 15344 7478
rect 15344 7420 15424 7426
rect 15292 7414 15424 7420
rect 15200 7404 15252 7410
rect 15304 7398 15424 7414
rect 15200 7346 15252 7352
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 14464 6928 14516 6934
rect 14464 6870 14516 6876
rect 14476 6798 14504 6870
rect 14844 6866 14872 7142
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14924 6724 14976 6730
rect 14924 6666 14976 6672
rect 14464 6384 14516 6390
rect 14464 6326 14516 6332
rect 14476 5710 14504 6326
rect 14936 5914 14964 6666
rect 15212 6662 15240 7346
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15304 7002 15332 7278
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 15396 6934 15424 7398
rect 15476 7336 15528 7342
rect 15476 7278 15528 7284
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15488 6322 15516 7278
rect 15580 6798 15608 7822
rect 16868 7750 16896 8434
rect 17052 8090 17080 8910
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 15784 7644 16092 7653
rect 15784 7642 15790 7644
rect 15846 7642 15870 7644
rect 15926 7642 15950 7644
rect 16006 7642 16030 7644
rect 16086 7642 16092 7644
rect 15846 7590 15848 7642
rect 16028 7590 16030 7642
rect 15784 7588 15790 7590
rect 15846 7588 15870 7590
rect 15926 7588 15950 7590
rect 16006 7588 16030 7590
rect 16086 7588 16092 7590
rect 15784 7579 16092 7588
rect 16960 7410 16988 7822
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 15580 6458 15608 6734
rect 15784 6556 16092 6565
rect 15784 6554 15790 6556
rect 15846 6554 15870 6556
rect 15926 6554 15950 6556
rect 16006 6554 16030 6556
rect 16086 6554 16092 6556
rect 15846 6502 15848 6554
rect 16028 6502 16030 6554
rect 15784 6500 15790 6502
rect 15846 6500 15870 6502
rect 15926 6500 15950 6502
rect 16006 6500 16030 6502
rect 16086 6500 16092 6502
rect 15784 6491 16092 6500
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 15016 5840 15068 5846
rect 15016 5782 15068 5788
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 15028 5234 15056 5782
rect 16132 5710 16160 6734
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16684 5778 16712 6054
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 15488 5302 15516 5510
rect 15784 5468 16092 5477
rect 15784 5466 15790 5468
rect 15846 5466 15870 5468
rect 15926 5466 15950 5468
rect 16006 5466 16030 5468
rect 16086 5466 16092 5468
rect 15846 5414 15848 5466
rect 16028 5414 16030 5466
rect 15784 5412 15790 5414
rect 15846 5412 15870 5414
rect 15926 5412 15950 5414
rect 16006 5412 16030 5414
rect 16086 5412 16092 5414
rect 15784 5403 16092 5412
rect 15476 5296 15528 5302
rect 16500 5273 16528 5510
rect 15476 5238 15528 5244
rect 16486 5264 16542 5273
rect 11150 5199 11206 5208
rect 11428 5228 11480 5234
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 8367 4924 8675 4933
rect 8367 4922 8373 4924
rect 8429 4922 8453 4924
rect 8509 4922 8533 4924
rect 8589 4922 8613 4924
rect 8669 4922 8675 4924
rect 8429 4870 8431 4922
rect 8611 4870 8613 4922
rect 8367 4868 8373 4870
rect 8429 4868 8453 4870
rect 8509 4868 8533 4870
rect 8589 4868 8613 4870
rect 8669 4868 8675 4870
rect 8367 4859 8675 4868
rect 9600 4622 9628 5102
rect 11164 5098 11192 5199
rect 11428 5170 11480 5176
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 15384 5228 15436 5234
rect 16486 5199 16542 5208
rect 15384 5170 15436 5176
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9600 4078 9628 4558
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 9876 4282 9904 4490
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8220 3602 8248 3878
rect 8367 3836 8675 3845
rect 8367 3834 8373 3836
rect 8429 3834 8453 3836
rect 8509 3834 8533 3836
rect 8589 3834 8613 3836
rect 8669 3834 8675 3836
rect 8429 3782 8431 3834
rect 8611 3782 8613 3834
rect 8367 3780 8373 3782
rect 8429 3780 8453 3782
rect 8509 3780 8533 3782
rect 8589 3780 8613 3782
rect 8669 3780 8675 3782
rect 8367 3771 8675 3780
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 9600 3534 9628 4014
rect 9692 3738 9720 4082
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 8772 2990 8800 3334
rect 9600 3126 9628 3470
rect 10428 3466 10456 4422
rect 10839 4380 11147 4389
rect 10839 4378 10845 4380
rect 10901 4378 10925 4380
rect 10981 4378 11005 4380
rect 11061 4378 11085 4380
rect 11141 4378 11147 4380
rect 10901 4326 10903 4378
rect 11083 4326 11085 4378
rect 10839 4324 10845 4326
rect 10901 4324 10925 4326
rect 10981 4324 11005 4326
rect 11061 4324 11085 4326
rect 11141 4324 11147 4326
rect 10839 4315 11147 4324
rect 11256 3534 11284 5034
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12636 4826 12664 4966
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12820 4622 12848 5102
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 9784 3194 9812 3402
rect 10839 3292 11147 3301
rect 10839 3290 10845 3292
rect 10901 3290 10925 3292
rect 10981 3290 11005 3292
rect 11061 3290 11085 3292
rect 11141 3290 11147 3292
rect 10901 3238 10903 3290
rect 11083 3238 11085 3290
rect 10839 3236 10845 3238
rect 10901 3236 10925 3238
rect 10981 3236 11005 3238
rect 11061 3236 11085 3238
rect 11141 3236 11147 3238
rect 10839 3227 11147 3236
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8367 2748 8675 2757
rect 8367 2746 8373 2748
rect 8429 2746 8453 2748
rect 8509 2746 8533 2748
rect 8589 2746 8613 2748
rect 8669 2746 8675 2748
rect 8429 2694 8431 2746
rect 8611 2694 8613 2746
rect 8367 2692 8373 2694
rect 8429 2692 8453 2694
rect 8509 2692 8533 2694
rect 8589 2692 8613 2694
rect 8669 2692 8675 2694
rect 8367 2683 8675 2692
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 8772 2378 8800 2926
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 8864 2446 8892 2790
rect 9600 2514 9628 3062
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10244 2650 10272 2994
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 11716 2582 11744 4082
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11808 3534 11836 3878
rect 11888 3664 11940 3670
rect 11888 3606 11940 3612
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11808 3058 11836 3470
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 11900 2446 11928 3606
rect 12820 3602 12848 4558
rect 12912 4214 12940 5170
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 13312 4924 13620 4933
rect 13312 4922 13318 4924
rect 13374 4922 13398 4924
rect 13454 4922 13478 4924
rect 13534 4922 13558 4924
rect 13614 4922 13620 4924
rect 13374 4870 13376 4922
rect 13556 4870 13558 4922
rect 13312 4868 13318 4870
rect 13374 4868 13398 4870
rect 13454 4868 13478 4870
rect 13534 4868 13558 4870
rect 13614 4868 13620 4870
rect 13312 4859 13620 4868
rect 12992 4276 13044 4282
rect 12992 4218 13044 4224
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 13004 3738 13032 4218
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13312 3836 13620 3845
rect 13312 3834 13318 3836
rect 13374 3834 13398 3836
rect 13454 3834 13478 3836
rect 13534 3834 13558 3836
rect 13614 3834 13620 3836
rect 13374 3782 13376 3834
rect 13556 3782 13558 3834
rect 13312 3780 13318 3782
rect 13374 3780 13398 3782
rect 13454 3780 13478 3782
rect 13534 3780 13558 3782
rect 13614 3780 13620 3782
rect 13312 3771 13620 3780
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 13740 3534 13768 4150
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 11992 2990 12020 3470
rect 12084 3126 12112 3470
rect 13372 3194 13400 3470
rect 14188 3460 14240 3466
rect 14188 3402 14240 3408
rect 14200 3194 14228 3402
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 12084 2854 12112 3062
rect 13188 2922 13492 2938
rect 13176 2916 13504 2922
rect 13228 2910 13452 2916
rect 13176 2858 13228 2864
rect 13452 2858 13504 2864
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 13312 2748 13620 2757
rect 13312 2746 13318 2748
rect 13374 2746 13398 2748
rect 13454 2746 13478 2748
rect 13534 2746 13558 2748
rect 13614 2746 13620 2748
rect 13374 2694 13376 2746
rect 13556 2694 13558 2746
rect 13312 2692 13318 2694
rect 13374 2692 13398 2694
rect 13454 2692 13478 2694
rect 13534 2692 13558 2694
rect 13614 2692 13620 2694
rect 13312 2683 13620 2692
rect 13648 2582 13676 3130
rect 14292 3058 14320 5102
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14660 4622 14688 4762
rect 14648 4616 14700 4622
rect 14844 4570 14872 5102
rect 14924 4752 14976 4758
rect 15108 4752 15160 4758
rect 14976 4712 15108 4740
rect 14924 4694 14976 4700
rect 15108 4694 15160 4700
rect 15212 4690 15240 5170
rect 15396 4826 15424 5170
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 14648 4558 14700 4564
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14568 3466 14596 4014
rect 14660 3738 14688 4558
rect 14752 4554 14872 4570
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 14740 4548 14872 4554
rect 14792 4542 14872 4548
rect 14740 4490 14792 4496
rect 14844 4146 14872 4542
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 15016 4140 15068 4146
rect 15016 4082 15068 4088
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14936 3534 14964 3946
rect 15028 3602 15056 4082
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 14924 3528 14976 3534
rect 14844 3488 14924 3516
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 14292 2446 14320 2994
rect 14568 2854 14596 3402
rect 14844 2990 14872 3488
rect 14924 3470 14976 3476
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14936 2650 14964 2994
rect 15028 2990 15056 3538
rect 15396 3398 15424 4558
rect 15784 4380 16092 4389
rect 15784 4378 15790 4380
rect 15846 4378 15870 4380
rect 15926 4378 15950 4380
rect 16006 4378 16030 4380
rect 16086 4378 16092 4380
rect 15846 4326 15848 4378
rect 16028 4326 16030 4378
rect 15784 4324 15790 4326
rect 15846 4324 15870 4326
rect 15926 4324 15950 4326
rect 16006 4324 16030 4326
rect 16086 4324 16092 4326
rect 15784 4315 16092 4324
rect 16500 3942 16528 5199
rect 16684 4622 16712 5714
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 16868 4146 16896 4490
rect 16960 4282 16988 7346
rect 17052 6798 17080 8026
rect 17144 7886 17172 8366
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 6322 17264 6598
rect 17420 6390 17448 6938
rect 17880 6798 17908 9998
rect 17960 9988 18012 9994
rect 17960 9930 18012 9936
rect 17972 9110 18000 9930
rect 18064 9586 18092 9998
rect 18892 9586 18920 10202
rect 19260 10198 19288 10610
rect 19248 10192 19300 10198
rect 19248 10134 19300 10140
rect 19444 9994 19472 10678
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 18064 9178 18092 9522
rect 19536 9450 19564 10798
rect 19812 10742 19840 12294
rect 19892 12232 19944 12238
rect 19892 12174 19944 12180
rect 19904 11558 19932 12174
rect 19996 11898 20024 13738
rect 20088 13258 20116 13806
rect 20076 13252 20128 13258
rect 20076 13194 20128 13200
rect 20729 13084 21037 13093
rect 20729 13082 20735 13084
rect 20791 13082 20815 13084
rect 20871 13082 20895 13084
rect 20951 13082 20975 13084
rect 21031 13082 21037 13084
rect 20791 13030 20793 13082
rect 20973 13030 20975 13082
rect 20729 13028 20735 13030
rect 20791 13028 20815 13030
rect 20871 13028 20895 13030
rect 20951 13028 20975 13030
rect 21031 13028 21037 13030
rect 20729 13019 21037 13028
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19800 10736 19852 10742
rect 19800 10678 19852 10684
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19628 10266 19656 10610
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19524 9444 19576 9450
rect 19524 9386 19576 9392
rect 18257 9276 18565 9285
rect 18257 9274 18263 9276
rect 18319 9274 18343 9276
rect 18399 9274 18423 9276
rect 18479 9274 18503 9276
rect 18559 9274 18565 9276
rect 18319 9222 18321 9274
rect 18501 9222 18503 9274
rect 18257 9220 18263 9222
rect 18319 9220 18343 9222
rect 18399 9220 18423 9222
rect 18479 9220 18503 9222
rect 18559 9220 18565 9222
rect 18257 9211 18565 9220
rect 19904 9178 19932 11494
rect 19996 11082 20024 11834
rect 20180 11218 20208 12378
rect 20729 11996 21037 12005
rect 20729 11994 20735 11996
rect 20791 11994 20815 11996
rect 20871 11994 20895 11996
rect 20951 11994 20975 11996
rect 21031 11994 21037 11996
rect 20791 11942 20793 11994
rect 20973 11942 20975 11994
rect 20729 11940 20735 11942
rect 20791 11940 20815 11942
rect 20871 11940 20895 11942
rect 20951 11940 20975 11942
rect 21031 11940 21037 11942
rect 20729 11931 21037 11940
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 19984 11076 20036 11082
rect 19984 11018 20036 11024
rect 20729 10908 21037 10917
rect 20729 10906 20735 10908
rect 20791 10906 20815 10908
rect 20871 10906 20895 10908
rect 20951 10906 20975 10908
rect 21031 10906 21037 10908
rect 20791 10854 20793 10906
rect 20973 10854 20975 10906
rect 20729 10852 20735 10854
rect 20791 10852 20815 10854
rect 20871 10852 20895 10854
rect 20951 10852 20975 10854
rect 21031 10852 21037 10854
rect 20729 10843 21037 10852
rect 20729 9820 21037 9829
rect 20729 9818 20735 9820
rect 20791 9818 20815 9820
rect 20871 9818 20895 9820
rect 20951 9818 20975 9820
rect 21031 9818 21037 9820
rect 20791 9766 20793 9818
rect 20973 9766 20975 9818
rect 20729 9764 20735 9766
rect 20791 9764 20815 9766
rect 20871 9764 20895 9766
rect 20951 9764 20975 9766
rect 21031 9764 21037 9766
rect 20729 9755 21037 9764
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 19892 9172 19944 9178
rect 19892 9114 19944 9120
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 17972 8634 18000 9046
rect 18064 9042 18092 9114
rect 18052 9036 18104 9042
rect 18052 8978 18104 8984
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 18616 8498 18644 8910
rect 18880 8900 18932 8906
rect 18880 8842 18932 8848
rect 18696 8560 18748 8566
rect 18696 8502 18748 8508
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18257 8188 18565 8197
rect 18257 8186 18263 8188
rect 18319 8186 18343 8188
rect 18399 8186 18423 8188
rect 18479 8186 18503 8188
rect 18559 8186 18565 8188
rect 18319 8134 18321 8186
rect 18501 8134 18503 8186
rect 18257 8132 18263 8134
rect 18319 8132 18343 8134
rect 18399 8132 18423 8134
rect 18479 8132 18503 8134
rect 18559 8132 18565 8134
rect 18257 8123 18565 8132
rect 18616 7970 18644 8298
rect 18708 8022 18736 8502
rect 18892 8362 18920 8842
rect 20729 8732 21037 8741
rect 20729 8730 20735 8732
rect 20791 8730 20815 8732
rect 20871 8730 20895 8732
rect 20951 8730 20975 8732
rect 21031 8730 21037 8732
rect 20791 8678 20793 8730
rect 20973 8678 20975 8730
rect 20729 8676 20735 8678
rect 20791 8676 20815 8678
rect 20871 8676 20895 8678
rect 20951 8676 20975 8678
rect 21031 8676 21037 8678
rect 20729 8667 21037 8676
rect 18880 8356 18932 8362
rect 18880 8298 18932 8304
rect 18892 8022 18920 8298
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 18524 7942 18644 7970
rect 18696 8016 18748 8022
rect 18696 7958 18748 7964
rect 18880 8016 18932 8022
rect 18880 7958 18932 7964
rect 18524 7886 18552 7942
rect 18892 7886 18920 7958
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18524 7546 18552 7822
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18257 7100 18565 7109
rect 18257 7098 18263 7100
rect 18319 7098 18343 7100
rect 18399 7098 18423 7100
rect 18479 7098 18503 7100
rect 18559 7098 18565 7100
rect 18319 7046 18321 7098
rect 18501 7046 18503 7098
rect 18257 7044 18263 7046
rect 18319 7044 18343 7046
rect 18399 7044 18423 7046
rect 18479 7044 18503 7046
rect 18559 7044 18565 7046
rect 18257 7035 18565 7044
rect 18616 6798 18644 7686
rect 18800 6866 18828 7686
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 17408 6384 17460 6390
rect 17408 6326 17460 6332
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 17236 5846 17264 6258
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17512 5370 17540 5646
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 17052 4570 17080 5170
rect 17512 4690 17540 5306
rect 17972 5137 18000 6258
rect 17958 5128 18014 5137
rect 17958 5063 18014 5072
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 18064 4622 18092 6598
rect 18340 6186 18368 6598
rect 18708 6458 18736 6734
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18800 6322 18828 6802
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18328 6180 18380 6186
rect 18328 6122 18380 6128
rect 18257 6012 18565 6021
rect 18257 6010 18263 6012
rect 18319 6010 18343 6012
rect 18399 6010 18423 6012
rect 18479 6010 18503 6012
rect 18559 6010 18565 6012
rect 18319 5958 18321 6010
rect 18501 5958 18503 6010
rect 18257 5956 18263 5958
rect 18319 5956 18343 5958
rect 18399 5956 18423 5958
rect 18479 5956 18503 5958
rect 18559 5956 18565 5958
rect 18257 5947 18565 5956
rect 18892 5642 18920 7822
rect 19628 7750 19656 8230
rect 19616 7744 19668 7750
rect 19616 7686 19668 7692
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18984 5846 19012 6258
rect 18972 5840 19024 5846
rect 18972 5782 19024 5788
rect 19628 5710 19656 7686
rect 20729 7644 21037 7653
rect 20729 7642 20735 7644
rect 20791 7642 20815 7644
rect 20871 7642 20895 7644
rect 20951 7642 20975 7644
rect 21031 7642 21037 7644
rect 20791 7590 20793 7642
rect 20973 7590 20975 7642
rect 20729 7588 20735 7590
rect 20791 7588 20815 7590
rect 20871 7588 20895 7590
rect 20951 7588 20975 7590
rect 21031 7588 21037 7590
rect 20729 7579 21037 7588
rect 20729 6556 21037 6565
rect 20729 6554 20735 6556
rect 20791 6554 20815 6556
rect 20871 6554 20895 6556
rect 20951 6554 20975 6556
rect 21031 6554 21037 6556
rect 20791 6502 20793 6554
rect 20973 6502 20975 6554
rect 20729 6500 20735 6502
rect 20791 6500 20815 6502
rect 20871 6500 20895 6502
rect 20951 6500 20975 6502
rect 21031 6500 21037 6502
rect 20729 6491 21037 6500
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 18880 5636 18932 5642
rect 18880 5578 18932 5584
rect 18257 4924 18565 4933
rect 18257 4922 18263 4924
rect 18319 4922 18343 4924
rect 18399 4922 18423 4924
rect 18479 4922 18503 4924
rect 18559 4922 18565 4924
rect 18319 4870 18321 4922
rect 18501 4870 18503 4922
rect 18257 4868 18263 4870
rect 18319 4868 18343 4870
rect 18399 4868 18423 4870
rect 18479 4868 18503 4870
rect 18559 4868 18565 4870
rect 18257 4859 18565 4868
rect 19628 4758 19656 5646
rect 20729 5468 21037 5477
rect 20729 5466 20735 5468
rect 20791 5466 20815 5468
rect 20871 5466 20895 5468
rect 20951 5466 20975 5468
rect 21031 5466 21037 5468
rect 20791 5414 20793 5466
rect 20973 5414 20975 5466
rect 20729 5412 20735 5414
rect 20791 5412 20815 5414
rect 20871 5412 20895 5414
rect 20951 5412 20975 5414
rect 21031 5412 21037 5414
rect 20729 5403 21037 5412
rect 19616 4752 19668 4758
rect 19616 4694 19668 4700
rect 17224 4616 17276 4622
rect 17052 4542 17172 4570
rect 18052 4616 18104 4622
rect 17224 4558 17276 4564
rect 17972 4564 18052 4570
rect 17972 4558 18104 4564
rect 17144 4486 17172 4542
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 16948 4276 17000 4282
rect 16948 4218 17000 4224
rect 17144 4146 17172 4422
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 15384 3392 15436 3398
rect 15384 3334 15436 3340
rect 15396 3058 15424 3334
rect 15784 3292 16092 3301
rect 15784 3290 15790 3292
rect 15846 3290 15870 3292
rect 15926 3290 15950 3292
rect 16006 3290 16030 3292
rect 16086 3290 16092 3292
rect 15846 3238 15848 3290
rect 16028 3238 16030 3290
rect 15784 3236 15790 3238
rect 15846 3236 15870 3238
rect 15926 3236 15950 3238
rect 16006 3236 16030 3238
rect 16086 3236 16092 3238
rect 15784 3227 16092 3236
rect 16316 3126 16344 3470
rect 16868 3466 16896 4082
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 17052 3534 17080 3878
rect 17236 3738 17264 4558
rect 17972 4542 18092 4558
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17328 3534 17356 4014
rect 17972 3534 18000 4542
rect 20729 4380 21037 4389
rect 20729 4378 20735 4380
rect 20791 4378 20815 4380
rect 20871 4378 20895 4380
rect 20951 4378 20975 4380
rect 21031 4378 21037 4380
rect 20791 4326 20793 4378
rect 20973 4326 20975 4378
rect 20729 4324 20735 4326
rect 20791 4324 20815 4326
rect 20871 4324 20895 4326
rect 20951 4324 20975 4326
rect 21031 4324 21037 4326
rect 20729 4315 21037 4324
rect 18257 3836 18565 3845
rect 18257 3834 18263 3836
rect 18319 3834 18343 3836
rect 18399 3834 18423 3836
rect 18479 3834 18503 3836
rect 18559 3834 18565 3836
rect 18319 3782 18321 3834
rect 18501 3782 18503 3834
rect 18257 3780 18263 3782
rect 18319 3780 18343 3782
rect 18399 3780 18423 3782
rect 18479 3780 18503 3782
rect 18559 3780 18565 3782
rect 18257 3771 18565 3780
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 15304 2446 15332 2994
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 3332 2372 3384 2378
rect 3332 2314 3384 2320
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 8760 2372 8812 2378
rect 8760 2314 8812 2320
rect 14292 2310 14320 2382
rect 15396 2310 15424 2994
rect 16868 2378 16896 3402
rect 17052 3058 17080 3470
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17328 2990 17356 3470
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 17788 2514 17816 3334
rect 18064 2990 18092 3470
rect 20729 3292 21037 3301
rect 20729 3290 20735 3292
rect 20791 3290 20815 3292
rect 20871 3290 20895 3292
rect 20951 3290 20975 3292
rect 21031 3290 21037 3292
rect 20791 3238 20793 3290
rect 20973 3238 20975 3290
rect 20729 3236 20735 3238
rect 20791 3236 20815 3238
rect 20871 3236 20895 3238
rect 20951 3236 20975 3238
rect 21031 3236 21037 3238
rect 20729 3227 21037 3236
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 18257 2748 18565 2757
rect 18257 2746 18263 2748
rect 18319 2746 18343 2748
rect 18399 2746 18423 2748
rect 18479 2746 18503 2748
rect 18559 2746 18565 2748
rect 18319 2694 18321 2746
rect 18501 2694 18503 2746
rect 18257 2692 18263 2694
rect 18319 2692 18343 2694
rect 18399 2692 18423 2694
rect 18479 2692 18503 2694
rect 18559 2692 18565 2694
rect 18257 2683 18565 2692
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 16856 2372 16908 2378
rect 16856 2314 16908 2320
rect 1952 2304 2004 2310
rect 1952 2246 2004 2252
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 5894 2204 6202 2213
rect 5894 2202 5900 2204
rect 5956 2202 5980 2204
rect 6036 2202 6060 2204
rect 6116 2202 6140 2204
rect 6196 2202 6202 2204
rect 5956 2150 5958 2202
rect 6138 2150 6140 2202
rect 5894 2148 5900 2150
rect 5956 2148 5980 2150
rect 6036 2148 6060 2150
rect 6116 2148 6140 2150
rect 6196 2148 6202 2150
rect 5894 2139 6202 2148
rect 10839 2204 11147 2213
rect 10839 2202 10845 2204
rect 10901 2202 10925 2204
rect 10981 2202 11005 2204
rect 11061 2202 11085 2204
rect 11141 2202 11147 2204
rect 10901 2150 10903 2202
rect 11083 2150 11085 2202
rect 10839 2148 10845 2150
rect 10901 2148 10925 2150
rect 10981 2148 11005 2150
rect 11061 2148 11085 2150
rect 11141 2148 11147 2150
rect 10839 2139 11147 2148
rect 15784 2204 16092 2213
rect 15784 2202 15790 2204
rect 15846 2202 15870 2204
rect 15926 2202 15950 2204
rect 16006 2202 16030 2204
rect 16086 2202 16092 2204
rect 15846 2150 15848 2202
rect 16028 2150 16030 2202
rect 15784 2148 15790 2150
rect 15846 2148 15870 2150
rect 15926 2148 15950 2150
rect 16006 2148 16030 2150
rect 16086 2148 16092 2150
rect 15784 2139 16092 2148
rect 20729 2204 21037 2213
rect 20729 2202 20735 2204
rect 20791 2202 20815 2204
rect 20871 2202 20895 2204
rect 20951 2202 20975 2204
rect 21031 2202 21037 2204
rect 20791 2150 20793 2202
rect 20973 2150 20975 2202
rect 20729 2148 20735 2150
rect 20791 2148 20815 2150
rect 20871 2148 20895 2150
rect 20951 2148 20975 2150
rect 21031 2148 21037 2150
rect 20729 2139 21037 2148
<< via2 >>
rect 5900 19610 5956 19612
rect 5980 19610 6036 19612
rect 6060 19610 6116 19612
rect 6140 19610 6196 19612
rect 5900 19558 5946 19610
rect 5946 19558 5956 19610
rect 5980 19558 6010 19610
rect 6010 19558 6022 19610
rect 6022 19558 6036 19610
rect 6060 19558 6074 19610
rect 6074 19558 6086 19610
rect 6086 19558 6116 19610
rect 6140 19558 6150 19610
rect 6150 19558 6196 19610
rect 5900 19556 5956 19558
rect 5980 19556 6036 19558
rect 6060 19556 6116 19558
rect 6140 19556 6196 19558
rect 10845 19610 10901 19612
rect 10925 19610 10981 19612
rect 11005 19610 11061 19612
rect 11085 19610 11141 19612
rect 10845 19558 10891 19610
rect 10891 19558 10901 19610
rect 10925 19558 10955 19610
rect 10955 19558 10967 19610
rect 10967 19558 10981 19610
rect 11005 19558 11019 19610
rect 11019 19558 11031 19610
rect 11031 19558 11061 19610
rect 11085 19558 11095 19610
rect 11095 19558 11141 19610
rect 10845 19556 10901 19558
rect 10925 19556 10981 19558
rect 11005 19556 11061 19558
rect 11085 19556 11141 19558
rect 15790 19610 15846 19612
rect 15870 19610 15926 19612
rect 15950 19610 16006 19612
rect 16030 19610 16086 19612
rect 15790 19558 15836 19610
rect 15836 19558 15846 19610
rect 15870 19558 15900 19610
rect 15900 19558 15912 19610
rect 15912 19558 15926 19610
rect 15950 19558 15964 19610
rect 15964 19558 15976 19610
rect 15976 19558 16006 19610
rect 16030 19558 16040 19610
rect 16040 19558 16086 19610
rect 15790 19556 15846 19558
rect 15870 19556 15926 19558
rect 15950 19556 16006 19558
rect 16030 19556 16086 19558
rect 20735 19610 20791 19612
rect 20815 19610 20871 19612
rect 20895 19610 20951 19612
rect 20975 19610 21031 19612
rect 20735 19558 20781 19610
rect 20781 19558 20791 19610
rect 20815 19558 20845 19610
rect 20845 19558 20857 19610
rect 20857 19558 20871 19610
rect 20895 19558 20909 19610
rect 20909 19558 20921 19610
rect 20921 19558 20951 19610
rect 20975 19558 20985 19610
rect 20985 19558 21031 19610
rect 20735 19556 20791 19558
rect 20815 19556 20871 19558
rect 20895 19556 20951 19558
rect 20975 19556 21031 19558
rect 3428 19066 3484 19068
rect 3508 19066 3564 19068
rect 3588 19066 3644 19068
rect 3668 19066 3724 19068
rect 3428 19014 3474 19066
rect 3474 19014 3484 19066
rect 3508 19014 3538 19066
rect 3538 19014 3550 19066
rect 3550 19014 3564 19066
rect 3588 19014 3602 19066
rect 3602 19014 3614 19066
rect 3614 19014 3644 19066
rect 3668 19014 3678 19066
rect 3678 19014 3724 19066
rect 3428 19012 3484 19014
rect 3508 19012 3564 19014
rect 3588 19012 3644 19014
rect 3668 19012 3724 19014
rect 8373 19066 8429 19068
rect 8453 19066 8509 19068
rect 8533 19066 8589 19068
rect 8613 19066 8669 19068
rect 8373 19014 8419 19066
rect 8419 19014 8429 19066
rect 8453 19014 8483 19066
rect 8483 19014 8495 19066
rect 8495 19014 8509 19066
rect 8533 19014 8547 19066
rect 8547 19014 8559 19066
rect 8559 19014 8589 19066
rect 8613 19014 8623 19066
rect 8623 19014 8669 19066
rect 8373 19012 8429 19014
rect 8453 19012 8509 19014
rect 8533 19012 8589 19014
rect 8613 19012 8669 19014
rect 13318 19066 13374 19068
rect 13398 19066 13454 19068
rect 13478 19066 13534 19068
rect 13558 19066 13614 19068
rect 13318 19014 13364 19066
rect 13364 19014 13374 19066
rect 13398 19014 13428 19066
rect 13428 19014 13440 19066
rect 13440 19014 13454 19066
rect 13478 19014 13492 19066
rect 13492 19014 13504 19066
rect 13504 19014 13534 19066
rect 13558 19014 13568 19066
rect 13568 19014 13614 19066
rect 13318 19012 13374 19014
rect 13398 19012 13454 19014
rect 13478 19012 13534 19014
rect 13558 19012 13614 19014
rect 18263 19066 18319 19068
rect 18343 19066 18399 19068
rect 18423 19066 18479 19068
rect 18503 19066 18559 19068
rect 18263 19014 18309 19066
rect 18309 19014 18319 19066
rect 18343 19014 18373 19066
rect 18373 19014 18385 19066
rect 18385 19014 18399 19066
rect 18423 19014 18437 19066
rect 18437 19014 18449 19066
rect 18449 19014 18479 19066
rect 18503 19014 18513 19066
rect 18513 19014 18559 19066
rect 18263 19012 18319 19014
rect 18343 19012 18399 19014
rect 18423 19012 18479 19014
rect 18503 19012 18559 19014
rect 1858 18264 1914 18320
rect 1674 10920 1730 10976
rect 5900 18522 5956 18524
rect 5980 18522 6036 18524
rect 6060 18522 6116 18524
rect 6140 18522 6196 18524
rect 5900 18470 5946 18522
rect 5946 18470 5956 18522
rect 5980 18470 6010 18522
rect 6010 18470 6022 18522
rect 6022 18470 6036 18522
rect 6060 18470 6074 18522
rect 6074 18470 6086 18522
rect 6086 18470 6116 18522
rect 6140 18470 6150 18522
rect 6150 18470 6196 18522
rect 5900 18468 5956 18470
rect 5980 18468 6036 18470
rect 6060 18468 6116 18470
rect 6140 18468 6196 18470
rect 10845 18522 10901 18524
rect 10925 18522 10981 18524
rect 11005 18522 11061 18524
rect 11085 18522 11141 18524
rect 10845 18470 10891 18522
rect 10891 18470 10901 18522
rect 10925 18470 10955 18522
rect 10955 18470 10967 18522
rect 10967 18470 10981 18522
rect 11005 18470 11019 18522
rect 11019 18470 11031 18522
rect 11031 18470 11061 18522
rect 11085 18470 11095 18522
rect 11095 18470 11141 18522
rect 10845 18468 10901 18470
rect 10925 18468 10981 18470
rect 11005 18468 11061 18470
rect 11085 18468 11141 18470
rect 15790 18522 15846 18524
rect 15870 18522 15926 18524
rect 15950 18522 16006 18524
rect 16030 18522 16086 18524
rect 15790 18470 15836 18522
rect 15836 18470 15846 18522
rect 15870 18470 15900 18522
rect 15900 18470 15912 18522
rect 15912 18470 15926 18522
rect 15950 18470 15964 18522
rect 15964 18470 15976 18522
rect 15976 18470 16006 18522
rect 16030 18470 16040 18522
rect 16040 18470 16086 18522
rect 15790 18468 15846 18470
rect 15870 18468 15926 18470
rect 15950 18468 16006 18470
rect 16030 18468 16086 18470
rect 20735 18522 20791 18524
rect 20815 18522 20871 18524
rect 20895 18522 20951 18524
rect 20975 18522 21031 18524
rect 20735 18470 20781 18522
rect 20781 18470 20791 18522
rect 20815 18470 20845 18522
rect 20845 18470 20857 18522
rect 20857 18470 20871 18522
rect 20895 18470 20909 18522
rect 20909 18470 20921 18522
rect 20921 18470 20951 18522
rect 20975 18470 20985 18522
rect 20985 18470 21031 18522
rect 20735 18468 20791 18470
rect 20815 18468 20871 18470
rect 20895 18468 20951 18470
rect 20975 18468 21031 18470
rect 3428 17978 3484 17980
rect 3508 17978 3564 17980
rect 3588 17978 3644 17980
rect 3668 17978 3724 17980
rect 3428 17926 3474 17978
rect 3474 17926 3484 17978
rect 3508 17926 3538 17978
rect 3538 17926 3550 17978
rect 3550 17926 3564 17978
rect 3588 17926 3602 17978
rect 3602 17926 3614 17978
rect 3614 17926 3644 17978
rect 3668 17926 3678 17978
rect 3678 17926 3724 17978
rect 3428 17924 3484 17926
rect 3508 17924 3564 17926
rect 3588 17924 3644 17926
rect 3668 17924 3724 17926
rect 8373 17978 8429 17980
rect 8453 17978 8509 17980
rect 8533 17978 8589 17980
rect 8613 17978 8669 17980
rect 8373 17926 8419 17978
rect 8419 17926 8429 17978
rect 8453 17926 8483 17978
rect 8483 17926 8495 17978
rect 8495 17926 8509 17978
rect 8533 17926 8547 17978
rect 8547 17926 8559 17978
rect 8559 17926 8589 17978
rect 8613 17926 8623 17978
rect 8623 17926 8669 17978
rect 8373 17924 8429 17926
rect 8453 17924 8509 17926
rect 8533 17924 8589 17926
rect 8613 17924 8669 17926
rect 13318 17978 13374 17980
rect 13398 17978 13454 17980
rect 13478 17978 13534 17980
rect 13558 17978 13614 17980
rect 13318 17926 13364 17978
rect 13364 17926 13374 17978
rect 13398 17926 13428 17978
rect 13428 17926 13440 17978
rect 13440 17926 13454 17978
rect 13478 17926 13492 17978
rect 13492 17926 13504 17978
rect 13504 17926 13534 17978
rect 13558 17926 13568 17978
rect 13568 17926 13614 17978
rect 13318 17924 13374 17926
rect 13398 17924 13454 17926
rect 13478 17924 13534 17926
rect 13558 17924 13614 17926
rect 18263 17978 18319 17980
rect 18343 17978 18399 17980
rect 18423 17978 18479 17980
rect 18503 17978 18559 17980
rect 18263 17926 18309 17978
rect 18309 17926 18319 17978
rect 18343 17926 18373 17978
rect 18373 17926 18385 17978
rect 18385 17926 18399 17978
rect 18423 17926 18437 17978
rect 18437 17926 18449 17978
rect 18449 17926 18479 17978
rect 18503 17926 18513 17978
rect 18513 17926 18559 17978
rect 18263 17924 18319 17926
rect 18343 17924 18399 17926
rect 18423 17924 18479 17926
rect 18503 17924 18559 17926
rect 5900 17434 5956 17436
rect 5980 17434 6036 17436
rect 6060 17434 6116 17436
rect 6140 17434 6196 17436
rect 5900 17382 5946 17434
rect 5946 17382 5956 17434
rect 5980 17382 6010 17434
rect 6010 17382 6022 17434
rect 6022 17382 6036 17434
rect 6060 17382 6074 17434
rect 6074 17382 6086 17434
rect 6086 17382 6116 17434
rect 6140 17382 6150 17434
rect 6150 17382 6196 17434
rect 5900 17380 5956 17382
rect 5980 17380 6036 17382
rect 6060 17380 6116 17382
rect 6140 17380 6196 17382
rect 10845 17434 10901 17436
rect 10925 17434 10981 17436
rect 11005 17434 11061 17436
rect 11085 17434 11141 17436
rect 10845 17382 10891 17434
rect 10891 17382 10901 17434
rect 10925 17382 10955 17434
rect 10955 17382 10967 17434
rect 10967 17382 10981 17434
rect 11005 17382 11019 17434
rect 11019 17382 11031 17434
rect 11031 17382 11061 17434
rect 11085 17382 11095 17434
rect 11095 17382 11141 17434
rect 10845 17380 10901 17382
rect 10925 17380 10981 17382
rect 11005 17380 11061 17382
rect 11085 17380 11141 17382
rect 15790 17434 15846 17436
rect 15870 17434 15926 17436
rect 15950 17434 16006 17436
rect 16030 17434 16086 17436
rect 15790 17382 15836 17434
rect 15836 17382 15846 17434
rect 15870 17382 15900 17434
rect 15900 17382 15912 17434
rect 15912 17382 15926 17434
rect 15950 17382 15964 17434
rect 15964 17382 15976 17434
rect 15976 17382 16006 17434
rect 16030 17382 16040 17434
rect 16040 17382 16086 17434
rect 15790 17380 15846 17382
rect 15870 17380 15926 17382
rect 15950 17380 16006 17382
rect 16030 17380 16086 17382
rect 20735 17434 20791 17436
rect 20815 17434 20871 17436
rect 20895 17434 20951 17436
rect 20975 17434 21031 17436
rect 20735 17382 20781 17434
rect 20781 17382 20791 17434
rect 20815 17382 20845 17434
rect 20845 17382 20857 17434
rect 20857 17382 20871 17434
rect 20895 17382 20909 17434
rect 20909 17382 20921 17434
rect 20921 17382 20951 17434
rect 20975 17382 20985 17434
rect 20985 17382 21031 17434
rect 20735 17380 20791 17382
rect 20815 17380 20871 17382
rect 20895 17380 20951 17382
rect 20975 17380 21031 17382
rect 3428 16890 3484 16892
rect 3508 16890 3564 16892
rect 3588 16890 3644 16892
rect 3668 16890 3724 16892
rect 3428 16838 3474 16890
rect 3474 16838 3484 16890
rect 3508 16838 3538 16890
rect 3538 16838 3550 16890
rect 3550 16838 3564 16890
rect 3588 16838 3602 16890
rect 3602 16838 3614 16890
rect 3614 16838 3644 16890
rect 3668 16838 3678 16890
rect 3678 16838 3724 16890
rect 3428 16836 3484 16838
rect 3508 16836 3564 16838
rect 3588 16836 3644 16838
rect 3668 16836 3724 16838
rect 3428 15802 3484 15804
rect 3508 15802 3564 15804
rect 3588 15802 3644 15804
rect 3668 15802 3724 15804
rect 3428 15750 3474 15802
rect 3474 15750 3484 15802
rect 3508 15750 3538 15802
rect 3538 15750 3550 15802
rect 3550 15750 3564 15802
rect 3588 15750 3602 15802
rect 3602 15750 3614 15802
rect 3614 15750 3644 15802
rect 3668 15750 3678 15802
rect 3678 15750 3724 15802
rect 3428 15748 3484 15750
rect 3508 15748 3564 15750
rect 3588 15748 3644 15750
rect 3668 15748 3724 15750
rect 3428 14714 3484 14716
rect 3508 14714 3564 14716
rect 3588 14714 3644 14716
rect 3668 14714 3724 14716
rect 3428 14662 3474 14714
rect 3474 14662 3484 14714
rect 3508 14662 3538 14714
rect 3538 14662 3550 14714
rect 3550 14662 3564 14714
rect 3588 14662 3602 14714
rect 3602 14662 3614 14714
rect 3614 14662 3644 14714
rect 3668 14662 3678 14714
rect 3678 14662 3724 14714
rect 3428 14660 3484 14662
rect 3508 14660 3564 14662
rect 3588 14660 3644 14662
rect 3668 14660 3724 14662
rect 3428 13626 3484 13628
rect 3508 13626 3564 13628
rect 3588 13626 3644 13628
rect 3668 13626 3724 13628
rect 3428 13574 3474 13626
rect 3474 13574 3484 13626
rect 3508 13574 3538 13626
rect 3538 13574 3550 13626
rect 3550 13574 3564 13626
rect 3588 13574 3602 13626
rect 3602 13574 3614 13626
rect 3614 13574 3644 13626
rect 3668 13574 3678 13626
rect 3678 13574 3724 13626
rect 3428 13572 3484 13574
rect 3508 13572 3564 13574
rect 3588 13572 3644 13574
rect 3668 13572 3724 13574
rect 3428 12538 3484 12540
rect 3508 12538 3564 12540
rect 3588 12538 3644 12540
rect 3668 12538 3724 12540
rect 3428 12486 3474 12538
rect 3474 12486 3484 12538
rect 3508 12486 3538 12538
rect 3538 12486 3550 12538
rect 3550 12486 3564 12538
rect 3588 12486 3602 12538
rect 3602 12486 3614 12538
rect 3614 12486 3644 12538
rect 3668 12486 3678 12538
rect 3678 12486 3724 12538
rect 3428 12484 3484 12486
rect 3508 12484 3564 12486
rect 3588 12484 3644 12486
rect 3668 12484 3724 12486
rect 3428 11450 3484 11452
rect 3508 11450 3564 11452
rect 3588 11450 3644 11452
rect 3668 11450 3724 11452
rect 3428 11398 3474 11450
rect 3474 11398 3484 11450
rect 3508 11398 3538 11450
rect 3538 11398 3550 11450
rect 3550 11398 3564 11450
rect 3588 11398 3602 11450
rect 3602 11398 3614 11450
rect 3614 11398 3644 11450
rect 3668 11398 3678 11450
rect 3678 11398 3724 11450
rect 3428 11396 3484 11398
rect 3508 11396 3564 11398
rect 3588 11396 3644 11398
rect 3668 11396 3724 11398
rect 3428 10362 3484 10364
rect 3508 10362 3564 10364
rect 3588 10362 3644 10364
rect 3668 10362 3724 10364
rect 3428 10310 3474 10362
rect 3474 10310 3484 10362
rect 3508 10310 3538 10362
rect 3538 10310 3550 10362
rect 3550 10310 3564 10362
rect 3588 10310 3602 10362
rect 3602 10310 3614 10362
rect 3614 10310 3644 10362
rect 3668 10310 3678 10362
rect 3678 10310 3724 10362
rect 3428 10308 3484 10310
rect 3508 10308 3564 10310
rect 3588 10308 3644 10310
rect 3668 10308 3724 10310
rect 3428 9274 3484 9276
rect 3508 9274 3564 9276
rect 3588 9274 3644 9276
rect 3668 9274 3724 9276
rect 3428 9222 3474 9274
rect 3474 9222 3484 9274
rect 3508 9222 3538 9274
rect 3538 9222 3550 9274
rect 3550 9222 3564 9274
rect 3588 9222 3602 9274
rect 3602 9222 3614 9274
rect 3614 9222 3644 9274
rect 3668 9222 3678 9274
rect 3678 9222 3724 9274
rect 3428 9220 3484 9222
rect 3508 9220 3564 9222
rect 3588 9220 3644 9222
rect 3668 9220 3724 9222
rect 3428 8186 3484 8188
rect 3508 8186 3564 8188
rect 3588 8186 3644 8188
rect 3668 8186 3724 8188
rect 3428 8134 3474 8186
rect 3474 8134 3484 8186
rect 3508 8134 3538 8186
rect 3538 8134 3550 8186
rect 3550 8134 3564 8186
rect 3588 8134 3602 8186
rect 3602 8134 3614 8186
rect 3614 8134 3644 8186
rect 3668 8134 3678 8186
rect 3678 8134 3724 8186
rect 3428 8132 3484 8134
rect 3508 8132 3564 8134
rect 3588 8132 3644 8134
rect 3668 8132 3724 8134
rect 3428 7098 3484 7100
rect 3508 7098 3564 7100
rect 3588 7098 3644 7100
rect 3668 7098 3724 7100
rect 3428 7046 3474 7098
rect 3474 7046 3484 7098
rect 3508 7046 3538 7098
rect 3538 7046 3550 7098
rect 3550 7046 3564 7098
rect 3588 7046 3602 7098
rect 3602 7046 3614 7098
rect 3614 7046 3644 7098
rect 3668 7046 3678 7098
rect 3678 7046 3724 7098
rect 3428 7044 3484 7046
rect 3508 7044 3564 7046
rect 3588 7044 3644 7046
rect 3668 7044 3724 7046
rect 5900 16346 5956 16348
rect 5980 16346 6036 16348
rect 6060 16346 6116 16348
rect 6140 16346 6196 16348
rect 5900 16294 5946 16346
rect 5946 16294 5956 16346
rect 5980 16294 6010 16346
rect 6010 16294 6022 16346
rect 6022 16294 6036 16346
rect 6060 16294 6074 16346
rect 6074 16294 6086 16346
rect 6086 16294 6116 16346
rect 6140 16294 6150 16346
rect 6150 16294 6196 16346
rect 5900 16292 5956 16294
rect 5980 16292 6036 16294
rect 6060 16292 6116 16294
rect 6140 16292 6196 16294
rect 5900 15258 5956 15260
rect 5980 15258 6036 15260
rect 6060 15258 6116 15260
rect 6140 15258 6196 15260
rect 5900 15206 5946 15258
rect 5946 15206 5956 15258
rect 5980 15206 6010 15258
rect 6010 15206 6022 15258
rect 6022 15206 6036 15258
rect 6060 15206 6074 15258
rect 6074 15206 6086 15258
rect 6086 15206 6116 15258
rect 6140 15206 6150 15258
rect 6150 15206 6196 15258
rect 5900 15204 5956 15206
rect 5980 15204 6036 15206
rect 6060 15204 6116 15206
rect 6140 15204 6196 15206
rect 5900 14170 5956 14172
rect 5980 14170 6036 14172
rect 6060 14170 6116 14172
rect 6140 14170 6196 14172
rect 5900 14118 5946 14170
rect 5946 14118 5956 14170
rect 5980 14118 6010 14170
rect 6010 14118 6022 14170
rect 6022 14118 6036 14170
rect 6060 14118 6074 14170
rect 6074 14118 6086 14170
rect 6086 14118 6116 14170
rect 6140 14118 6150 14170
rect 6150 14118 6196 14170
rect 5900 14116 5956 14118
rect 5980 14116 6036 14118
rect 6060 14116 6116 14118
rect 6140 14116 6196 14118
rect 8373 16890 8429 16892
rect 8453 16890 8509 16892
rect 8533 16890 8589 16892
rect 8613 16890 8669 16892
rect 8373 16838 8419 16890
rect 8419 16838 8429 16890
rect 8453 16838 8483 16890
rect 8483 16838 8495 16890
rect 8495 16838 8509 16890
rect 8533 16838 8547 16890
rect 8547 16838 8559 16890
rect 8559 16838 8589 16890
rect 8613 16838 8623 16890
rect 8623 16838 8669 16890
rect 8373 16836 8429 16838
rect 8453 16836 8509 16838
rect 8533 16836 8589 16838
rect 8613 16836 8669 16838
rect 13318 16890 13374 16892
rect 13398 16890 13454 16892
rect 13478 16890 13534 16892
rect 13558 16890 13614 16892
rect 13318 16838 13364 16890
rect 13364 16838 13374 16890
rect 13398 16838 13428 16890
rect 13428 16838 13440 16890
rect 13440 16838 13454 16890
rect 13478 16838 13492 16890
rect 13492 16838 13504 16890
rect 13504 16838 13534 16890
rect 13558 16838 13568 16890
rect 13568 16838 13614 16890
rect 13318 16836 13374 16838
rect 13398 16836 13454 16838
rect 13478 16836 13534 16838
rect 13558 16836 13614 16838
rect 18263 16890 18319 16892
rect 18343 16890 18399 16892
rect 18423 16890 18479 16892
rect 18503 16890 18559 16892
rect 18263 16838 18309 16890
rect 18309 16838 18319 16890
rect 18343 16838 18373 16890
rect 18373 16838 18385 16890
rect 18385 16838 18399 16890
rect 18423 16838 18437 16890
rect 18437 16838 18449 16890
rect 18449 16838 18479 16890
rect 18503 16838 18513 16890
rect 18513 16838 18559 16890
rect 18263 16836 18319 16838
rect 18343 16836 18399 16838
rect 18423 16836 18479 16838
rect 18503 16836 18559 16838
rect 5900 13082 5956 13084
rect 5980 13082 6036 13084
rect 6060 13082 6116 13084
rect 6140 13082 6196 13084
rect 5900 13030 5946 13082
rect 5946 13030 5956 13082
rect 5980 13030 6010 13082
rect 6010 13030 6022 13082
rect 6022 13030 6036 13082
rect 6060 13030 6074 13082
rect 6074 13030 6086 13082
rect 6086 13030 6116 13082
rect 6140 13030 6150 13082
rect 6150 13030 6196 13082
rect 5900 13028 5956 13030
rect 5980 13028 6036 13030
rect 6060 13028 6116 13030
rect 6140 13028 6196 13030
rect 5900 11994 5956 11996
rect 5980 11994 6036 11996
rect 6060 11994 6116 11996
rect 6140 11994 6196 11996
rect 5900 11942 5946 11994
rect 5946 11942 5956 11994
rect 5980 11942 6010 11994
rect 6010 11942 6022 11994
rect 6022 11942 6036 11994
rect 6060 11942 6074 11994
rect 6074 11942 6086 11994
rect 6086 11942 6116 11994
rect 6140 11942 6150 11994
rect 6150 11942 6196 11994
rect 5900 11940 5956 11942
rect 5980 11940 6036 11942
rect 6060 11940 6116 11942
rect 6140 11940 6196 11942
rect 3428 6010 3484 6012
rect 3508 6010 3564 6012
rect 3588 6010 3644 6012
rect 3668 6010 3724 6012
rect 3428 5958 3474 6010
rect 3474 5958 3484 6010
rect 3508 5958 3538 6010
rect 3538 5958 3550 6010
rect 3550 5958 3564 6010
rect 3588 5958 3602 6010
rect 3602 5958 3614 6010
rect 3614 5958 3644 6010
rect 3668 5958 3678 6010
rect 3678 5958 3724 6010
rect 3428 5956 3484 5958
rect 3508 5956 3564 5958
rect 3588 5956 3644 5958
rect 3668 5956 3724 5958
rect 2778 5092 2834 5128
rect 2778 5072 2780 5092
rect 2780 5072 2832 5092
rect 2832 5072 2834 5092
rect 2962 5072 3018 5128
rect 3428 4922 3484 4924
rect 3508 4922 3564 4924
rect 3588 4922 3644 4924
rect 3668 4922 3724 4924
rect 3428 4870 3474 4922
rect 3474 4870 3484 4922
rect 3508 4870 3538 4922
rect 3538 4870 3550 4922
rect 3550 4870 3564 4922
rect 3588 4870 3602 4922
rect 3602 4870 3614 4922
rect 3614 4870 3644 4922
rect 3668 4870 3678 4922
rect 3678 4870 3724 4922
rect 3428 4868 3484 4870
rect 3508 4868 3564 4870
rect 3588 4868 3644 4870
rect 3668 4868 3724 4870
rect 3428 3834 3484 3836
rect 3508 3834 3564 3836
rect 3588 3834 3644 3836
rect 3668 3834 3724 3836
rect 3428 3782 3474 3834
rect 3474 3782 3484 3834
rect 3508 3782 3538 3834
rect 3538 3782 3550 3834
rect 3550 3782 3564 3834
rect 3588 3782 3602 3834
rect 3602 3782 3614 3834
rect 3614 3782 3644 3834
rect 3668 3782 3678 3834
rect 3678 3782 3724 3834
rect 3428 3780 3484 3782
rect 3508 3780 3564 3782
rect 3588 3780 3644 3782
rect 3668 3780 3724 3782
rect 3146 3576 3202 3632
rect 3428 2746 3484 2748
rect 3508 2746 3564 2748
rect 3588 2746 3644 2748
rect 3668 2746 3724 2748
rect 3428 2694 3474 2746
rect 3474 2694 3484 2746
rect 3508 2694 3538 2746
rect 3538 2694 3550 2746
rect 3550 2694 3564 2746
rect 3588 2694 3602 2746
rect 3602 2694 3614 2746
rect 3614 2694 3644 2746
rect 3668 2694 3678 2746
rect 3678 2694 3724 2746
rect 3428 2692 3484 2694
rect 3508 2692 3564 2694
rect 3588 2692 3644 2694
rect 3668 2692 3724 2694
rect 5900 10906 5956 10908
rect 5980 10906 6036 10908
rect 6060 10906 6116 10908
rect 6140 10906 6196 10908
rect 5900 10854 5946 10906
rect 5946 10854 5956 10906
rect 5980 10854 6010 10906
rect 6010 10854 6022 10906
rect 6022 10854 6036 10906
rect 6060 10854 6074 10906
rect 6074 10854 6086 10906
rect 6086 10854 6116 10906
rect 6140 10854 6150 10906
rect 6150 10854 6196 10906
rect 5900 10852 5956 10854
rect 5980 10852 6036 10854
rect 6060 10852 6116 10854
rect 6140 10852 6196 10854
rect 5900 9818 5956 9820
rect 5980 9818 6036 9820
rect 6060 9818 6116 9820
rect 6140 9818 6196 9820
rect 5900 9766 5946 9818
rect 5946 9766 5956 9818
rect 5980 9766 6010 9818
rect 6010 9766 6022 9818
rect 6022 9766 6036 9818
rect 6060 9766 6074 9818
rect 6074 9766 6086 9818
rect 6086 9766 6116 9818
rect 6140 9766 6150 9818
rect 6150 9766 6196 9818
rect 5900 9764 5956 9766
rect 5980 9764 6036 9766
rect 6060 9764 6116 9766
rect 6140 9764 6196 9766
rect 5900 8730 5956 8732
rect 5980 8730 6036 8732
rect 6060 8730 6116 8732
rect 6140 8730 6196 8732
rect 5900 8678 5946 8730
rect 5946 8678 5956 8730
rect 5980 8678 6010 8730
rect 6010 8678 6022 8730
rect 6022 8678 6036 8730
rect 6060 8678 6074 8730
rect 6074 8678 6086 8730
rect 6086 8678 6116 8730
rect 6140 8678 6150 8730
rect 6150 8678 6196 8730
rect 5900 8676 5956 8678
rect 5980 8676 6036 8678
rect 6060 8676 6116 8678
rect 6140 8676 6196 8678
rect 10845 16346 10901 16348
rect 10925 16346 10981 16348
rect 11005 16346 11061 16348
rect 11085 16346 11141 16348
rect 10845 16294 10891 16346
rect 10891 16294 10901 16346
rect 10925 16294 10955 16346
rect 10955 16294 10967 16346
rect 10967 16294 10981 16346
rect 11005 16294 11019 16346
rect 11019 16294 11031 16346
rect 11031 16294 11061 16346
rect 11085 16294 11095 16346
rect 11095 16294 11141 16346
rect 10845 16292 10901 16294
rect 10925 16292 10981 16294
rect 11005 16292 11061 16294
rect 11085 16292 11141 16294
rect 8373 15802 8429 15804
rect 8453 15802 8509 15804
rect 8533 15802 8589 15804
rect 8613 15802 8669 15804
rect 8373 15750 8419 15802
rect 8419 15750 8429 15802
rect 8453 15750 8483 15802
rect 8483 15750 8495 15802
rect 8495 15750 8509 15802
rect 8533 15750 8547 15802
rect 8547 15750 8559 15802
rect 8559 15750 8589 15802
rect 8613 15750 8623 15802
rect 8623 15750 8669 15802
rect 8373 15748 8429 15750
rect 8453 15748 8509 15750
rect 8533 15748 8589 15750
rect 8613 15748 8669 15750
rect 8373 14714 8429 14716
rect 8453 14714 8509 14716
rect 8533 14714 8589 14716
rect 8613 14714 8669 14716
rect 8373 14662 8419 14714
rect 8419 14662 8429 14714
rect 8453 14662 8483 14714
rect 8483 14662 8495 14714
rect 8495 14662 8509 14714
rect 8533 14662 8547 14714
rect 8547 14662 8559 14714
rect 8559 14662 8589 14714
rect 8613 14662 8623 14714
rect 8623 14662 8669 14714
rect 8373 14660 8429 14662
rect 8453 14660 8509 14662
rect 8533 14660 8589 14662
rect 8613 14660 8669 14662
rect 5900 7642 5956 7644
rect 5980 7642 6036 7644
rect 6060 7642 6116 7644
rect 6140 7642 6196 7644
rect 5900 7590 5946 7642
rect 5946 7590 5956 7642
rect 5980 7590 6010 7642
rect 6010 7590 6022 7642
rect 6022 7590 6036 7642
rect 6060 7590 6074 7642
rect 6074 7590 6086 7642
rect 6086 7590 6116 7642
rect 6140 7590 6150 7642
rect 6150 7590 6196 7642
rect 5900 7588 5956 7590
rect 5980 7588 6036 7590
rect 6060 7588 6116 7590
rect 6140 7588 6196 7590
rect 5900 6554 5956 6556
rect 5980 6554 6036 6556
rect 6060 6554 6116 6556
rect 6140 6554 6196 6556
rect 5900 6502 5946 6554
rect 5946 6502 5956 6554
rect 5980 6502 6010 6554
rect 6010 6502 6022 6554
rect 6022 6502 6036 6554
rect 6060 6502 6074 6554
rect 6074 6502 6086 6554
rect 6086 6502 6116 6554
rect 6140 6502 6150 6554
rect 6150 6502 6196 6554
rect 5900 6500 5956 6502
rect 5980 6500 6036 6502
rect 6060 6500 6116 6502
rect 6140 6500 6196 6502
rect 5900 5466 5956 5468
rect 5980 5466 6036 5468
rect 6060 5466 6116 5468
rect 6140 5466 6196 5468
rect 5900 5414 5946 5466
rect 5946 5414 5956 5466
rect 5980 5414 6010 5466
rect 6010 5414 6022 5466
rect 6022 5414 6036 5466
rect 6060 5414 6074 5466
rect 6074 5414 6086 5466
rect 6086 5414 6116 5466
rect 6140 5414 6150 5466
rect 6150 5414 6196 5466
rect 5900 5412 5956 5414
rect 5980 5412 6036 5414
rect 6060 5412 6116 5414
rect 6140 5412 6196 5414
rect 8373 13626 8429 13628
rect 8453 13626 8509 13628
rect 8533 13626 8589 13628
rect 8613 13626 8669 13628
rect 8373 13574 8419 13626
rect 8419 13574 8429 13626
rect 8453 13574 8483 13626
rect 8483 13574 8495 13626
rect 8495 13574 8509 13626
rect 8533 13574 8547 13626
rect 8547 13574 8559 13626
rect 8559 13574 8589 13626
rect 8613 13574 8623 13626
rect 8623 13574 8669 13626
rect 8373 13572 8429 13574
rect 8453 13572 8509 13574
rect 8533 13572 8589 13574
rect 8613 13572 8669 13574
rect 8373 12538 8429 12540
rect 8453 12538 8509 12540
rect 8533 12538 8589 12540
rect 8613 12538 8669 12540
rect 8373 12486 8419 12538
rect 8419 12486 8429 12538
rect 8453 12486 8483 12538
rect 8483 12486 8495 12538
rect 8495 12486 8509 12538
rect 8533 12486 8547 12538
rect 8547 12486 8559 12538
rect 8559 12486 8589 12538
rect 8613 12486 8623 12538
rect 8623 12486 8669 12538
rect 8373 12484 8429 12486
rect 8453 12484 8509 12486
rect 8533 12484 8589 12486
rect 8613 12484 8669 12486
rect 8373 11450 8429 11452
rect 8453 11450 8509 11452
rect 8533 11450 8589 11452
rect 8613 11450 8669 11452
rect 8373 11398 8419 11450
rect 8419 11398 8429 11450
rect 8453 11398 8483 11450
rect 8483 11398 8495 11450
rect 8495 11398 8509 11450
rect 8533 11398 8547 11450
rect 8547 11398 8559 11450
rect 8559 11398 8589 11450
rect 8613 11398 8623 11450
rect 8623 11398 8669 11450
rect 8373 11396 8429 11398
rect 8453 11396 8509 11398
rect 8533 11396 8589 11398
rect 8613 11396 8669 11398
rect 8373 10362 8429 10364
rect 8453 10362 8509 10364
rect 8533 10362 8589 10364
rect 8613 10362 8669 10364
rect 8373 10310 8419 10362
rect 8419 10310 8429 10362
rect 8453 10310 8483 10362
rect 8483 10310 8495 10362
rect 8495 10310 8509 10362
rect 8533 10310 8547 10362
rect 8547 10310 8559 10362
rect 8559 10310 8589 10362
rect 8613 10310 8623 10362
rect 8623 10310 8669 10362
rect 8373 10308 8429 10310
rect 8453 10308 8509 10310
rect 8533 10308 8589 10310
rect 8613 10308 8669 10310
rect 8373 9274 8429 9276
rect 8453 9274 8509 9276
rect 8533 9274 8589 9276
rect 8613 9274 8669 9276
rect 8373 9222 8419 9274
rect 8419 9222 8429 9274
rect 8453 9222 8483 9274
rect 8483 9222 8495 9274
rect 8495 9222 8509 9274
rect 8533 9222 8547 9274
rect 8547 9222 8559 9274
rect 8559 9222 8589 9274
rect 8613 9222 8623 9274
rect 8623 9222 8669 9274
rect 8373 9220 8429 9222
rect 8453 9220 8509 9222
rect 8533 9220 8589 9222
rect 8613 9220 8669 9222
rect 8373 8186 8429 8188
rect 8453 8186 8509 8188
rect 8533 8186 8589 8188
rect 8613 8186 8669 8188
rect 8373 8134 8419 8186
rect 8419 8134 8429 8186
rect 8453 8134 8483 8186
rect 8483 8134 8495 8186
rect 8495 8134 8509 8186
rect 8533 8134 8547 8186
rect 8547 8134 8559 8186
rect 8559 8134 8589 8186
rect 8613 8134 8623 8186
rect 8623 8134 8669 8186
rect 8373 8132 8429 8134
rect 8453 8132 8509 8134
rect 8533 8132 8589 8134
rect 8613 8132 8669 8134
rect 8373 7098 8429 7100
rect 8453 7098 8509 7100
rect 8533 7098 8589 7100
rect 8613 7098 8669 7100
rect 8373 7046 8419 7098
rect 8419 7046 8429 7098
rect 8453 7046 8483 7098
rect 8483 7046 8495 7098
rect 8495 7046 8509 7098
rect 8533 7046 8547 7098
rect 8547 7046 8559 7098
rect 8559 7046 8589 7098
rect 8613 7046 8623 7098
rect 8623 7046 8669 7098
rect 8373 7044 8429 7046
rect 8453 7044 8509 7046
rect 8533 7044 8589 7046
rect 8613 7044 8669 7046
rect 5900 4378 5956 4380
rect 5980 4378 6036 4380
rect 6060 4378 6116 4380
rect 6140 4378 6196 4380
rect 5900 4326 5946 4378
rect 5946 4326 5956 4378
rect 5980 4326 6010 4378
rect 6010 4326 6022 4378
rect 6022 4326 6036 4378
rect 6060 4326 6074 4378
rect 6074 4326 6086 4378
rect 6086 4326 6116 4378
rect 6140 4326 6150 4378
rect 6150 4326 6196 4378
rect 5900 4324 5956 4326
rect 5980 4324 6036 4326
rect 6060 4324 6116 4326
rect 6140 4324 6196 4326
rect 5900 3290 5956 3292
rect 5980 3290 6036 3292
rect 6060 3290 6116 3292
rect 6140 3290 6196 3292
rect 5900 3238 5946 3290
rect 5946 3238 5956 3290
rect 5980 3238 6010 3290
rect 6010 3238 6022 3290
rect 6022 3238 6036 3290
rect 6060 3238 6074 3290
rect 6074 3238 6086 3290
rect 6086 3238 6116 3290
rect 6140 3238 6150 3290
rect 6150 3238 6196 3290
rect 5900 3236 5956 3238
rect 5980 3236 6036 3238
rect 6060 3236 6116 3238
rect 6140 3236 6196 3238
rect 9678 12164 9734 12200
rect 9678 12144 9680 12164
rect 9680 12144 9732 12164
rect 9732 12144 9734 12164
rect 10845 15258 10901 15260
rect 10925 15258 10981 15260
rect 11005 15258 11061 15260
rect 11085 15258 11141 15260
rect 10845 15206 10891 15258
rect 10891 15206 10901 15258
rect 10925 15206 10955 15258
rect 10955 15206 10967 15258
rect 10967 15206 10981 15258
rect 11005 15206 11019 15258
rect 11019 15206 11031 15258
rect 11031 15206 11061 15258
rect 11085 15206 11095 15258
rect 11095 15206 11141 15258
rect 10845 15204 10901 15206
rect 10925 15204 10981 15206
rect 11005 15204 11061 15206
rect 11085 15204 11141 15206
rect 10845 14170 10901 14172
rect 10925 14170 10981 14172
rect 11005 14170 11061 14172
rect 11085 14170 11141 14172
rect 10845 14118 10891 14170
rect 10891 14118 10901 14170
rect 10925 14118 10955 14170
rect 10955 14118 10967 14170
rect 10967 14118 10981 14170
rect 11005 14118 11019 14170
rect 11019 14118 11031 14170
rect 11031 14118 11061 14170
rect 11085 14118 11095 14170
rect 11095 14118 11141 14170
rect 10845 14116 10901 14118
rect 10925 14116 10981 14118
rect 11005 14116 11061 14118
rect 11085 14116 11141 14118
rect 10845 13082 10901 13084
rect 10925 13082 10981 13084
rect 11005 13082 11061 13084
rect 11085 13082 11141 13084
rect 10845 13030 10891 13082
rect 10891 13030 10901 13082
rect 10925 13030 10955 13082
rect 10955 13030 10967 13082
rect 10967 13030 10981 13082
rect 11005 13030 11019 13082
rect 11019 13030 11031 13082
rect 11031 13030 11061 13082
rect 11085 13030 11095 13082
rect 11095 13030 11141 13082
rect 10845 13028 10901 13030
rect 10925 13028 10981 13030
rect 11005 13028 11061 13030
rect 11085 13028 11141 13030
rect 10845 11994 10901 11996
rect 10925 11994 10981 11996
rect 11005 11994 11061 11996
rect 11085 11994 11141 11996
rect 10845 11942 10891 11994
rect 10891 11942 10901 11994
rect 10925 11942 10955 11994
rect 10955 11942 10967 11994
rect 10967 11942 10981 11994
rect 11005 11942 11019 11994
rect 11019 11942 11031 11994
rect 11031 11942 11061 11994
rect 11085 11942 11095 11994
rect 11095 11942 11141 11994
rect 10845 11940 10901 11942
rect 10925 11940 10981 11942
rect 11005 11940 11061 11942
rect 11085 11940 11141 11942
rect 10845 10906 10901 10908
rect 10925 10906 10981 10908
rect 11005 10906 11061 10908
rect 11085 10906 11141 10908
rect 10845 10854 10891 10906
rect 10891 10854 10901 10906
rect 10925 10854 10955 10906
rect 10955 10854 10967 10906
rect 10967 10854 10981 10906
rect 11005 10854 11019 10906
rect 11019 10854 11031 10906
rect 11031 10854 11061 10906
rect 11085 10854 11095 10906
rect 11095 10854 11141 10906
rect 10845 10852 10901 10854
rect 10925 10852 10981 10854
rect 11005 10852 11061 10854
rect 11085 10852 11141 10854
rect 13318 15802 13374 15804
rect 13398 15802 13454 15804
rect 13478 15802 13534 15804
rect 13558 15802 13614 15804
rect 13318 15750 13364 15802
rect 13364 15750 13374 15802
rect 13398 15750 13428 15802
rect 13428 15750 13440 15802
rect 13440 15750 13454 15802
rect 13478 15750 13492 15802
rect 13492 15750 13504 15802
rect 13504 15750 13534 15802
rect 13558 15750 13568 15802
rect 13568 15750 13614 15802
rect 13318 15748 13374 15750
rect 13398 15748 13454 15750
rect 13478 15748 13534 15750
rect 13558 15748 13614 15750
rect 10845 9818 10901 9820
rect 10925 9818 10981 9820
rect 11005 9818 11061 9820
rect 11085 9818 11141 9820
rect 10845 9766 10891 9818
rect 10891 9766 10901 9818
rect 10925 9766 10955 9818
rect 10955 9766 10967 9818
rect 10967 9766 10981 9818
rect 11005 9766 11019 9818
rect 11019 9766 11031 9818
rect 11031 9766 11061 9818
rect 11085 9766 11095 9818
rect 11095 9766 11141 9818
rect 10845 9764 10901 9766
rect 10925 9764 10981 9766
rect 11005 9764 11061 9766
rect 11085 9764 11141 9766
rect 13318 14714 13374 14716
rect 13398 14714 13454 14716
rect 13478 14714 13534 14716
rect 13558 14714 13614 14716
rect 13318 14662 13364 14714
rect 13364 14662 13374 14714
rect 13398 14662 13428 14714
rect 13428 14662 13440 14714
rect 13440 14662 13454 14714
rect 13478 14662 13492 14714
rect 13492 14662 13504 14714
rect 13504 14662 13534 14714
rect 13558 14662 13568 14714
rect 13568 14662 13614 14714
rect 13318 14660 13374 14662
rect 13398 14660 13454 14662
rect 13478 14660 13534 14662
rect 13558 14660 13614 14662
rect 13358 14356 13360 14376
rect 13360 14356 13412 14376
rect 13412 14356 13414 14376
rect 13358 14320 13414 14356
rect 13318 13626 13374 13628
rect 13398 13626 13454 13628
rect 13478 13626 13534 13628
rect 13558 13626 13614 13628
rect 13318 13574 13364 13626
rect 13364 13574 13374 13626
rect 13398 13574 13428 13626
rect 13428 13574 13440 13626
rect 13440 13574 13454 13626
rect 13478 13574 13492 13626
rect 13492 13574 13504 13626
rect 13504 13574 13534 13626
rect 13558 13574 13568 13626
rect 13568 13574 13614 13626
rect 13318 13572 13374 13574
rect 13398 13572 13454 13574
rect 13478 13572 13534 13574
rect 13558 13572 13614 13574
rect 13318 12538 13374 12540
rect 13398 12538 13454 12540
rect 13478 12538 13534 12540
rect 13558 12538 13614 12540
rect 13318 12486 13364 12538
rect 13364 12486 13374 12538
rect 13398 12486 13428 12538
rect 13428 12486 13440 12538
rect 13440 12486 13454 12538
rect 13478 12486 13492 12538
rect 13492 12486 13504 12538
rect 13504 12486 13534 12538
rect 13558 12486 13568 12538
rect 13568 12486 13614 12538
rect 13318 12484 13374 12486
rect 13398 12484 13454 12486
rect 13478 12484 13534 12486
rect 13558 12484 13614 12486
rect 13450 12280 13506 12336
rect 13318 11450 13374 11452
rect 13398 11450 13454 11452
rect 13478 11450 13534 11452
rect 13558 11450 13614 11452
rect 13318 11398 13364 11450
rect 13364 11398 13374 11450
rect 13398 11398 13428 11450
rect 13428 11398 13440 11450
rect 13440 11398 13454 11450
rect 13478 11398 13492 11450
rect 13492 11398 13504 11450
rect 13504 11398 13534 11450
rect 13558 11398 13568 11450
rect 13568 11398 13614 11450
rect 13318 11396 13374 11398
rect 13398 11396 13454 11398
rect 13478 11396 13534 11398
rect 13558 11396 13614 11398
rect 13318 10362 13374 10364
rect 13398 10362 13454 10364
rect 13478 10362 13534 10364
rect 13558 10362 13614 10364
rect 13318 10310 13364 10362
rect 13364 10310 13374 10362
rect 13398 10310 13428 10362
rect 13428 10310 13440 10362
rect 13440 10310 13454 10362
rect 13478 10310 13492 10362
rect 13492 10310 13504 10362
rect 13504 10310 13534 10362
rect 13558 10310 13568 10362
rect 13568 10310 13614 10362
rect 13318 10308 13374 10310
rect 13398 10308 13454 10310
rect 13478 10308 13534 10310
rect 13558 10308 13614 10310
rect 10845 8730 10901 8732
rect 10925 8730 10981 8732
rect 11005 8730 11061 8732
rect 11085 8730 11141 8732
rect 10845 8678 10891 8730
rect 10891 8678 10901 8730
rect 10925 8678 10955 8730
rect 10955 8678 10967 8730
rect 10967 8678 10981 8730
rect 11005 8678 11019 8730
rect 11019 8678 11031 8730
rect 11031 8678 11061 8730
rect 11085 8678 11095 8730
rect 11095 8678 11141 8730
rect 10845 8676 10901 8678
rect 10925 8676 10981 8678
rect 11005 8676 11061 8678
rect 11085 8676 11141 8678
rect 13318 9274 13374 9276
rect 13398 9274 13454 9276
rect 13478 9274 13534 9276
rect 13558 9274 13614 9276
rect 13318 9222 13364 9274
rect 13364 9222 13374 9274
rect 13398 9222 13428 9274
rect 13428 9222 13440 9274
rect 13440 9222 13454 9274
rect 13478 9222 13492 9274
rect 13492 9222 13504 9274
rect 13504 9222 13534 9274
rect 13558 9222 13568 9274
rect 13568 9222 13614 9274
rect 13318 9220 13374 9222
rect 13398 9220 13454 9222
rect 13478 9220 13534 9222
rect 13558 9220 13614 9222
rect 10845 7642 10901 7644
rect 10925 7642 10981 7644
rect 11005 7642 11061 7644
rect 11085 7642 11141 7644
rect 10845 7590 10891 7642
rect 10891 7590 10901 7642
rect 10925 7590 10955 7642
rect 10955 7590 10967 7642
rect 10967 7590 10981 7642
rect 11005 7590 11019 7642
rect 11019 7590 11031 7642
rect 11031 7590 11061 7642
rect 11085 7590 11095 7642
rect 11095 7590 11141 7642
rect 10845 7588 10901 7590
rect 10925 7588 10981 7590
rect 11005 7588 11061 7590
rect 11085 7588 11141 7590
rect 10845 6554 10901 6556
rect 10925 6554 10981 6556
rect 11005 6554 11061 6556
rect 11085 6554 11141 6556
rect 10845 6502 10891 6554
rect 10891 6502 10901 6554
rect 10925 6502 10955 6554
rect 10955 6502 10967 6554
rect 10967 6502 10981 6554
rect 11005 6502 11019 6554
rect 11019 6502 11031 6554
rect 11031 6502 11061 6554
rect 11085 6502 11095 6554
rect 11095 6502 11141 6554
rect 10845 6500 10901 6502
rect 10925 6500 10981 6502
rect 11005 6500 11061 6502
rect 11085 6500 11141 6502
rect 8373 6010 8429 6012
rect 8453 6010 8509 6012
rect 8533 6010 8589 6012
rect 8613 6010 8669 6012
rect 8373 5958 8419 6010
rect 8419 5958 8429 6010
rect 8453 5958 8483 6010
rect 8483 5958 8495 6010
rect 8495 5958 8509 6010
rect 8533 5958 8547 6010
rect 8547 5958 8559 6010
rect 8559 5958 8589 6010
rect 8613 5958 8623 6010
rect 8623 5958 8669 6010
rect 8373 5956 8429 5958
rect 8453 5956 8509 5958
rect 8533 5956 8589 5958
rect 8613 5956 8669 5958
rect 10845 5466 10901 5468
rect 10925 5466 10981 5468
rect 11005 5466 11061 5468
rect 11085 5466 11141 5468
rect 10845 5414 10891 5466
rect 10891 5414 10901 5466
rect 10925 5414 10955 5466
rect 10955 5414 10967 5466
rect 10967 5414 10981 5466
rect 11005 5414 11019 5466
rect 11019 5414 11031 5466
rect 11031 5414 11061 5466
rect 11085 5414 11095 5466
rect 11095 5414 11141 5466
rect 10845 5412 10901 5414
rect 10925 5412 10981 5414
rect 11005 5412 11061 5414
rect 11085 5412 11141 5414
rect 11150 5208 11206 5264
rect 13318 8186 13374 8188
rect 13398 8186 13454 8188
rect 13478 8186 13534 8188
rect 13558 8186 13614 8188
rect 13318 8134 13364 8186
rect 13364 8134 13374 8186
rect 13398 8134 13428 8186
rect 13428 8134 13440 8186
rect 13440 8134 13454 8186
rect 13478 8134 13492 8186
rect 13492 8134 13504 8186
rect 13504 8134 13534 8186
rect 13558 8134 13568 8186
rect 13568 8134 13614 8186
rect 13318 8132 13374 8134
rect 13398 8132 13454 8134
rect 13478 8132 13534 8134
rect 13558 8132 13614 8134
rect 13318 7098 13374 7100
rect 13398 7098 13454 7100
rect 13478 7098 13534 7100
rect 13558 7098 13614 7100
rect 13318 7046 13364 7098
rect 13364 7046 13374 7098
rect 13398 7046 13428 7098
rect 13428 7046 13440 7098
rect 13440 7046 13454 7098
rect 13478 7046 13492 7098
rect 13492 7046 13504 7098
rect 13504 7046 13534 7098
rect 13558 7046 13568 7098
rect 13568 7046 13614 7098
rect 13318 7044 13374 7046
rect 13398 7044 13454 7046
rect 13478 7044 13534 7046
rect 13558 7044 13614 7046
rect 13318 6010 13374 6012
rect 13398 6010 13454 6012
rect 13478 6010 13534 6012
rect 13558 6010 13614 6012
rect 13318 5958 13364 6010
rect 13364 5958 13374 6010
rect 13398 5958 13428 6010
rect 13428 5958 13440 6010
rect 13440 5958 13454 6010
rect 13478 5958 13492 6010
rect 13492 5958 13504 6010
rect 13504 5958 13534 6010
rect 13558 5958 13568 6010
rect 13568 5958 13614 6010
rect 13318 5956 13374 5958
rect 13398 5956 13454 5958
rect 13478 5956 13534 5958
rect 13558 5956 13614 5958
rect 15790 16346 15846 16348
rect 15870 16346 15926 16348
rect 15950 16346 16006 16348
rect 16030 16346 16086 16348
rect 15790 16294 15836 16346
rect 15836 16294 15846 16346
rect 15870 16294 15900 16346
rect 15900 16294 15912 16346
rect 15912 16294 15926 16346
rect 15950 16294 15964 16346
rect 15964 16294 15976 16346
rect 15976 16294 16006 16346
rect 16030 16294 16040 16346
rect 16040 16294 16086 16346
rect 15790 16292 15846 16294
rect 15870 16292 15926 16294
rect 15950 16292 16006 16294
rect 16030 16292 16086 16294
rect 20735 16346 20791 16348
rect 20815 16346 20871 16348
rect 20895 16346 20951 16348
rect 20975 16346 21031 16348
rect 20735 16294 20781 16346
rect 20781 16294 20791 16346
rect 20815 16294 20845 16346
rect 20845 16294 20857 16346
rect 20857 16294 20871 16346
rect 20895 16294 20909 16346
rect 20909 16294 20921 16346
rect 20921 16294 20951 16346
rect 20975 16294 20985 16346
rect 20985 16294 21031 16346
rect 20735 16292 20791 16294
rect 20815 16292 20871 16294
rect 20895 16292 20951 16294
rect 20975 16292 21031 16294
rect 15290 14048 15346 14104
rect 15790 15258 15846 15260
rect 15870 15258 15926 15260
rect 15950 15258 16006 15260
rect 16030 15258 16086 15260
rect 15790 15206 15836 15258
rect 15836 15206 15846 15258
rect 15870 15206 15900 15258
rect 15900 15206 15912 15258
rect 15912 15206 15926 15258
rect 15950 15206 15964 15258
rect 15964 15206 15976 15258
rect 15976 15206 16006 15258
rect 16030 15206 16040 15258
rect 16040 15206 16086 15258
rect 15790 15204 15846 15206
rect 15870 15204 15926 15206
rect 15950 15204 16006 15206
rect 16030 15204 16086 15206
rect 15790 14170 15846 14172
rect 15870 14170 15926 14172
rect 15950 14170 16006 14172
rect 16030 14170 16086 14172
rect 15790 14118 15836 14170
rect 15836 14118 15846 14170
rect 15870 14118 15900 14170
rect 15900 14118 15912 14170
rect 15912 14118 15926 14170
rect 15950 14118 15964 14170
rect 15964 14118 15976 14170
rect 15976 14118 16006 14170
rect 16030 14118 16040 14170
rect 16040 14118 16086 14170
rect 15790 14116 15846 14118
rect 15870 14116 15926 14118
rect 15950 14116 16006 14118
rect 16030 14116 16086 14118
rect 15658 13776 15714 13832
rect 15790 13082 15846 13084
rect 15870 13082 15926 13084
rect 15950 13082 16006 13084
rect 16030 13082 16086 13084
rect 15790 13030 15836 13082
rect 15836 13030 15846 13082
rect 15870 13030 15900 13082
rect 15900 13030 15912 13082
rect 15912 13030 15926 13082
rect 15950 13030 15964 13082
rect 15964 13030 15976 13082
rect 15976 13030 16006 13082
rect 16030 13030 16040 13082
rect 16040 13030 16086 13082
rect 15790 13028 15846 13030
rect 15870 13028 15926 13030
rect 15950 13028 16006 13030
rect 16030 13028 16086 13030
rect 15790 11994 15846 11996
rect 15870 11994 15926 11996
rect 15950 11994 16006 11996
rect 16030 11994 16086 11996
rect 15790 11942 15836 11994
rect 15836 11942 15846 11994
rect 15870 11942 15900 11994
rect 15900 11942 15912 11994
rect 15912 11942 15926 11994
rect 15950 11942 15964 11994
rect 15964 11942 15976 11994
rect 15976 11942 16006 11994
rect 16030 11942 16040 11994
rect 16040 11942 16086 11994
rect 15790 11940 15846 11942
rect 15870 11940 15926 11942
rect 15950 11940 16006 11942
rect 16030 11940 16086 11942
rect 15790 10906 15846 10908
rect 15870 10906 15926 10908
rect 15950 10906 16006 10908
rect 16030 10906 16086 10908
rect 15790 10854 15836 10906
rect 15836 10854 15846 10906
rect 15870 10854 15900 10906
rect 15900 10854 15912 10906
rect 15912 10854 15926 10906
rect 15950 10854 15964 10906
rect 15964 10854 15976 10906
rect 15976 10854 16006 10906
rect 16030 10854 16040 10906
rect 16040 10854 16086 10906
rect 15790 10852 15846 10854
rect 15870 10852 15926 10854
rect 15950 10852 16006 10854
rect 16030 10852 16086 10854
rect 15790 9818 15846 9820
rect 15870 9818 15926 9820
rect 15950 9818 16006 9820
rect 16030 9818 16086 9820
rect 15790 9766 15836 9818
rect 15836 9766 15846 9818
rect 15870 9766 15900 9818
rect 15900 9766 15912 9818
rect 15912 9766 15926 9818
rect 15950 9766 15964 9818
rect 15964 9766 15976 9818
rect 15976 9766 16006 9818
rect 16030 9766 16040 9818
rect 16040 9766 16086 9818
rect 15790 9764 15846 9766
rect 15870 9764 15926 9766
rect 15950 9764 16006 9766
rect 16030 9764 16086 9766
rect 15790 8730 15846 8732
rect 15870 8730 15926 8732
rect 15950 8730 16006 8732
rect 16030 8730 16086 8732
rect 15790 8678 15836 8730
rect 15836 8678 15846 8730
rect 15870 8678 15900 8730
rect 15900 8678 15912 8730
rect 15912 8678 15926 8730
rect 15950 8678 15964 8730
rect 15964 8678 15976 8730
rect 15976 8678 16006 8730
rect 16030 8678 16040 8730
rect 16040 8678 16086 8730
rect 15790 8676 15846 8678
rect 15870 8676 15926 8678
rect 15950 8676 16006 8678
rect 16030 8676 16086 8678
rect 18263 15802 18319 15804
rect 18343 15802 18399 15804
rect 18423 15802 18479 15804
rect 18503 15802 18559 15804
rect 18263 15750 18309 15802
rect 18309 15750 18319 15802
rect 18343 15750 18373 15802
rect 18373 15750 18385 15802
rect 18385 15750 18399 15802
rect 18423 15750 18437 15802
rect 18437 15750 18449 15802
rect 18449 15750 18479 15802
rect 18503 15750 18513 15802
rect 18513 15750 18559 15802
rect 18263 15748 18319 15750
rect 18343 15748 18399 15750
rect 18423 15748 18479 15750
rect 18503 15748 18559 15750
rect 16578 12300 16634 12336
rect 16578 12280 16580 12300
rect 16580 12280 16632 12300
rect 16632 12280 16634 12300
rect 20735 15258 20791 15260
rect 20815 15258 20871 15260
rect 20895 15258 20951 15260
rect 20975 15258 21031 15260
rect 20735 15206 20781 15258
rect 20781 15206 20791 15258
rect 20815 15206 20845 15258
rect 20845 15206 20857 15258
rect 20857 15206 20871 15258
rect 20895 15206 20909 15258
rect 20909 15206 20921 15258
rect 20921 15206 20951 15258
rect 20975 15206 20985 15258
rect 20985 15206 21031 15258
rect 20735 15204 20791 15206
rect 20815 15204 20871 15206
rect 20895 15204 20951 15206
rect 20975 15204 21031 15206
rect 17866 14320 17922 14376
rect 18263 14714 18319 14716
rect 18343 14714 18399 14716
rect 18423 14714 18479 14716
rect 18503 14714 18559 14716
rect 18263 14662 18309 14714
rect 18309 14662 18319 14714
rect 18343 14662 18373 14714
rect 18373 14662 18385 14714
rect 18385 14662 18399 14714
rect 18423 14662 18437 14714
rect 18437 14662 18449 14714
rect 18449 14662 18479 14714
rect 18503 14662 18513 14714
rect 18513 14662 18559 14714
rect 18263 14660 18319 14662
rect 18343 14660 18399 14662
rect 18423 14660 18479 14662
rect 18503 14660 18559 14662
rect 18234 14356 18236 14376
rect 18236 14356 18288 14376
rect 18288 14356 18290 14376
rect 18234 14320 18290 14356
rect 18263 13626 18319 13628
rect 18343 13626 18399 13628
rect 18423 13626 18479 13628
rect 18503 13626 18559 13628
rect 18263 13574 18309 13626
rect 18309 13574 18319 13626
rect 18343 13574 18373 13626
rect 18373 13574 18385 13626
rect 18385 13574 18399 13626
rect 18423 13574 18437 13626
rect 18437 13574 18449 13626
rect 18449 13574 18479 13626
rect 18503 13574 18513 13626
rect 18513 13574 18559 13626
rect 18263 13572 18319 13574
rect 18343 13572 18399 13574
rect 18423 13572 18479 13574
rect 18503 13572 18559 13574
rect 18263 12538 18319 12540
rect 18343 12538 18399 12540
rect 18423 12538 18479 12540
rect 18503 12538 18559 12540
rect 18263 12486 18309 12538
rect 18309 12486 18319 12538
rect 18343 12486 18373 12538
rect 18373 12486 18385 12538
rect 18385 12486 18399 12538
rect 18423 12486 18437 12538
rect 18437 12486 18449 12538
rect 18449 12486 18479 12538
rect 18503 12486 18513 12538
rect 18513 12486 18559 12538
rect 18263 12484 18319 12486
rect 18343 12484 18399 12486
rect 18423 12484 18479 12486
rect 18503 12484 18559 12486
rect 19430 12144 19486 12200
rect 18263 11450 18319 11452
rect 18343 11450 18399 11452
rect 18423 11450 18479 11452
rect 18503 11450 18559 11452
rect 18263 11398 18309 11450
rect 18309 11398 18319 11450
rect 18343 11398 18373 11450
rect 18373 11398 18385 11450
rect 18385 11398 18399 11450
rect 18423 11398 18437 11450
rect 18437 11398 18449 11450
rect 18449 11398 18479 11450
rect 18503 11398 18513 11450
rect 18513 11398 18559 11450
rect 18263 11396 18319 11398
rect 18343 11396 18399 11398
rect 18423 11396 18479 11398
rect 18503 11396 18559 11398
rect 20735 14170 20791 14172
rect 20815 14170 20871 14172
rect 20895 14170 20951 14172
rect 20975 14170 21031 14172
rect 20735 14118 20781 14170
rect 20781 14118 20791 14170
rect 20815 14118 20845 14170
rect 20845 14118 20857 14170
rect 20857 14118 20871 14170
rect 20895 14118 20909 14170
rect 20909 14118 20921 14170
rect 20921 14118 20951 14170
rect 20975 14118 20985 14170
rect 20985 14118 21031 14170
rect 20735 14116 20791 14118
rect 20815 14116 20871 14118
rect 20895 14116 20951 14118
rect 20975 14116 21031 14118
rect 18263 10362 18319 10364
rect 18343 10362 18399 10364
rect 18423 10362 18479 10364
rect 18503 10362 18559 10364
rect 18263 10310 18309 10362
rect 18309 10310 18319 10362
rect 18343 10310 18373 10362
rect 18373 10310 18385 10362
rect 18385 10310 18399 10362
rect 18423 10310 18437 10362
rect 18437 10310 18449 10362
rect 18449 10310 18479 10362
rect 18503 10310 18513 10362
rect 18513 10310 18559 10362
rect 18263 10308 18319 10310
rect 18343 10308 18399 10310
rect 18423 10308 18479 10310
rect 18503 10308 18559 10310
rect 15790 7642 15846 7644
rect 15870 7642 15926 7644
rect 15950 7642 16006 7644
rect 16030 7642 16086 7644
rect 15790 7590 15836 7642
rect 15836 7590 15846 7642
rect 15870 7590 15900 7642
rect 15900 7590 15912 7642
rect 15912 7590 15926 7642
rect 15950 7590 15964 7642
rect 15964 7590 15976 7642
rect 15976 7590 16006 7642
rect 16030 7590 16040 7642
rect 16040 7590 16086 7642
rect 15790 7588 15846 7590
rect 15870 7588 15926 7590
rect 15950 7588 16006 7590
rect 16030 7588 16086 7590
rect 15790 6554 15846 6556
rect 15870 6554 15926 6556
rect 15950 6554 16006 6556
rect 16030 6554 16086 6556
rect 15790 6502 15836 6554
rect 15836 6502 15846 6554
rect 15870 6502 15900 6554
rect 15900 6502 15912 6554
rect 15912 6502 15926 6554
rect 15950 6502 15964 6554
rect 15964 6502 15976 6554
rect 15976 6502 16006 6554
rect 16030 6502 16040 6554
rect 16040 6502 16086 6554
rect 15790 6500 15846 6502
rect 15870 6500 15926 6502
rect 15950 6500 16006 6502
rect 16030 6500 16086 6502
rect 15790 5466 15846 5468
rect 15870 5466 15926 5468
rect 15950 5466 16006 5468
rect 16030 5466 16086 5468
rect 15790 5414 15836 5466
rect 15836 5414 15846 5466
rect 15870 5414 15900 5466
rect 15900 5414 15912 5466
rect 15912 5414 15926 5466
rect 15950 5414 15964 5466
rect 15964 5414 15976 5466
rect 15976 5414 16006 5466
rect 16030 5414 16040 5466
rect 16040 5414 16086 5466
rect 15790 5412 15846 5414
rect 15870 5412 15926 5414
rect 15950 5412 16006 5414
rect 16030 5412 16086 5414
rect 8373 4922 8429 4924
rect 8453 4922 8509 4924
rect 8533 4922 8589 4924
rect 8613 4922 8669 4924
rect 8373 4870 8419 4922
rect 8419 4870 8429 4922
rect 8453 4870 8483 4922
rect 8483 4870 8495 4922
rect 8495 4870 8509 4922
rect 8533 4870 8547 4922
rect 8547 4870 8559 4922
rect 8559 4870 8589 4922
rect 8613 4870 8623 4922
rect 8623 4870 8669 4922
rect 8373 4868 8429 4870
rect 8453 4868 8509 4870
rect 8533 4868 8589 4870
rect 8613 4868 8669 4870
rect 16486 5208 16542 5264
rect 8373 3834 8429 3836
rect 8453 3834 8509 3836
rect 8533 3834 8589 3836
rect 8613 3834 8669 3836
rect 8373 3782 8419 3834
rect 8419 3782 8429 3834
rect 8453 3782 8483 3834
rect 8483 3782 8495 3834
rect 8495 3782 8509 3834
rect 8533 3782 8547 3834
rect 8547 3782 8559 3834
rect 8559 3782 8589 3834
rect 8613 3782 8623 3834
rect 8623 3782 8669 3834
rect 8373 3780 8429 3782
rect 8453 3780 8509 3782
rect 8533 3780 8589 3782
rect 8613 3780 8669 3782
rect 10845 4378 10901 4380
rect 10925 4378 10981 4380
rect 11005 4378 11061 4380
rect 11085 4378 11141 4380
rect 10845 4326 10891 4378
rect 10891 4326 10901 4378
rect 10925 4326 10955 4378
rect 10955 4326 10967 4378
rect 10967 4326 10981 4378
rect 11005 4326 11019 4378
rect 11019 4326 11031 4378
rect 11031 4326 11061 4378
rect 11085 4326 11095 4378
rect 11095 4326 11141 4378
rect 10845 4324 10901 4326
rect 10925 4324 10981 4326
rect 11005 4324 11061 4326
rect 11085 4324 11141 4326
rect 10845 3290 10901 3292
rect 10925 3290 10981 3292
rect 11005 3290 11061 3292
rect 11085 3290 11141 3292
rect 10845 3238 10891 3290
rect 10891 3238 10901 3290
rect 10925 3238 10955 3290
rect 10955 3238 10967 3290
rect 10967 3238 10981 3290
rect 11005 3238 11019 3290
rect 11019 3238 11031 3290
rect 11031 3238 11061 3290
rect 11085 3238 11095 3290
rect 11095 3238 11141 3290
rect 10845 3236 10901 3238
rect 10925 3236 10981 3238
rect 11005 3236 11061 3238
rect 11085 3236 11141 3238
rect 8373 2746 8429 2748
rect 8453 2746 8509 2748
rect 8533 2746 8589 2748
rect 8613 2746 8669 2748
rect 8373 2694 8419 2746
rect 8419 2694 8429 2746
rect 8453 2694 8483 2746
rect 8483 2694 8495 2746
rect 8495 2694 8509 2746
rect 8533 2694 8547 2746
rect 8547 2694 8559 2746
rect 8559 2694 8589 2746
rect 8613 2694 8623 2746
rect 8623 2694 8669 2746
rect 8373 2692 8429 2694
rect 8453 2692 8509 2694
rect 8533 2692 8589 2694
rect 8613 2692 8669 2694
rect 13318 4922 13374 4924
rect 13398 4922 13454 4924
rect 13478 4922 13534 4924
rect 13558 4922 13614 4924
rect 13318 4870 13364 4922
rect 13364 4870 13374 4922
rect 13398 4870 13428 4922
rect 13428 4870 13440 4922
rect 13440 4870 13454 4922
rect 13478 4870 13492 4922
rect 13492 4870 13504 4922
rect 13504 4870 13534 4922
rect 13558 4870 13568 4922
rect 13568 4870 13614 4922
rect 13318 4868 13374 4870
rect 13398 4868 13454 4870
rect 13478 4868 13534 4870
rect 13558 4868 13614 4870
rect 13318 3834 13374 3836
rect 13398 3834 13454 3836
rect 13478 3834 13534 3836
rect 13558 3834 13614 3836
rect 13318 3782 13364 3834
rect 13364 3782 13374 3834
rect 13398 3782 13428 3834
rect 13428 3782 13440 3834
rect 13440 3782 13454 3834
rect 13478 3782 13492 3834
rect 13492 3782 13504 3834
rect 13504 3782 13534 3834
rect 13558 3782 13568 3834
rect 13568 3782 13614 3834
rect 13318 3780 13374 3782
rect 13398 3780 13454 3782
rect 13478 3780 13534 3782
rect 13558 3780 13614 3782
rect 13318 2746 13374 2748
rect 13398 2746 13454 2748
rect 13478 2746 13534 2748
rect 13558 2746 13614 2748
rect 13318 2694 13364 2746
rect 13364 2694 13374 2746
rect 13398 2694 13428 2746
rect 13428 2694 13440 2746
rect 13440 2694 13454 2746
rect 13478 2694 13492 2746
rect 13492 2694 13504 2746
rect 13504 2694 13534 2746
rect 13558 2694 13568 2746
rect 13568 2694 13614 2746
rect 13318 2692 13374 2694
rect 13398 2692 13454 2694
rect 13478 2692 13534 2694
rect 13558 2692 13614 2694
rect 15790 4378 15846 4380
rect 15870 4378 15926 4380
rect 15950 4378 16006 4380
rect 16030 4378 16086 4380
rect 15790 4326 15836 4378
rect 15836 4326 15846 4378
rect 15870 4326 15900 4378
rect 15900 4326 15912 4378
rect 15912 4326 15926 4378
rect 15950 4326 15964 4378
rect 15964 4326 15976 4378
rect 15976 4326 16006 4378
rect 16030 4326 16040 4378
rect 16040 4326 16086 4378
rect 15790 4324 15846 4326
rect 15870 4324 15926 4326
rect 15950 4324 16006 4326
rect 16030 4324 16086 4326
rect 20735 13082 20791 13084
rect 20815 13082 20871 13084
rect 20895 13082 20951 13084
rect 20975 13082 21031 13084
rect 20735 13030 20781 13082
rect 20781 13030 20791 13082
rect 20815 13030 20845 13082
rect 20845 13030 20857 13082
rect 20857 13030 20871 13082
rect 20895 13030 20909 13082
rect 20909 13030 20921 13082
rect 20921 13030 20951 13082
rect 20975 13030 20985 13082
rect 20985 13030 21031 13082
rect 20735 13028 20791 13030
rect 20815 13028 20871 13030
rect 20895 13028 20951 13030
rect 20975 13028 21031 13030
rect 18263 9274 18319 9276
rect 18343 9274 18399 9276
rect 18423 9274 18479 9276
rect 18503 9274 18559 9276
rect 18263 9222 18309 9274
rect 18309 9222 18319 9274
rect 18343 9222 18373 9274
rect 18373 9222 18385 9274
rect 18385 9222 18399 9274
rect 18423 9222 18437 9274
rect 18437 9222 18449 9274
rect 18449 9222 18479 9274
rect 18503 9222 18513 9274
rect 18513 9222 18559 9274
rect 18263 9220 18319 9222
rect 18343 9220 18399 9222
rect 18423 9220 18479 9222
rect 18503 9220 18559 9222
rect 20735 11994 20791 11996
rect 20815 11994 20871 11996
rect 20895 11994 20951 11996
rect 20975 11994 21031 11996
rect 20735 11942 20781 11994
rect 20781 11942 20791 11994
rect 20815 11942 20845 11994
rect 20845 11942 20857 11994
rect 20857 11942 20871 11994
rect 20895 11942 20909 11994
rect 20909 11942 20921 11994
rect 20921 11942 20951 11994
rect 20975 11942 20985 11994
rect 20985 11942 21031 11994
rect 20735 11940 20791 11942
rect 20815 11940 20871 11942
rect 20895 11940 20951 11942
rect 20975 11940 21031 11942
rect 20735 10906 20791 10908
rect 20815 10906 20871 10908
rect 20895 10906 20951 10908
rect 20975 10906 21031 10908
rect 20735 10854 20781 10906
rect 20781 10854 20791 10906
rect 20815 10854 20845 10906
rect 20845 10854 20857 10906
rect 20857 10854 20871 10906
rect 20895 10854 20909 10906
rect 20909 10854 20921 10906
rect 20921 10854 20951 10906
rect 20975 10854 20985 10906
rect 20985 10854 21031 10906
rect 20735 10852 20791 10854
rect 20815 10852 20871 10854
rect 20895 10852 20951 10854
rect 20975 10852 21031 10854
rect 20735 9818 20791 9820
rect 20815 9818 20871 9820
rect 20895 9818 20951 9820
rect 20975 9818 21031 9820
rect 20735 9766 20781 9818
rect 20781 9766 20791 9818
rect 20815 9766 20845 9818
rect 20845 9766 20857 9818
rect 20857 9766 20871 9818
rect 20895 9766 20909 9818
rect 20909 9766 20921 9818
rect 20921 9766 20951 9818
rect 20975 9766 20985 9818
rect 20985 9766 21031 9818
rect 20735 9764 20791 9766
rect 20815 9764 20871 9766
rect 20895 9764 20951 9766
rect 20975 9764 21031 9766
rect 18263 8186 18319 8188
rect 18343 8186 18399 8188
rect 18423 8186 18479 8188
rect 18503 8186 18559 8188
rect 18263 8134 18309 8186
rect 18309 8134 18319 8186
rect 18343 8134 18373 8186
rect 18373 8134 18385 8186
rect 18385 8134 18399 8186
rect 18423 8134 18437 8186
rect 18437 8134 18449 8186
rect 18449 8134 18479 8186
rect 18503 8134 18513 8186
rect 18513 8134 18559 8186
rect 18263 8132 18319 8134
rect 18343 8132 18399 8134
rect 18423 8132 18479 8134
rect 18503 8132 18559 8134
rect 20735 8730 20791 8732
rect 20815 8730 20871 8732
rect 20895 8730 20951 8732
rect 20975 8730 21031 8732
rect 20735 8678 20781 8730
rect 20781 8678 20791 8730
rect 20815 8678 20845 8730
rect 20845 8678 20857 8730
rect 20857 8678 20871 8730
rect 20895 8678 20909 8730
rect 20909 8678 20921 8730
rect 20921 8678 20951 8730
rect 20975 8678 20985 8730
rect 20985 8678 21031 8730
rect 20735 8676 20791 8678
rect 20815 8676 20871 8678
rect 20895 8676 20951 8678
rect 20975 8676 21031 8678
rect 18263 7098 18319 7100
rect 18343 7098 18399 7100
rect 18423 7098 18479 7100
rect 18503 7098 18559 7100
rect 18263 7046 18309 7098
rect 18309 7046 18319 7098
rect 18343 7046 18373 7098
rect 18373 7046 18385 7098
rect 18385 7046 18399 7098
rect 18423 7046 18437 7098
rect 18437 7046 18449 7098
rect 18449 7046 18479 7098
rect 18503 7046 18513 7098
rect 18513 7046 18559 7098
rect 18263 7044 18319 7046
rect 18343 7044 18399 7046
rect 18423 7044 18479 7046
rect 18503 7044 18559 7046
rect 17958 5072 18014 5128
rect 18263 6010 18319 6012
rect 18343 6010 18399 6012
rect 18423 6010 18479 6012
rect 18503 6010 18559 6012
rect 18263 5958 18309 6010
rect 18309 5958 18319 6010
rect 18343 5958 18373 6010
rect 18373 5958 18385 6010
rect 18385 5958 18399 6010
rect 18423 5958 18437 6010
rect 18437 5958 18449 6010
rect 18449 5958 18479 6010
rect 18503 5958 18513 6010
rect 18513 5958 18559 6010
rect 18263 5956 18319 5958
rect 18343 5956 18399 5958
rect 18423 5956 18479 5958
rect 18503 5956 18559 5958
rect 20735 7642 20791 7644
rect 20815 7642 20871 7644
rect 20895 7642 20951 7644
rect 20975 7642 21031 7644
rect 20735 7590 20781 7642
rect 20781 7590 20791 7642
rect 20815 7590 20845 7642
rect 20845 7590 20857 7642
rect 20857 7590 20871 7642
rect 20895 7590 20909 7642
rect 20909 7590 20921 7642
rect 20921 7590 20951 7642
rect 20975 7590 20985 7642
rect 20985 7590 21031 7642
rect 20735 7588 20791 7590
rect 20815 7588 20871 7590
rect 20895 7588 20951 7590
rect 20975 7588 21031 7590
rect 20735 6554 20791 6556
rect 20815 6554 20871 6556
rect 20895 6554 20951 6556
rect 20975 6554 21031 6556
rect 20735 6502 20781 6554
rect 20781 6502 20791 6554
rect 20815 6502 20845 6554
rect 20845 6502 20857 6554
rect 20857 6502 20871 6554
rect 20895 6502 20909 6554
rect 20909 6502 20921 6554
rect 20921 6502 20951 6554
rect 20975 6502 20985 6554
rect 20985 6502 21031 6554
rect 20735 6500 20791 6502
rect 20815 6500 20871 6502
rect 20895 6500 20951 6502
rect 20975 6500 21031 6502
rect 18263 4922 18319 4924
rect 18343 4922 18399 4924
rect 18423 4922 18479 4924
rect 18503 4922 18559 4924
rect 18263 4870 18309 4922
rect 18309 4870 18319 4922
rect 18343 4870 18373 4922
rect 18373 4870 18385 4922
rect 18385 4870 18399 4922
rect 18423 4870 18437 4922
rect 18437 4870 18449 4922
rect 18449 4870 18479 4922
rect 18503 4870 18513 4922
rect 18513 4870 18559 4922
rect 18263 4868 18319 4870
rect 18343 4868 18399 4870
rect 18423 4868 18479 4870
rect 18503 4868 18559 4870
rect 20735 5466 20791 5468
rect 20815 5466 20871 5468
rect 20895 5466 20951 5468
rect 20975 5466 21031 5468
rect 20735 5414 20781 5466
rect 20781 5414 20791 5466
rect 20815 5414 20845 5466
rect 20845 5414 20857 5466
rect 20857 5414 20871 5466
rect 20895 5414 20909 5466
rect 20909 5414 20921 5466
rect 20921 5414 20951 5466
rect 20975 5414 20985 5466
rect 20985 5414 21031 5466
rect 20735 5412 20791 5414
rect 20815 5412 20871 5414
rect 20895 5412 20951 5414
rect 20975 5412 21031 5414
rect 15790 3290 15846 3292
rect 15870 3290 15926 3292
rect 15950 3290 16006 3292
rect 16030 3290 16086 3292
rect 15790 3238 15836 3290
rect 15836 3238 15846 3290
rect 15870 3238 15900 3290
rect 15900 3238 15912 3290
rect 15912 3238 15926 3290
rect 15950 3238 15964 3290
rect 15964 3238 15976 3290
rect 15976 3238 16006 3290
rect 16030 3238 16040 3290
rect 16040 3238 16086 3290
rect 15790 3236 15846 3238
rect 15870 3236 15926 3238
rect 15950 3236 16006 3238
rect 16030 3236 16086 3238
rect 20735 4378 20791 4380
rect 20815 4378 20871 4380
rect 20895 4378 20951 4380
rect 20975 4378 21031 4380
rect 20735 4326 20781 4378
rect 20781 4326 20791 4378
rect 20815 4326 20845 4378
rect 20845 4326 20857 4378
rect 20857 4326 20871 4378
rect 20895 4326 20909 4378
rect 20909 4326 20921 4378
rect 20921 4326 20951 4378
rect 20975 4326 20985 4378
rect 20985 4326 21031 4378
rect 20735 4324 20791 4326
rect 20815 4324 20871 4326
rect 20895 4324 20951 4326
rect 20975 4324 21031 4326
rect 18263 3834 18319 3836
rect 18343 3834 18399 3836
rect 18423 3834 18479 3836
rect 18503 3834 18559 3836
rect 18263 3782 18309 3834
rect 18309 3782 18319 3834
rect 18343 3782 18373 3834
rect 18373 3782 18385 3834
rect 18385 3782 18399 3834
rect 18423 3782 18437 3834
rect 18437 3782 18449 3834
rect 18449 3782 18479 3834
rect 18503 3782 18513 3834
rect 18513 3782 18559 3834
rect 18263 3780 18319 3782
rect 18343 3780 18399 3782
rect 18423 3780 18479 3782
rect 18503 3780 18559 3782
rect 20735 3290 20791 3292
rect 20815 3290 20871 3292
rect 20895 3290 20951 3292
rect 20975 3290 21031 3292
rect 20735 3238 20781 3290
rect 20781 3238 20791 3290
rect 20815 3238 20845 3290
rect 20845 3238 20857 3290
rect 20857 3238 20871 3290
rect 20895 3238 20909 3290
rect 20909 3238 20921 3290
rect 20921 3238 20951 3290
rect 20975 3238 20985 3290
rect 20985 3238 21031 3290
rect 20735 3236 20791 3238
rect 20815 3236 20871 3238
rect 20895 3236 20951 3238
rect 20975 3236 21031 3238
rect 18263 2746 18319 2748
rect 18343 2746 18399 2748
rect 18423 2746 18479 2748
rect 18503 2746 18559 2748
rect 18263 2694 18309 2746
rect 18309 2694 18319 2746
rect 18343 2694 18373 2746
rect 18373 2694 18385 2746
rect 18385 2694 18399 2746
rect 18423 2694 18437 2746
rect 18437 2694 18449 2746
rect 18449 2694 18479 2746
rect 18503 2694 18513 2746
rect 18513 2694 18559 2746
rect 18263 2692 18319 2694
rect 18343 2692 18399 2694
rect 18423 2692 18479 2694
rect 18503 2692 18559 2694
rect 5900 2202 5956 2204
rect 5980 2202 6036 2204
rect 6060 2202 6116 2204
rect 6140 2202 6196 2204
rect 5900 2150 5946 2202
rect 5946 2150 5956 2202
rect 5980 2150 6010 2202
rect 6010 2150 6022 2202
rect 6022 2150 6036 2202
rect 6060 2150 6074 2202
rect 6074 2150 6086 2202
rect 6086 2150 6116 2202
rect 6140 2150 6150 2202
rect 6150 2150 6196 2202
rect 5900 2148 5956 2150
rect 5980 2148 6036 2150
rect 6060 2148 6116 2150
rect 6140 2148 6196 2150
rect 10845 2202 10901 2204
rect 10925 2202 10981 2204
rect 11005 2202 11061 2204
rect 11085 2202 11141 2204
rect 10845 2150 10891 2202
rect 10891 2150 10901 2202
rect 10925 2150 10955 2202
rect 10955 2150 10967 2202
rect 10967 2150 10981 2202
rect 11005 2150 11019 2202
rect 11019 2150 11031 2202
rect 11031 2150 11061 2202
rect 11085 2150 11095 2202
rect 11095 2150 11141 2202
rect 10845 2148 10901 2150
rect 10925 2148 10981 2150
rect 11005 2148 11061 2150
rect 11085 2148 11141 2150
rect 15790 2202 15846 2204
rect 15870 2202 15926 2204
rect 15950 2202 16006 2204
rect 16030 2202 16086 2204
rect 15790 2150 15836 2202
rect 15836 2150 15846 2202
rect 15870 2150 15900 2202
rect 15900 2150 15912 2202
rect 15912 2150 15926 2202
rect 15950 2150 15964 2202
rect 15964 2150 15976 2202
rect 15976 2150 16006 2202
rect 16030 2150 16040 2202
rect 16040 2150 16086 2202
rect 15790 2148 15846 2150
rect 15870 2148 15926 2150
rect 15950 2148 16006 2150
rect 16030 2148 16086 2150
rect 20735 2202 20791 2204
rect 20815 2202 20871 2204
rect 20895 2202 20951 2204
rect 20975 2202 21031 2204
rect 20735 2150 20781 2202
rect 20781 2150 20791 2202
rect 20815 2150 20845 2202
rect 20845 2150 20857 2202
rect 20857 2150 20871 2202
rect 20895 2150 20909 2202
rect 20909 2150 20921 2202
rect 20921 2150 20951 2202
rect 20975 2150 20985 2202
rect 20985 2150 21031 2202
rect 20735 2148 20791 2150
rect 20815 2148 20871 2150
rect 20895 2148 20951 2150
rect 20975 2148 21031 2150
<< metal3 >>
rect 5890 19616 6206 19617
rect 5890 19552 5896 19616
rect 5960 19552 5976 19616
rect 6040 19552 6056 19616
rect 6120 19552 6136 19616
rect 6200 19552 6206 19616
rect 5890 19551 6206 19552
rect 10835 19616 11151 19617
rect 10835 19552 10841 19616
rect 10905 19552 10921 19616
rect 10985 19552 11001 19616
rect 11065 19552 11081 19616
rect 11145 19552 11151 19616
rect 10835 19551 11151 19552
rect 15780 19616 16096 19617
rect 15780 19552 15786 19616
rect 15850 19552 15866 19616
rect 15930 19552 15946 19616
rect 16010 19552 16026 19616
rect 16090 19552 16096 19616
rect 15780 19551 16096 19552
rect 20725 19616 21041 19617
rect 20725 19552 20731 19616
rect 20795 19552 20811 19616
rect 20875 19552 20891 19616
rect 20955 19552 20971 19616
rect 21035 19552 21041 19616
rect 20725 19551 21041 19552
rect 3418 19072 3734 19073
rect 3418 19008 3424 19072
rect 3488 19008 3504 19072
rect 3568 19008 3584 19072
rect 3648 19008 3664 19072
rect 3728 19008 3734 19072
rect 3418 19007 3734 19008
rect 8363 19072 8679 19073
rect 8363 19008 8369 19072
rect 8433 19008 8449 19072
rect 8513 19008 8529 19072
rect 8593 19008 8609 19072
rect 8673 19008 8679 19072
rect 8363 19007 8679 19008
rect 13308 19072 13624 19073
rect 13308 19008 13314 19072
rect 13378 19008 13394 19072
rect 13458 19008 13474 19072
rect 13538 19008 13554 19072
rect 13618 19008 13624 19072
rect 13308 19007 13624 19008
rect 18253 19072 18569 19073
rect 18253 19008 18259 19072
rect 18323 19008 18339 19072
rect 18403 19008 18419 19072
rect 18483 19008 18499 19072
rect 18563 19008 18569 19072
rect 18253 19007 18569 19008
rect 5890 18528 6206 18529
rect 5890 18464 5896 18528
rect 5960 18464 5976 18528
rect 6040 18464 6056 18528
rect 6120 18464 6136 18528
rect 6200 18464 6206 18528
rect 5890 18463 6206 18464
rect 10835 18528 11151 18529
rect 10835 18464 10841 18528
rect 10905 18464 10921 18528
rect 10985 18464 11001 18528
rect 11065 18464 11081 18528
rect 11145 18464 11151 18528
rect 10835 18463 11151 18464
rect 15780 18528 16096 18529
rect 15780 18464 15786 18528
rect 15850 18464 15866 18528
rect 15930 18464 15946 18528
rect 16010 18464 16026 18528
rect 16090 18464 16096 18528
rect 15780 18463 16096 18464
rect 20725 18528 21041 18529
rect 20725 18464 20731 18528
rect 20795 18464 20811 18528
rect 20875 18464 20891 18528
rect 20955 18464 20971 18528
rect 21035 18464 21041 18528
rect 20725 18463 21041 18464
rect 0 18322 800 18352
rect 1853 18322 1919 18325
rect 0 18320 1919 18322
rect 0 18264 1858 18320
rect 1914 18264 1919 18320
rect 0 18262 1919 18264
rect 0 18232 800 18262
rect 1853 18259 1919 18262
rect 3418 17984 3734 17985
rect 3418 17920 3424 17984
rect 3488 17920 3504 17984
rect 3568 17920 3584 17984
rect 3648 17920 3664 17984
rect 3728 17920 3734 17984
rect 3418 17919 3734 17920
rect 8363 17984 8679 17985
rect 8363 17920 8369 17984
rect 8433 17920 8449 17984
rect 8513 17920 8529 17984
rect 8593 17920 8609 17984
rect 8673 17920 8679 17984
rect 8363 17919 8679 17920
rect 13308 17984 13624 17985
rect 13308 17920 13314 17984
rect 13378 17920 13394 17984
rect 13458 17920 13474 17984
rect 13538 17920 13554 17984
rect 13618 17920 13624 17984
rect 13308 17919 13624 17920
rect 18253 17984 18569 17985
rect 18253 17920 18259 17984
rect 18323 17920 18339 17984
rect 18403 17920 18419 17984
rect 18483 17920 18499 17984
rect 18563 17920 18569 17984
rect 18253 17919 18569 17920
rect 5890 17440 6206 17441
rect 5890 17376 5896 17440
rect 5960 17376 5976 17440
rect 6040 17376 6056 17440
rect 6120 17376 6136 17440
rect 6200 17376 6206 17440
rect 5890 17375 6206 17376
rect 10835 17440 11151 17441
rect 10835 17376 10841 17440
rect 10905 17376 10921 17440
rect 10985 17376 11001 17440
rect 11065 17376 11081 17440
rect 11145 17376 11151 17440
rect 10835 17375 11151 17376
rect 15780 17440 16096 17441
rect 15780 17376 15786 17440
rect 15850 17376 15866 17440
rect 15930 17376 15946 17440
rect 16010 17376 16026 17440
rect 16090 17376 16096 17440
rect 15780 17375 16096 17376
rect 20725 17440 21041 17441
rect 20725 17376 20731 17440
rect 20795 17376 20811 17440
rect 20875 17376 20891 17440
rect 20955 17376 20971 17440
rect 21035 17376 21041 17440
rect 20725 17375 21041 17376
rect 3418 16896 3734 16897
rect 3418 16832 3424 16896
rect 3488 16832 3504 16896
rect 3568 16832 3584 16896
rect 3648 16832 3664 16896
rect 3728 16832 3734 16896
rect 3418 16831 3734 16832
rect 8363 16896 8679 16897
rect 8363 16832 8369 16896
rect 8433 16832 8449 16896
rect 8513 16832 8529 16896
rect 8593 16832 8609 16896
rect 8673 16832 8679 16896
rect 8363 16831 8679 16832
rect 13308 16896 13624 16897
rect 13308 16832 13314 16896
rect 13378 16832 13394 16896
rect 13458 16832 13474 16896
rect 13538 16832 13554 16896
rect 13618 16832 13624 16896
rect 13308 16831 13624 16832
rect 18253 16896 18569 16897
rect 18253 16832 18259 16896
rect 18323 16832 18339 16896
rect 18403 16832 18419 16896
rect 18483 16832 18499 16896
rect 18563 16832 18569 16896
rect 18253 16831 18569 16832
rect 5890 16352 6206 16353
rect 5890 16288 5896 16352
rect 5960 16288 5976 16352
rect 6040 16288 6056 16352
rect 6120 16288 6136 16352
rect 6200 16288 6206 16352
rect 5890 16287 6206 16288
rect 10835 16352 11151 16353
rect 10835 16288 10841 16352
rect 10905 16288 10921 16352
rect 10985 16288 11001 16352
rect 11065 16288 11081 16352
rect 11145 16288 11151 16352
rect 10835 16287 11151 16288
rect 15780 16352 16096 16353
rect 15780 16288 15786 16352
rect 15850 16288 15866 16352
rect 15930 16288 15946 16352
rect 16010 16288 16026 16352
rect 16090 16288 16096 16352
rect 15780 16287 16096 16288
rect 20725 16352 21041 16353
rect 20725 16288 20731 16352
rect 20795 16288 20811 16352
rect 20875 16288 20891 16352
rect 20955 16288 20971 16352
rect 21035 16288 21041 16352
rect 20725 16287 21041 16288
rect 3418 15808 3734 15809
rect 3418 15744 3424 15808
rect 3488 15744 3504 15808
rect 3568 15744 3584 15808
rect 3648 15744 3664 15808
rect 3728 15744 3734 15808
rect 3418 15743 3734 15744
rect 8363 15808 8679 15809
rect 8363 15744 8369 15808
rect 8433 15744 8449 15808
rect 8513 15744 8529 15808
rect 8593 15744 8609 15808
rect 8673 15744 8679 15808
rect 8363 15743 8679 15744
rect 13308 15808 13624 15809
rect 13308 15744 13314 15808
rect 13378 15744 13394 15808
rect 13458 15744 13474 15808
rect 13538 15744 13554 15808
rect 13618 15744 13624 15808
rect 13308 15743 13624 15744
rect 18253 15808 18569 15809
rect 18253 15744 18259 15808
rect 18323 15744 18339 15808
rect 18403 15744 18419 15808
rect 18483 15744 18499 15808
rect 18563 15744 18569 15808
rect 18253 15743 18569 15744
rect 5890 15264 6206 15265
rect 5890 15200 5896 15264
rect 5960 15200 5976 15264
rect 6040 15200 6056 15264
rect 6120 15200 6136 15264
rect 6200 15200 6206 15264
rect 5890 15199 6206 15200
rect 10835 15264 11151 15265
rect 10835 15200 10841 15264
rect 10905 15200 10921 15264
rect 10985 15200 11001 15264
rect 11065 15200 11081 15264
rect 11145 15200 11151 15264
rect 10835 15199 11151 15200
rect 15780 15264 16096 15265
rect 15780 15200 15786 15264
rect 15850 15200 15866 15264
rect 15930 15200 15946 15264
rect 16010 15200 16026 15264
rect 16090 15200 16096 15264
rect 15780 15199 16096 15200
rect 20725 15264 21041 15265
rect 20725 15200 20731 15264
rect 20795 15200 20811 15264
rect 20875 15200 20891 15264
rect 20955 15200 20971 15264
rect 21035 15200 21041 15264
rect 20725 15199 21041 15200
rect 3418 14720 3734 14721
rect 3418 14656 3424 14720
rect 3488 14656 3504 14720
rect 3568 14656 3584 14720
rect 3648 14656 3664 14720
rect 3728 14656 3734 14720
rect 3418 14655 3734 14656
rect 8363 14720 8679 14721
rect 8363 14656 8369 14720
rect 8433 14656 8449 14720
rect 8513 14656 8529 14720
rect 8593 14656 8609 14720
rect 8673 14656 8679 14720
rect 8363 14655 8679 14656
rect 13308 14720 13624 14721
rect 13308 14656 13314 14720
rect 13378 14656 13394 14720
rect 13458 14656 13474 14720
rect 13538 14656 13554 14720
rect 13618 14656 13624 14720
rect 13308 14655 13624 14656
rect 18253 14720 18569 14721
rect 18253 14656 18259 14720
rect 18323 14656 18339 14720
rect 18403 14656 18419 14720
rect 18483 14656 18499 14720
rect 18563 14656 18569 14720
rect 18253 14655 18569 14656
rect 13353 14378 13419 14381
rect 17861 14378 17927 14381
rect 18229 14378 18295 14381
rect 13353 14376 18295 14378
rect 13353 14320 13358 14376
rect 13414 14320 17866 14376
rect 17922 14320 18234 14376
rect 18290 14320 18295 14376
rect 13353 14318 18295 14320
rect 13353 14315 13419 14318
rect 17861 14315 17927 14318
rect 18229 14315 18295 14318
rect 5890 14176 6206 14177
rect 5890 14112 5896 14176
rect 5960 14112 5976 14176
rect 6040 14112 6056 14176
rect 6120 14112 6136 14176
rect 6200 14112 6206 14176
rect 5890 14111 6206 14112
rect 10835 14176 11151 14177
rect 10835 14112 10841 14176
rect 10905 14112 10921 14176
rect 10985 14112 11001 14176
rect 11065 14112 11081 14176
rect 11145 14112 11151 14176
rect 10835 14111 11151 14112
rect 15780 14176 16096 14177
rect 15780 14112 15786 14176
rect 15850 14112 15866 14176
rect 15930 14112 15946 14176
rect 16010 14112 16026 14176
rect 16090 14112 16096 14176
rect 15780 14111 16096 14112
rect 20725 14176 21041 14177
rect 20725 14112 20731 14176
rect 20795 14112 20811 14176
rect 20875 14112 20891 14176
rect 20955 14112 20971 14176
rect 21035 14112 21041 14176
rect 20725 14111 21041 14112
rect 15285 14106 15351 14109
rect 15285 14104 15394 14106
rect 15285 14048 15290 14104
rect 15346 14048 15394 14104
rect 15285 14043 15394 14048
rect 15334 13834 15394 14043
rect 15653 13834 15719 13837
rect 15334 13832 15719 13834
rect 15334 13776 15658 13832
rect 15714 13776 15719 13832
rect 15334 13774 15719 13776
rect 15653 13771 15719 13774
rect 3418 13632 3734 13633
rect 3418 13568 3424 13632
rect 3488 13568 3504 13632
rect 3568 13568 3584 13632
rect 3648 13568 3664 13632
rect 3728 13568 3734 13632
rect 3418 13567 3734 13568
rect 8363 13632 8679 13633
rect 8363 13568 8369 13632
rect 8433 13568 8449 13632
rect 8513 13568 8529 13632
rect 8593 13568 8609 13632
rect 8673 13568 8679 13632
rect 8363 13567 8679 13568
rect 13308 13632 13624 13633
rect 13308 13568 13314 13632
rect 13378 13568 13394 13632
rect 13458 13568 13474 13632
rect 13538 13568 13554 13632
rect 13618 13568 13624 13632
rect 13308 13567 13624 13568
rect 18253 13632 18569 13633
rect 18253 13568 18259 13632
rect 18323 13568 18339 13632
rect 18403 13568 18419 13632
rect 18483 13568 18499 13632
rect 18563 13568 18569 13632
rect 18253 13567 18569 13568
rect 5890 13088 6206 13089
rect 5890 13024 5896 13088
rect 5960 13024 5976 13088
rect 6040 13024 6056 13088
rect 6120 13024 6136 13088
rect 6200 13024 6206 13088
rect 5890 13023 6206 13024
rect 10835 13088 11151 13089
rect 10835 13024 10841 13088
rect 10905 13024 10921 13088
rect 10985 13024 11001 13088
rect 11065 13024 11081 13088
rect 11145 13024 11151 13088
rect 10835 13023 11151 13024
rect 15780 13088 16096 13089
rect 15780 13024 15786 13088
rect 15850 13024 15866 13088
rect 15930 13024 15946 13088
rect 16010 13024 16026 13088
rect 16090 13024 16096 13088
rect 15780 13023 16096 13024
rect 20725 13088 21041 13089
rect 20725 13024 20731 13088
rect 20795 13024 20811 13088
rect 20875 13024 20891 13088
rect 20955 13024 20971 13088
rect 21035 13024 21041 13088
rect 20725 13023 21041 13024
rect 3418 12544 3734 12545
rect 3418 12480 3424 12544
rect 3488 12480 3504 12544
rect 3568 12480 3584 12544
rect 3648 12480 3664 12544
rect 3728 12480 3734 12544
rect 3418 12479 3734 12480
rect 8363 12544 8679 12545
rect 8363 12480 8369 12544
rect 8433 12480 8449 12544
rect 8513 12480 8529 12544
rect 8593 12480 8609 12544
rect 8673 12480 8679 12544
rect 8363 12479 8679 12480
rect 13308 12544 13624 12545
rect 13308 12480 13314 12544
rect 13378 12480 13394 12544
rect 13458 12480 13474 12544
rect 13538 12480 13554 12544
rect 13618 12480 13624 12544
rect 13308 12479 13624 12480
rect 18253 12544 18569 12545
rect 18253 12480 18259 12544
rect 18323 12480 18339 12544
rect 18403 12480 18419 12544
rect 18483 12480 18499 12544
rect 18563 12480 18569 12544
rect 18253 12479 18569 12480
rect 13445 12338 13511 12341
rect 16573 12338 16639 12341
rect 13445 12336 16639 12338
rect 13445 12280 13450 12336
rect 13506 12280 16578 12336
rect 16634 12280 16639 12336
rect 13445 12278 16639 12280
rect 13445 12275 13511 12278
rect 16573 12275 16639 12278
rect 9673 12202 9739 12205
rect 19425 12202 19491 12205
rect 9673 12200 19491 12202
rect 9673 12144 9678 12200
rect 9734 12144 19430 12200
rect 19486 12144 19491 12200
rect 9673 12142 19491 12144
rect 9673 12139 9739 12142
rect 19425 12139 19491 12142
rect 5890 12000 6206 12001
rect 5890 11936 5896 12000
rect 5960 11936 5976 12000
rect 6040 11936 6056 12000
rect 6120 11936 6136 12000
rect 6200 11936 6206 12000
rect 5890 11935 6206 11936
rect 10835 12000 11151 12001
rect 10835 11936 10841 12000
rect 10905 11936 10921 12000
rect 10985 11936 11001 12000
rect 11065 11936 11081 12000
rect 11145 11936 11151 12000
rect 10835 11935 11151 11936
rect 15780 12000 16096 12001
rect 15780 11936 15786 12000
rect 15850 11936 15866 12000
rect 15930 11936 15946 12000
rect 16010 11936 16026 12000
rect 16090 11936 16096 12000
rect 15780 11935 16096 11936
rect 20725 12000 21041 12001
rect 20725 11936 20731 12000
rect 20795 11936 20811 12000
rect 20875 11936 20891 12000
rect 20955 11936 20971 12000
rect 21035 11936 21041 12000
rect 20725 11935 21041 11936
rect 3418 11456 3734 11457
rect 3418 11392 3424 11456
rect 3488 11392 3504 11456
rect 3568 11392 3584 11456
rect 3648 11392 3664 11456
rect 3728 11392 3734 11456
rect 3418 11391 3734 11392
rect 8363 11456 8679 11457
rect 8363 11392 8369 11456
rect 8433 11392 8449 11456
rect 8513 11392 8529 11456
rect 8593 11392 8609 11456
rect 8673 11392 8679 11456
rect 8363 11391 8679 11392
rect 13308 11456 13624 11457
rect 13308 11392 13314 11456
rect 13378 11392 13394 11456
rect 13458 11392 13474 11456
rect 13538 11392 13554 11456
rect 13618 11392 13624 11456
rect 13308 11391 13624 11392
rect 18253 11456 18569 11457
rect 18253 11392 18259 11456
rect 18323 11392 18339 11456
rect 18403 11392 18419 11456
rect 18483 11392 18499 11456
rect 18563 11392 18569 11456
rect 18253 11391 18569 11392
rect 0 10978 800 11008
rect 1669 10978 1735 10981
rect 0 10976 1735 10978
rect 0 10920 1674 10976
rect 1730 10920 1735 10976
rect 0 10918 1735 10920
rect 0 10888 800 10918
rect 1669 10915 1735 10918
rect 5890 10912 6206 10913
rect 5890 10848 5896 10912
rect 5960 10848 5976 10912
rect 6040 10848 6056 10912
rect 6120 10848 6136 10912
rect 6200 10848 6206 10912
rect 5890 10847 6206 10848
rect 10835 10912 11151 10913
rect 10835 10848 10841 10912
rect 10905 10848 10921 10912
rect 10985 10848 11001 10912
rect 11065 10848 11081 10912
rect 11145 10848 11151 10912
rect 10835 10847 11151 10848
rect 15780 10912 16096 10913
rect 15780 10848 15786 10912
rect 15850 10848 15866 10912
rect 15930 10848 15946 10912
rect 16010 10848 16026 10912
rect 16090 10848 16096 10912
rect 15780 10847 16096 10848
rect 20725 10912 21041 10913
rect 20725 10848 20731 10912
rect 20795 10848 20811 10912
rect 20875 10848 20891 10912
rect 20955 10848 20971 10912
rect 21035 10848 21041 10912
rect 20725 10847 21041 10848
rect 3418 10368 3734 10369
rect 3418 10304 3424 10368
rect 3488 10304 3504 10368
rect 3568 10304 3584 10368
rect 3648 10304 3664 10368
rect 3728 10304 3734 10368
rect 3418 10303 3734 10304
rect 8363 10368 8679 10369
rect 8363 10304 8369 10368
rect 8433 10304 8449 10368
rect 8513 10304 8529 10368
rect 8593 10304 8609 10368
rect 8673 10304 8679 10368
rect 8363 10303 8679 10304
rect 13308 10368 13624 10369
rect 13308 10304 13314 10368
rect 13378 10304 13394 10368
rect 13458 10304 13474 10368
rect 13538 10304 13554 10368
rect 13618 10304 13624 10368
rect 13308 10303 13624 10304
rect 18253 10368 18569 10369
rect 18253 10304 18259 10368
rect 18323 10304 18339 10368
rect 18403 10304 18419 10368
rect 18483 10304 18499 10368
rect 18563 10304 18569 10368
rect 18253 10303 18569 10304
rect 5890 9824 6206 9825
rect 5890 9760 5896 9824
rect 5960 9760 5976 9824
rect 6040 9760 6056 9824
rect 6120 9760 6136 9824
rect 6200 9760 6206 9824
rect 5890 9759 6206 9760
rect 10835 9824 11151 9825
rect 10835 9760 10841 9824
rect 10905 9760 10921 9824
rect 10985 9760 11001 9824
rect 11065 9760 11081 9824
rect 11145 9760 11151 9824
rect 10835 9759 11151 9760
rect 15780 9824 16096 9825
rect 15780 9760 15786 9824
rect 15850 9760 15866 9824
rect 15930 9760 15946 9824
rect 16010 9760 16026 9824
rect 16090 9760 16096 9824
rect 15780 9759 16096 9760
rect 20725 9824 21041 9825
rect 20725 9760 20731 9824
rect 20795 9760 20811 9824
rect 20875 9760 20891 9824
rect 20955 9760 20971 9824
rect 21035 9760 21041 9824
rect 20725 9759 21041 9760
rect 3418 9280 3734 9281
rect 3418 9216 3424 9280
rect 3488 9216 3504 9280
rect 3568 9216 3584 9280
rect 3648 9216 3664 9280
rect 3728 9216 3734 9280
rect 3418 9215 3734 9216
rect 8363 9280 8679 9281
rect 8363 9216 8369 9280
rect 8433 9216 8449 9280
rect 8513 9216 8529 9280
rect 8593 9216 8609 9280
rect 8673 9216 8679 9280
rect 8363 9215 8679 9216
rect 13308 9280 13624 9281
rect 13308 9216 13314 9280
rect 13378 9216 13394 9280
rect 13458 9216 13474 9280
rect 13538 9216 13554 9280
rect 13618 9216 13624 9280
rect 13308 9215 13624 9216
rect 18253 9280 18569 9281
rect 18253 9216 18259 9280
rect 18323 9216 18339 9280
rect 18403 9216 18419 9280
rect 18483 9216 18499 9280
rect 18563 9216 18569 9280
rect 18253 9215 18569 9216
rect 5890 8736 6206 8737
rect 5890 8672 5896 8736
rect 5960 8672 5976 8736
rect 6040 8672 6056 8736
rect 6120 8672 6136 8736
rect 6200 8672 6206 8736
rect 5890 8671 6206 8672
rect 10835 8736 11151 8737
rect 10835 8672 10841 8736
rect 10905 8672 10921 8736
rect 10985 8672 11001 8736
rect 11065 8672 11081 8736
rect 11145 8672 11151 8736
rect 10835 8671 11151 8672
rect 15780 8736 16096 8737
rect 15780 8672 15786 8736
rect 15850 8672 15866 8736
rect 15930 8672 15946 8736
rect 16010 8672 16026 8736
rect 16090 8672 16096 8736
rect 15780 8671 16096 8672
rect 20725 8736 21041 8737
rect 20725 8672 20731 8736
rect 20795 8672 20811 8736
rect 20875 8672 20891 8736
rect 20955 8672 20971 8736
rect 21035 8672 21041 8736
rect 20725 8671 21041 8672
rect 3418 8192 3734 8193
rect 3418 8128 3424 8192
rect 3488 8128 3504 8192
rect 3568 8128 3584 8192
rect 3648 8128 3664 8192
rect 3728 8128 3734 8192
rect 3418 8127 3734 8128
rect 8363 8192 8679 8193
rect 8363 8128 8369 8192
rect 8433 8128 8449 8192
rect 8513 8128 8529 8192
rect 8593 8128 8609 8192
rect 8673 8128 8679 8192
rect 8363 8127 8679 8128
rect 13308 8192 13624 8193
rect 13308 8128 13314 8192
rect 13378 8128 13394 8192
rect 13458 8128 13474 8192
rect 13538 8128 13554 8192
rect 13618 8128 13624 8192
rect 13308 8127 13624 8128
rect 18253 8192 18569 8193
rect 18253 8128 18259 8192
rect 18323 8128 18339 8192
rect 18403 8128 18419 8192
rect 18483 8128 18499 8192
rect 18563 8128 18569 8192
rect 18253 8127 18569 8128
rect 5890 7648 6206 7649
rect 5890 7584 5896 7648
rect 5960 7584 5976 7648
rect 6040 7584 6056 7648
rect 6120 7584 6136 7648
rect 6200 7584 6206 7648
rect 5890 7583 6206 7584
rect 10835 7648 11151 7649
rect 10835 7584 10841 7648
rect 10905 7584 10921 7648
rect 10985 7584 11001 7648
rect 11065 7584 11081 7648
rect 11145 7584 11151 7648
rect 10835 7583 11151 7584
rect 15780 7648 16096 7649
rect 15780 7584 15786 7648
rect 15850 7584 15866 7648
rect 15930 7584 15946 7648
rect 16010 7584 16026 7648
rect 16090 7584 16096 7648
rect 15780 7583 16096 7584
rect 20725 7648 21041 7649
rect 20725 7584 20731 7648
rect 20795 7584 20811 7648
rect 20875 7584 20891 7648
rect 20955 7584 20971 7648
rect 21035 7584 21041 7648
rect 20725 7583 21041 7584
rect 3418 7104 3734 7105
rect 3418 7040 3424 7104
rect 3488 7040 3504 7104
rect 3568 7040 3584 7104
rect 3648 7040 3664 7104
rect 3728 7040 3734 7104
rect 3418 7039 3734 7040
rect 8363 7104 8679 7105
rect 8363 7040 8369 7104
rect 8433 7040 8449 7104
rect 8513 7040 8529 7104
rect 8593 7040 8609 7104
rect 8673 7040 8679 7104
rect 8363 7039 8679 7040
rect 13308 7104 13624 7105
rect 13308 7040 13314 7104
rect 13378 7040 13394 7104
rect 13458 7040 13474 7104
rect 13538 7040 13554 7104
rect 13618 7040 13624 7104
rect 13308 7039 13624 7040
rect 18253 7104 18569 7105
rect 18253 7040 18259 7104
rect 18323 7040 18339 7104
rect 18403 7040 18419 7104
rect 18483 7040 18499 7104
rect 18563 7040 18569 7104
rect 18253 7039 18569 7040
rect 5890 6560 6206 6561
rect 5890 6496 5896 6560
rect 5960 6496 5976 6560
rect 6040 6496 6056 6560
rect 6120 6496 6136 6560
rect 6200 6496 6206 6560
rect 5890 6495 6206 6496
rect 10835 6560 11151 6561
rect 10835 6496 10841 6560
rect 10905 6496 10921 6560
rect 10985 6496 11001 6560
rect 11065 6496 11081 6560
rect 11145 6496 11151 6560
rect 10835 6495 11151 6496
rect 15780 6560 16096 6561
rect 15780 6496 15786 6560
rect 15850 6496 15866 6560
rect 15930 6496 15946 6560
rect 16010 6496 16026 6560
rect 16090 6496 16096 6560
rect 15780 6495 16096 6496
rect 20725 6560 21041 6561
rect 20725 6496 20731 6560
rect 20795 6496 20811 6560
rect 20875 6496 20891 6560
rect 20955 6496 20971 6560
rect 21035 6496 21041 6560
rect 20725 6495 21041 6496
rect 3418 6016 3734 6017
rect 3418 5952 3424 6016
rect 3488 5952 3504 6016
rect 3568 5952 3584 6016
rect 3648 5952 3664 6016
rect 3728 5952 3734 6016
rect 3418 5951 3734 5952
rect 8363 6016 8679 6017
rect 8363 5952 8369 6016
rect 8433 5952 8449 6016
rect 8513 5952 8529 6016
rect 8593 5952 8609 6016
rect 8673 5952 8679 6016
rect 8363 5951 8679 5952
rect 13308 6016 13624 6017
rect 13308 5952 13314 6016
rect 13378 5952 13394 6016
rect 13458 5952 13474 6016
rect 13538 5952 13554 6016
rect 13618 5952 13624 6016
rect 13308 5951 13624 5952
rect 18253 6016 18569 6017
rect 18253 5952 18259 6016
rect 18323 5952 18339 6016
rect 18403 5952 18419 6016
rect 18483 5952 18499 6016
rect 18563 5952 18569 6016
rect 18253 5951 18569 5952
rect 5890 5472 6206 5473
rect 5890 5408 5896 5472
rect 5960 5408 5976 5472
rect 6040 5408 6056 5472
rect 6120 5408 6136 5472
rect 6200 5408 6206 5472
rect 5890 5407 6206 5408
rect 10835 5472 11151 5473
rect 10835 5408 10841 5472
rect 10905 5408 10921 5472
rect 10985 5408 11001 5472
rect 11065 5408 11081 5472
rect 11145 5408 11151 5472
rect 10835 5407 11151 5408
rect 15780 5472 16096 5473
rect 15780 5408 15786 5472
rect 15850 5408 15866 5472
rect 15930 5408 15946 5472
rect 16010 5408 16026 5472
rect 16090 5408 16096 5472
rect 15780 5407 16096 5408
rect 20725 5472 21041 5473
rect 20725 5408 20731 5472
rect 20795 5408 20811 5472
rect 20875 5408 20891 5472
rect 20955 5408 20971 5472
rect 21035 5408 21041 5472
rect 20725 5407 21041 5408
rect 11145 5266 11211 5269
rect 16481 5266 16547 5269
rect 11145 5264 16547 5266
rect 11145 5208 11150 5264
rect 11206 5208 16486 5264
rect 16542 5208 16547 5264
rect 11145 5206 16547 5208
rect 11145 5203 11211 5206
rect 16481 5203 16547 5206
rect 2773 5130 2839 5133
rect 2957 5130 3023 5133
rect 17953 5130 18019 5133
rect 2773 5128 18019 5130
rect 2773 5072 2778 5128
rect 2834 5072 2962 5128
rect 3018 5072 17958 5128
rect 18014 5072 18019 5128
rect 2773 5070 18019 5072
rect 2773 5067 2839 5070
rect 2957 5067 3023 5070
rect 17953 5067 18019 5070
rect 3418 4928 3734 4929
rect 3418 4864 3424 4928
rect 3488 4864 3504 4928
rect 3568 4864 3584 4928
rect 3648 4864 3664 4928
rect 3728 4864 3734 4928
rect 3418 4863 3734 4864
rect 8363 4928 8679 4929
rect 8363 4864 8369 4928
rect 8433 4864 8449 4928
rect 8513 4864 8529 4928
rect 8593 4864 8609 4928
rect 8673 4864 8679 4928
rect 8363 4863 8679 4864
rect 13308 4928 13624 4929
rect 13308 4864 13314 4928
rect 13378 4864 13394 4928
rect 13458 4864 13474 4928
rect 13538 4864 13554 4928
rect 13618 4864 13624 4928
rect 13308 4863 13624 4864
rect 18253 4928 18569 4929
rect 18253 4864 18259 4928
rect 18323 4864 18339 4928
rect 18403 4864 18419 4928
rect 18483 4864 18499 4928
rect 18563 4864 18569 4928
rect 18253 4863 18569 4864
rect 5890 4384 6206 4385
rect 5890 4320 5896 4384
rect 5960 4320 5976 4384
rect 6040 4320 6056 4384
rect 6120 4320 6136 4384
rect 6200 4320 6206 4384
rect 5890 4319 6206 4320
rect 10835 4384 11151 4385
rect 10835 4320 10841 4384
rect 10905 4320 10921 4384
rect 10985 4320 11001 4384
rect 11065 4320 11081 4384
rect 11145 4320 11151 4384
rect 10835 4319 11151 4320
rect 15780 4384 16096 4385
rect 15780 4320 15786 4384
rect 15850 4320 15866 4384
rect 15930 4320 15946 4384
rect 16010 4320 16026 4384
rect 16090 4320 16096 4384
rect 15780 4319 16096 4320
rect 20725 4384 21041 4385
rect 20725 4320 20731 4384
rect 20795 4320 20811 4384
rect 20875 4320 20891 4384
rect 20955 4320 20971 4384
rect 21035 4320 21041 4384
rect 20725 4319 21041 4320
rect 3418 3840 3734 3841
rect 3418 3776 3424 3840
rect 3488 3776 3504 3840
rect 3568 3776 3584 3840
rect 3648 3776 3664 3840
rect 3728 3776 3734 3840
rect 3418 3775 3734 3776
rect 8363 3840 8679 3841
rect 8363 3776 8369 3840
rect 8433 3776 8449 3840
rect 8513 3776 8529 3840
rect 8593 3776 8609 3840
rect 8673 3776 8679 3840
rect 8363 3775 8679 3776
rect 13308 3840 13624 3841
rect 13308 3776 13314 3840
rect 13378 3776 13394 3840
rect 13458 3776 13474 3840
rect 13538 3776 13554 3840
rect 13618 3776 13624 3840
rect 13308 3775 13624 3776
rect 18253 3840 18569 3841
rect 18253 3776 18259 3840
rect 18323 3776 18339 3840
rect 18403 3776 18419 3840
rect 18483 3776 18499 3840
rect 18563 3776 18569 3840
rect 18253 3775 18569 3776
rect 0 3634 800 3664
rect 3141 3634 3207 3637
rect 0 3632 3207 3634
rect 0 3576 3146 3632
rect 3202 3576 3207 3632
rect 0 3574 3207 3576
rect 0 3544 800 3574
rect 3141 3571 3207 3574
rect 5890 3296 6206 3297
rect 5890 3232 5896 3296
rect 5960 3232 5976 3296
rect 6040 3232 6056 3296
rect 6120 3232 6136 3296
rect 6200 3232 6206 3296
rect 5890 3231 6206 3232
rect 10835 3296 11151 3297
rect 10835 3232 10841 3296
rect 10905 3232 10921 3296
rect 10985 3232 11001 3296
rect 11065 3232 11081 3296
rect 11145 3232 11151 3296
rect 10835 3231 11151 3232
rect 15780 3296 16096 3297
rect 15780 3232 15786 3296
rect 15850 3232 15866 3296
rect 15930 3232 15946 3296
rect 16010 3232 16026 3296
rect 16090 3232 16096 3296
rect 15780 3231 16096 3232
rect 20725 3296 21041 3297
rect 20725 3232 20731 3296
rect 20795 3232 20811 3296
rect 20875 3232 20891 3296
rect 20955 3232 20971 3296
rect 21035 3232 21041 3296
rect 20725 3231 21041 3232
rect 3418 2752 3734 2753
rect 3418 2688 3424 2752
rect 3488 2688 3504 2752
rect 3568 2688 3584 2752
rect 3648 2688 3664 2752
rect 3728 2688 3734 2752
rect 3418 2687 3734 2688
rect 8363 2752 8679 2753
rect 8363 2688 8369 2752
rect 8433 2688 8449 2752
rect 8513 2688 8529 2752
rect 8593 2688 8609 2752
rect 8673 2688 8679 2752
rect 8363 2687 8679 2688
rect 13308 2752 13624 2753
rect 13308 2688 13314 2752
rect 13378 2688 13394 2752
rect 13458 2688 13474 2752
rect 13538 2688 13554 2752
rect 13618 2688 13624 2752
rect 13308 2687 13624 2688
rect 18253 2752 18569 2753
rect 18253 2688 18259 2752
rect 18323 2688 18339 2752
rect 18403 2688 18419 2752
rect 18483 2688 18499 2752
rect 18563 2688 18569 2752
rect 18253 2687 18569 2688
rect 5890 2208 6206 2209
rect 5890 2144 5896 2208
rect 5960 2144 5976 2208
rect 6040 2144 6056 2208
rect 6120 2144 6136 2208
rect 6200 2144 6206 2208
rect 5890 2143 6206 2144
rect 10835 2208 11151 2209
rect 10835 2144 10841 2208
rect 10905 2144 10921 2208
rect 10985 2144 11001 2208
rect 11065 2144 11081 2208
rect 11145 2144 11151 2208
rect 10835 2143 11151 2144
rect 15780 2208 16096 2209
rect 15780 2144 15786 2208
rect 15850 2144 15866 2208
rect 15930 2144 15946 2208
rect 16010 2144 16026 2208
rect 16090 2144 16096 2208
rect 15780 2143 16096 2144
rect 20725 2208 21041 2209
rect 20725 2144 20731 2208
rect 20795 2144 20811 2208
rect 20875 2144 20891 2208
rect 20955 2144 20971 2208
rect 21035 2144 21041 2208
rect 20725 2143 21041 2144
<< via3 >>
rect 5896 19612 5960 19616
rect 5896 19556 5900 19612
rect 5900 19556 5956 19612
rect 5956 19556 5960 19612
rect 5896 19552 5960 19556
rect 5976 19612 6040 19616
rect 5976 19556 5980 19612
rect 5980 19556 6036 19612
rect 6036 19556 6040 19612
rect 5976 19552 6040 19556
rect 6056 19612 6120 19616
rect 6056 19556 6060 19612
rect 6060 19556 6116 19612
rect 6116 19556 6120 19612
rect 6056 19552 6120 19556
rect 6136 19612 6200 19616
rect 6136 19556 6140 19612
rect 6140 19556 6196 19612
rect 6196 19556 6200 19612
rect 6136 19552 6200 19556
rect 10841 19612 10905 19616
rect 10841 19556 10845 19612
rect 10845 19556 10901 19612
rect 10901 19556 10905 19612
rect 10841 19552 10905 19556
rect 10921 19612 10985 19616
rect 10921 19556 10925 19612
rect 10925 19556 10981 19612
rect 10981 19556 10985 19612
rect 10921 19552 10985 19556
rect 11001 19612 11065 19616
rect 11001 19556 11005 19612
rect 11005 19556 11061 19612
rect 11061 19556 11065 19612
rect 11001 19552 11065 19556
rect 11081 19612 11145 19616
rect 11081 19556 11085 19612
rect 11085 19556 11141 19612
rect 11141 19556 11145 19612
rect 11081 19552 11145 19556
rect 15786 19612 15850 19616
rect 15786 19556 15790 19612
rect 15790 19556 15846 19612
rect 15846 19556 15850 19612
rect 15786 19552 15850 19556
rect 15866 19612 15930 19616
rect 15866 19556 15870 19612
rect 15870 19556 15926 19612
rect 15926 19556 15930 19612
rect 15866 19552 15930 19556
rect 15946 19612 16010 19616
rect 15946 19556 15950 19612
rect 15950 19556 16006 19612
rect 16006 19556 16010 19612
rect 15946 19552 16010 19556
rect 16026 19612 16090 19616
rect 16026 19556 16030 19612
rect 16030 19556 16086 19612
rect 16086 19556 16090 19612
rect 16026 19552 16090 19556
rect 20731 19612 20795 19616
rect 20731 19556 20735 19612
rect 20735 19556 20791 19612
rect 20791 19556 20795 19612
rect 20731 19552 20795 19556
rect 20811 19612 20875 19616
rect 20811 19556 20815 19612
rect 20815 19556 20871 19612
rect 20871 19556 20875 19612
rect 20811 19552 20875 19556
rect 20891 19612 20955 19616
rect 20891 19556 20895 19612
rect 20895 19556 20951 19612
rect 20951 19556 20955 19612
rect 20891 19552 20955 19556
rect 20971 19612 21035 19616
rect 20971 19556 20975 19612
rect 20975 19556 21031 19612
rect 21031 19556 21035 19612
rect 20971 19552 21035 19556
rect 3424 19068 3488 19072
rect 3424 19012 3428 19068
rect 3428 19012 3484 19068
rect 3484 19012 3488 19068
rect 3424 19008 3488 19012
rect 3504 19068 3568 19072
rect 3504 19012 3508 19068
rect 3508 19012 3564 19068
rect 3564 19012 3568 19068
rect 3504 19008 3568 19012
rect 3584 19068 3648 19072
rect 3584 19012 3588 19068
rect 3588 19012 3644 19068
rect 3644 19012 3648 19068
rect 3584 19008 3648 19012
rect 3664 19068 3728 19072
rect 3664 19012 3668 19068
rect 3668 19012 3724 19068
rect 3724 19012 3728 19068
rect 3664 19008 3728 19012
rect 8369 19068 8433 19072
rect 8369 19012 8373 19068
rect 8373 19012 8429 19068
rect 8429 19012 8433 19068
rect 8369 19008 8433 19012
rect 8449 19068 8513 19072
rect 8449 19012 8453 19068
rect 8453 19012 8509 19068
rect 8509 19012 8513 19068
rect 8449 19008 8513 19012
rect 8529 19068 8593 19072
rect 8529 19012 8533 19068
rect 8533 19012 8589 19068
rect 8589 19012 8593 19068
rect 8529 19008 8593 19012
rect 8609 19068 8673 19072
rect 8609 19012 8613 19068
rect 8613 19012 8669 19068
rect 8669 19012 8673 19068
rect 8609 19008 8673 19012
rect 13314 19068 13378 19072
rect 13314 19012 13318 19068
rect 13318 19012 13374 19068
rect 13374 19012 13378 19068
rect 13314 19008 13378 19012
rect 13394 19068 13458 19072
rect 13394 19012 13398 19068
rect 13398 19012 13454 19068
rect 13454 19012 13458 19068
rect 13394 19008 13458 19012
rect 13474 19068 13538 19072
rect 13474 19012 13478 19068
rect 13478 19012 13534 19068
rect 13534 19012 13538 19068
rect 13474 19008 13538 19012
rect 13554 19068 13618 19072
rect 13554 19012 13558 19068
rect 13558 19012 13614 19068
rect 13614 19012 13618 19068
rect 13554 19008 13618 19012
rect 18259 19068 18323 19072
rect 18259 19012 18263 19068
rect 18263 19012 18319 19068
rect 18319 19012 18323 19068
rect 18259 19008 18323 19012
rect 18339 19068 18403 19072
rect 18339 19012 18343 19068
rect 18343 19012 18399 19068
rect 18399 19012 18403 19068
rect 18339 19008 18403 19012
rect 18419 19068 18483 19072
rect 18419 19012 18423 19068
rect 18423 19012 18479 19068
rect 18479 19012 18483 19068
rect 18419 19008 18483 19012
rect 18499 19068 18563 19072
rect 18499 19012 18503 19068
rect 18503 19012 18559 19068
rect 18559 19012 18563 19068
rect 18499 19008 18563 19012
rect 5896 18524 5960 18528
rect 5896 18468 5900 18524
rect 5900 18468 5956 18524
rect 5956 18468 5960 18524
rect 5896 18464 5960 18468
rect 5976 18524 6040 18528
rect 5976 18468 5980 18524
rect 5980 18468 6036 18524
rect 6036 18468 6040 18524
rect 5976 18464 6040 18468
rect 6056 18524 6120 18528
rect 6056 18468 6060 18524
rect 6060 18468 6116 18524
rect 6116 18468 6120 18524
rect 6056 18464 6120 18468
rect 6136 18524 6200 18528
rect 6136 18468 6140 18524
rect 6140 18468 6196 18524
rect 6196 18468 6200 18524
rect 6136 18464 6200 18468
rect 10841 18524 10905 18528
rect 10841 18468 10845 18524
rect 10845 18468 10901 18524
rect 10901 18468 10905 18524
rect 10841 18464 10905 18468
rect 10921 18524 10985 18528
rect 10921 18468 10925 18524
rect 10925 18468 10981 18524
rect 10981 18468 10985 18524
rect 10921 18464 10985 18468
rect 11001 18524 11065 18528
rect 11001 18468 11005 18524
rect 11005 18468 11061 18524
rect 11061 18468 11065 18524
rect 11001 18464 11065 18468
rect 11081 18524 11145 18528
rect 11081 18468 11085 18524
rect 11085 18468 11141 18524
rect 11141 18468 11145 18524
rect 11081 18464 11145 18468
rect 15786 18524 15850 18528
rect 15786 18468 15790 18524
rect 15790 18468 15846 18524
rect 15846 18468 15850 18524
rect 15786 18464 15850 18468
rect 15866 18524 15930 18528
rect 15866 18468 15870 18524
rect 15870 18468 15926 18524
rect 15926 18468 15930 18524
rect 15866 18464 15930 18468
rect 15946 18524 16010 18528
rect 15946 18468 15950 18524
rect 15950 18468 16006 18524
rect 16006 18468 16010 18524
rect 15946 18464 16010 18468
rect 16026 18524 16090 18528
rect 16026 18468 16030 18524
rect 16030 18468 16086 18524
rect 16086 18468 16090 18524
rect 16026 18464 16090 18468
rect 20731 18524 20795 18528
rect 20731 18468 20735 18524
rect 20735 18468 20791 18524
rect 20791 18468 20795 18524
rect 20731 18464 20795 18468
rect 20811 18524 20875 18528
rect 20811 18468 20815 18524
rect 20815 18468 20871 18524
rect 20871 18468 20875 18524
rect 20811 18464 20875 18468
rect 20891 18524 20955 18528
rect 20891 18468 20895 18524
rect 20895 18468 20951 18524
rect 20951 18468 20955 18524
rect 20891 18464 20955 18468
rect 20971 18524 21035 18528
rect 20971 18468 20975 18524
rect 20975 18468 21031 18524
rect 21031 18468 21035 18524
rect 20971 18464 21035 18468
rect 3424 17980 3488 17984
rect 3424 17924 3428 17980
rect 3428 17924 3484 17980
rect 3484 17924 3488 17980
rect 3424 17920 3488 17924
rect 3504 17980 3568 17984
rect 3504 17924 3508 17980
rect 3508 17924 3564 17980
rect 3564 17924 3568 17980
rect 3504 17920 3568 17924
rect 3584 17980 3648 17984
rect 3584 17924 3588 17980
rect 3588 17924 3644 17980
rect 3644 17924 3648 17980
rect 3584 17920 3648 17924
rect 3664 17980 3728 17984
rect 3664 17924 3668 17980
rect 3668 17924 3724 17980
rect 3724 17924 3728 17980
rect 3664 17920 3728 17924
rect 8369 17980 8433 17984
rect 8369 17924 8373 17980
rect 8373 17924 8429 17980
rect 8429 17924 8433 17980
rect 8369 17920 8433 17924
rect 8449 17980 8513 17984
rect 8449 17924 8453 17980
rect 8453 17924 8509 17980
rect 8509 17924 8513 17980
rect 8449 17920 8513 17924
rect 8529 17980 8593 17984
rect 8529 17924 8533 17980
rect 8533 17924 8589 17980
rect 8589 17924 8593 17980
rect 8529 17920 8593 17924
rect 8609 17980 8673 17984
rect 8609 17924 8613 17980
rect 8613 17924 8669 17980
rect 8669 17924 8673 17980
rect 8609 17920 8673 17924
rect 13314 17980 13378 17984
rect 13314 17924 13318 17980
rect 13318 17924 13374 17980
rect 13374 17924 13378 17980
rect 13314 17920 13378 17924
rect 13394 17980 13458 17984
rect 13394 17924 13398 17980
rect 13398 17924 13454 17980
rect 13454 17924 13458 17980
rect 13394 17920 13458 17924
rect 13474 17980 13538 17984
rect 13474 17924 13478 17980
rect 13478 17924 13534 17980
rect 13534 17924 13538 17980
rect 13474 17920 13538 17924
rect 13554 17980 13618 17984
rect 13554 17924 13558 17980
rect 13558 17924 13614 17980
rect 13614 17924 13618 17980
rect 13554 17920 13618 17924
rect 18259 17980 18323 17984
rect 18259 17924 18263 17980
rect 18263 17924 18319 17980
rect 18319 17924 18323 17980
rect 18259 17920 18323 17924
rect 18339 17980 18403 17984
rect 18339 17924 18343 17980
rect 18343 17924 18399 17980
rect 18399 17924 18403 17980
rect 18339 17920 18403 17924
rect 18419 17980 18483 17984
rect 18419 17924 18423 17980
rect 18423 17924 18479 17980
rect 18479 17924 18483 17980
rect 18419 17920 18483 17924
rect 18499 17980 18563 17984
rect 18499 17924 18503 17980
rect 18503 17924 18559 17980
rect 18559 17924 18563 17980
rect 18499 17920 18563 17924
rect 5896 17436 5960 17440
rect 5896 17380 5900 17436
rect 5900 17380 5956 17436
rect 5956 17380 5960 17436
rect 5896 17376 5960 17380
rect 5976 17436 6040 17440
rect 5976 17380 5980 17436
rect 5980 17380 6036 17436
rect 6036 17380 6040 17436
rect 5976 17376 6040 17380
rect 6056 17436 6120 17440
rect 6056 17380 6060 17436
rect 6060 17380 6116 17436
rect 6116 17380 6120 17436
rect 6056 17376 6120 17380
rect 6136 17436 6200 17440
rect 6136 17380 6140 17436
rect 6140 17380 6196 17436
rect 6196 17380 6200 17436
rect 6136 17376 6200 17380
rect 10841 17436 10905 17440
rect 10841 17380 10845 17436
rect 10845 17380 10901 17436
rect 10901 17380 10905 17436
rect 10841 17376 10905 17380
rect 10921 17436 10985 17440
rect 10921 17380 10925 17436
rect 10925 17380 10981 17436
rect 10981 17380 10985 17436
rect 10921 17376 10985 17380
rect 11001 17436 11065 17440
rect 11001 17380 11005 17436
rect 11005 17380 11061 17436
rect 11061 17380 11065 17436
rect 11001 17376 11065 17380
rect 11081 17436 11145 17440
rect 11081 17380 11085 17436
rect 11085 17380 11141 17436
rect 11141 17380 11145 17436
rect 11081 17376 11145 17380
rect 15786 17436 15850 17440
rect 15786 17380 15790 17436
rect 15790 17380 15846 17436
rect 15846 17380 15850 17436
rect 15786 17376 15850 17380
rect 15866 17436 15930 17440
rect 15866 17380 15870 17436
rect 15870 17380 15926 17436
rect 15926 17380 15930 17436
rect 15866 17376 15930 17380
rect 15946 17436 16010 17440
rect 15946 17380 15950 17436
rect 15950 17380 16006 17436
rect 16006 17380 16010 17436
rect 15946 17376 16010 17380
rect 16026 17436 16090 17440
rect 16026 17380 16030 17436
rect 16030 17380 16086 17436
rect 16086 17380 16090 17436
rect 16026 17376 16090 17380
rect 20731 17436 20795 17440
rect 20731 17380 20735 17436
rect 20735 17380 20791 17436
rect 20791 17380 20795 17436
rect 20731 17376 20795 17380
rect 20811 17436 20875 17440
rect 20811 17380 20815 17436
rect 20815 17380 20871 17436
rect 20871 17380 20875 17436
rect 20811 17376 20875 17380
rect 20891 17436 20955 17440
rect 20891 17380 20895 17436
rect 20895 17380 20951 17436
rect 20951 17380 20955 17436
rect 20891 17376 20955 17380
rect 20971 17436 21035 17440
rect 20971 17380 20975 17436
rect 20975 17380 21031 17436
rect 21031 17380 21035 17436
rect 20971 17376 21035 17380
rect 3424 16892 3488 16896
rect 3424 16836 3428 16892
rect 3428 16836 3484 16892
rect 3484 16836 3488 16892
rect 3424 16832 3488 16836
rect 3504 16892 3568 16896
rect 3504 16836 3508 16892
rect 3508 16836 3564 16892
rect 3564 16836 3568 16892
rect 3504 16832 3568 16836
rect 3584 16892 3648 16896
rect 3584 16836 3588 16892
rect 3588 16836 3644 16892
rect 3644 16836 3648 16892
rect 3584 16832 3648 16836
rect 3664 16892 3728 16896
rect 3664 16836 3668 16892
rect 3668 16836 3724 16892
rect 3724 16836 3728 16892
rect 3664 16832 3728 16836
rect 8369 16892 8433 16896
rect 8369 16836 8373 16892
rect 8373 16836 8429 16892
rect 8429 16836 8433 16892
rect 8369 16832 8433 16836
rect 8449 16892 8513 16896
rect 8449 16836 8453 16892
rect 8453 16836 8509 16892
rect 8509 16836 8513 16892
rect 8449 16832 8513 16836
rect 8529 16892 8593 16896
rect 8529 16836 8533 16892
rect 8533 16836 8589 16892
rect 8589 16836 8593 16892
rect 8529 16832 8593 16836
rect 8609 16892 8673 16896
rect 8609 16836 8613 16892
rect 8613 16836 8669 16892
rect 8669 16836 8673 16892
rect 8609 16832 8673 16836
rect 13314 16892 13378 16896
rect 13314 16836 13318 16892
rect 13318 16836 13374 16892
rect 13374 16836 13378 16892
rect 13314 16832 13378 16836
rect 13394 16892 13458 16896
rect 13394 16836 13398 16892
rect 13398 16836 13454 16892
rect 13454 16836 13458 16892
rect 13394 16832 13458 16836
rect 13474 16892 13538 16896
rect 13474 16836 13478 16892
rect 13478 16836 13534 16892
rect 13534 16836 13538 16892
rect 13474 16832 13538 16836
rect 13554 16892 13618 16896
rect 13554 16836 13558 16892
rect 13558 16836 13614 16892
rect 13614 16836 13618 16892
rect 13554 16832 13618 16836
rect 18259 16892 18323 16896
rect 18259 16836 18263 16892
rect 18263 16836 18319 16892
rect 18319 16836 18323 16892
rect 18259 16832 18323 16836
rect 18339 16892 18403 16896
rect 18339 16836 18343 16892
rect 18343 16836 18399 16892
rect 18399 16836 18403 16892
rect 18339 16832 18403 16836
rect 18419 16892 18483 16896
rect 18419 16836 18423 16892
rect 18423 16836 18479 16892
rect 18479 16836 18483 16892
rect 18419 16832 18483 16836
rect 18499 16892 18563 16896
rect 18499 16836 18503 16892
rect 18503 16836 18559 16892
rect 18559 16836 18563 16892
rect 18499 16832 18563 16836
rect 5896 16348 5960 16352
rect 5896 16292 5900 16348
rect 5900 16292 5956 16348
rect 5956 16292 5960 16348
rect 5896 16288 5960 16292
rect 5976 16348 6040 16352
rect 5976 16292 5980 16348
rect 5980 16292 6036 16348
rect 6036 16292 6040 16348
rect 5976 16288 6040 16292
rect 6056 16348 6120 16352
rect 6056 16292 6060 16348
rect 6060 16292 6116 16348
rect 6116 16292 6120 16348
rect 6056 16288 6120 16292
rect 6136 16348 6200 16352
rect 6136 16292 6140 16348
rect 6140 16292 6196 16348
rect 6196 16292 6200 16348
rect 6136 16288 6200 16292
rect 10841 16348 10905 16352
rect 10841 16292 10845 16348
rect 10845 16292 10901 16348
rect 10901 16292 10905 16348
rect 10841 16288 10905 16292
rect 10921 16348 10985 16352
rect 10921 16292 10925 16348
rect 10925 16292 10981 16348
rect 10981 16292 10985 16348
rect 10921 16288 10985 16292
rect 11001 16348 11065 16352
rect 11001 16292 11005 16348
rect 11005 16292 11061 16348
rect 11061 16292 11065 16348
rect 11001 16288 11065 16292
rect 11081 16348 11145 16352
rect 11081 16292 11085 16348
rect 11085 16292 11141 16348
rect 11141 16292 11145 16348
rect 11081 16288 11145 16292
rect 15786 16348 15850 16352
rect 15786 16292 15790 16348
rect 15790 16292 15846 16348
rect 15846 16292 15850 16348
rect 15786 16288 15850 16292
rect 15866 16348 15930 16352
rect 15866 16292 15870 16348
rect 15870 16292 15926 16348
rect 15926 16292 15930 16348
rect 15866 16288 15930 16292
rect 15946 16348 16010 16352
rect 15946 16292 15950 16348
rect 15950 16292 16006 16348
rect 16006 16292 16010 16348
rect 15946 16288 16010 16292
rect 16026 16348 16090 16352
rect 16026 16292 16030 16348
rect 16030 16292 16086 16348
rect 16086 16292 16090 16348
rect 16026 16288 16090 16292
rect 20731 16348 20795 16352
rect 20731 16292 20735 16348
rect 20735 16292 20791 16348
rect 20791 16292 20795 16348
rect 20731 16288 20795 16292
rect 20811 16348 20875 16352
rect 20811 16292 20815 16348
rect 20815 16292 20871 16348
rect 20871 16292 20875 16348
rect 20811 16288 20875 16292
rect 20891 16348 20955 16352
rect 20891 16292 20895 16348
rect 20895 16292 20951 16348
rect 20951 16292 20955 16348
rect 20891 16288 20955 16292
rect 20971 16348 21035 16352
rect 20971 16292 20975 16348
rect 20975 16292 21031 16348
rect 21031 16292 21035 16348
rect 20971 16288 21035 16292
rect 3424 15804 3488 15808
rect 3424 15748 3428 15804
rect 3428 15748 3484 15804
rect 3484 15748 3488 15804
rect 3424 15744 3488 15748
rect 3504 15804 3568 15808
rect 3504 15748 3508 15804
rect 3508 15748 3564 15804
rect 3564 15748 3568 15804
rect 3504 15744 3568 15748
rect 3584 15804 3648 15808
rect 3584 15748 3588 15804
rect 3588 15748 3644 15804
rect 3644 15748 3648 15804
rect 3584 15744 3648 15748
rect 3664 15804 3728 15808
rect 3664 15748 3668 15804
rect 3668 15748 3724 15804
rect 3724 15748 3728 15804
rect 3664 15744 3728 15748
rect 8369 15804 8433 15808
rect 8369 15748 8373 15804
rect 8373 15748 8429 15804
rect 8429 15748 8433 15804
rect 8369 15744 8433 15748
rect 8449 15804 8513 15808
rect 8449 15748 8453 15804
rect 8453 15748 8509 15804
rect 8509 15748 8513 15804
rect 8449 15744 8513 15748
rect 8529 15804 8593 15808
rect 8529 15748 8533 15804
rect 8533 15748 8589 15804
rect 8589 15748 8593 15804
rect 8529 15744 8593 15748
rect 8609 15804 8673 15808
rect 8609 15748 8613 15804
rect 8613 15748 8669 15804
rect 8669 15748 8673 15804
rect 8609 15744 8673 15748
rect 13314 15804 13378 15808
rect 13314 15748 13318 15804
rect 13318 15748 13374 15804
rect 13374 15748 13378 15804
rect 13314 15744 13378 15748
rect 13394 15804 13458 15808
rect 13394 15748 13398 15804
rect 13398 15748 13454 15804
rect 13454 15748 13458 15804
rect 13394 15744 13458 15748
rect 13474 15804 13538 15808
rect 13474 15748 13478 15804
rect 13478 15748 13534 15804
rect 13534 15748 13538 15804
rect 13474 15744 13538 15748
rect 13554 15804 13618 15808
rect 13554 15748 13558 15804
rect 13558 15748 13614 15804
rect 13614 15748 13618 15804
rect 13554 15744 13618 15748
rect 18259 15804 18323 15808
rect 18259 15748 18263 15804
rect 18263 15748 18319 15804
rect 18319 15748 18323 15804
rect 18259 15744 18323 15748
rect 18339 15804 18403 15808
rect 18339 15748 18343 15804
rect 18343 15748 18399 15804
rect 18399 15748 18403 15804
rect 18339 15744 18403 15748
rect 18419 15804 18483 15808
rect 18419 15748 18423 15804
rect 18423 15748 18479 15804
rect 18479 15748 18483 15804
rect 18419 15744 18483 15748
rect 18499 15804 18563 15808
rect 18499 15748 18503 15804
rect 18503 15748 18559 15804
rect 18559 15748 18563 15804
rect 18499 15744 18563 15748
rect 5896 15260 5960 15264
rect 5896 15204 5900 15260
rect 5900 15204 5956 15260
rect 5956 15204 5960 15260
rect 5896 15200 5960 15204
rect 5976 15260 6040 15264
rect 5976 15204 5980 15260
rect 5980 15204 6036 15260
rect 6036 15204 6040 15260
rect 5976 15200 6040 15204
rect 6056 15260 6120 15264
rect 6056 15204 6060 15260
rect 6060 15204 6116 15260
rect 6116 15204 6120 15260
rect 6056 15200 6120 15204
rect 6136 15260 6200 15264
rect 6136 15204 6140 15260
rect 6140 15204 6196 15260
rect 6196 15204 6200 15260
rect 6136 15200 6200 15204
rect 10841 15260 10905 15264
rect 10841 15204 10845 15260
rect 10845 15204 10901 15260
rect 10901 15204 10905 15260
rect 10841 15200 10905 15204
rect 10921 15260 10985 15264
rect 10921 15204 10925 15260
rect 10925 15204 10981 15260
rect 10981 15204 10985 15260
rect 10921 15200 10985 15204
rect 11001 15260 11065 15264
rect 11001 15204 11005 15260
rect 11005 15204 11061 15260
rect 11061 15204 11065 15260
rect 11001 15200 11065 15204
rect 11081 15260 11145 15264
rect 11081 15204 11085 15260
rect 11085 15204 11141 15260
rect 11141 15204 11145 15260
rect 11081 15200 11145 15204
rect 15786 15260 15850 15264
rect 15786 15204 15790 15260
rect 15790 15204 15846 15260
rect 15846 15204 15850 15260
rect 15786 15200 15850 15204
rect 15866 15260 15930 15264
rect 15866 15204 15870 15260
rect 15870 15204 15926 15260
rect 15926 15204 15930 15260
rect 15866 15200 15930 15204
rect 15946 15260 16010 15264
rect 15946 15204 15950 15260
rect 15950 15204 16006 15260
rect 16006 15204 16010 15260
rect 15946 15200 16010 15204
rect 16026 15260 16090 15264
rect 16026 15204 16030 15260
rect 16030 15204 16086 15260
rect 16086 15204 16090 15260
rect 16026 15200 16090 15204
rect 20731 15260 20795 15264
rect 20731 15204 20735 15260
rect 20735 15204 20791 15260
rect 20791 15204 20795 15260
rect 20731 15200 20795 15204
rect 20811 15260 20875 15264
rect 20811 15204 20815 15260
rect 20815 15204 20871 15260
rect 20871 15204 20875 15260
rect 20811 15200 20875 15204
rect 20891 15260 20955 15264
rect 20891 15204 20895 15260
rect 20895 15204 20951 15260
rect 20951 15204 20955 15260
rect 20891 15200 20955 15204
rect 20971 15260 21035 15264
rect 20971 15204 20975 15260
rect 20975 15204 21031 15260
rect 21031 15204 21035 15260
rect 20971 15200 21035 15204
rect 3424 14716 3488 14720
rect 3424 14660 3428 14716
rect 3428 14660 3484 14716
rect 3484 14660 3488 14716
rect 3424 14656 3488 14660
rect 3504 14716 3568 14720
rect 3504 14660 3508 14716
rect 3508 14660 3564 14716
rect 3564 14660 3568 14716
rect 3504 14656 3568 14660
rect 3584 14716 3648 14720
rect 3584 14660 3588 14716
rect 3588 14660 3644 14716
rect 3644 14660 3648 14716
rect 3584 14656 3648 14660
rect 3664 14716 3728 14720
rect 3664 14660 3668 14716
rect 3668 14660 3724 14716
rect 3724 14660 3728 14716
rect 3664 14656 3728 14660
rect 8369 14716 8433 14720
rect 8369 14660 8373 14716
rect 8373 14660 8429 14716
rect 8429 14660 8433 14716
rect 8369 14656 8433 14660
rect 8449 14716 8513 14720
rect 8449 14660 8453 14716
rect 8453 14660 8509 14716
rect 8509 14660 8513 14716
rect 8449 14656 8513 14660
rect 8529 14716 8593 14720
rect 8529 14660 8533 14716
rect 8533 14660 8589 14716
rect 8589 14660 8593 14716
rect 8529 14656 8593 14660
rect 8609 14716 8673 14720
rect 8609 14660 8613 14716
rect 8613 14660 8669 14716
rect 8669 14660 8673 14716
rect 8609 14656 8673 14660
rect 13314 14716 13378 14720
rect 13314 14660 13318 14716
rect 13318 14660 13374 14716
rect 13374 14660 13378 14716
rect 13314 14656 13378 14660
rect 13394 14716 13458 14720
rect 13394 14660 13398 14716
rect 13398 14660 13454 14716
rect 13454 14660 13458 14716
rect 13394 14656 13458 14660
rect 13474 14716 13538 14720
rect 13474 14660 13478 14716
rect 13478 14660 13534 14716
rect 13534 14660 13538 14716
rect 13474 14656 13538 14660
rect 13554 14716 13618 14720
rect 13554 14660 13558 14716
rect 13558 14660 13614 14716
rect 13614 14660 13618 14716
rect 13554 14656 13618 14660
rect 18259 14716 18323 14720
rect 18259 14660 18263 14716
rect 18263 14660 18319 14716
rect 18319 14660 18323 14716
rect 18259 14656 18323 14660
rect 18339 14716 18403 14720
rect 18339 14660 18343 14716
rect 18343 14660 18399 14716
rect 18399 14660 18403 14716
rect 18339 14656 18403 14660
rect 18419 14716 18483 14720
rect 18419 14660 18423 14716
rect 18423 14660 18479 14716
rect 18479 14660 18483 14716
rect 18419 14656 18483 14660
rect 18499 14716 18563 14720
rect 18499 14660 18503 14716
rect 18503 14660 18559 14716
rect 18559 14660 18563 14716
rect 18499 14656 18563 14660
rect 5896 14172 5960 14176
rect 5896 14116 5900 14172
rect 5900 14116 5956 14172
rect 5956 14116 5960 14172
rect 5896 14112 5960 14116
rect 5976 14172 6040 14176
rect 5976 14116 5980 14172
rect 5980 14116 6036 14172
rect 6036 14116 6040 14172
rect 5976 14112 6040 14116
rect 6056 14172 6120 14176
rect 6056 14116 6060 14172
rect 6060 14116 6116 14172
rect 6116 14116 6120 14172
rect 6056 14112 6120 14116
rect 6136 14172 6200 14176
rect 6136 14116 6140 14172
rect 6140 14116 6196 14172
rect 6196 14116 6200 14172
rect 6136 14112 6200 14116
rect 10841 14172 10905 14176
rect 10841 14116 10845 14172
rect 10845 14116 10901 14172
rect 10901 14116 10905 14172
rect 10841 14112 10905 14116
rect 10921 14172 10985 14176
rect 10921 14116 10925 14172
rect 10925 14116 10981 14172
rect 10981 14116 10985 14172
rect 10921 14112 10985 14116
rect 11001 14172 11065 14176
rect 11001 14116 11005 14172
rect 11005 14116 11061 14172
rect 11061 14116 11065 14172
rect 11001 14112 11065 14116
rect 11081 14172 11145 14176
rect 11081 14116 11085 14172
rect 11085 14116 11141 14172
rect 11141 14116 11145 14172
rect 11081 14112 11145 14116
rect 15786 14172 15850 14176
rect 15786 14116 15790 14172
rect 15790 14116 15846 14172
rect 15846 14116 15850 14172
rect 15786 14112 15850 14116
rect 15866 14172 15930 14176
rect 15866 14116 15870 14172
rect 15870 14116 15926 14172
rect 15926 14116 15930 14172
rect 15866 14112 15930 14116
rect 15946 14172 16010 14176
rect 15946 14116 15950 14172
rect 15950 14116 16006 14172
rect 16006 14116 16010 14172
rect 15946 14112 16010 14116
rect 16026 14172 16090 14176
rect 16026 14116 16030 14172
rect 16030 14116 16086 14172
rect 16086 14116 16090 14172
rect 16026 14112 16090 14116
rect 20731 14172 20795 14176
rect 20731 14116 20735 14172
rect 20735 14116 20791 14172
rect 20791 14116 20795 14172
rect 20731 14112 20795 14116
rect 20811 14172 20875 14176
rect 20811 14116 20815 14172
rect 20815 14116 20871 14172
rect 20871 14116 20875 14172
rect 20811 14112 20875 14116
rect 20891 14172 20955 14176
rect 20891 14116 20895 14172
rect 20895 14116 20951 14172
rect 20951 14116 20955 14172
rect 20891 14112 20955 14116
rect 20971 14172 21035 14176
rect 20971 14116 20975 14172
rect 20975 14116 21031 14172
rect 21031 14116 21035 14172
rect 20971 14112 21035 14116
rect 3424 13628 3488 13632
rect 3424 13572 3428 13628
rect 3428 13572 3484 13628
rect 3484 13572 3488 13628
rect 3424 13568 3488 13572
rect 3504 13628 3568 13632
rect 3504 13572 3508 13628
rect 3508 13572 3564 13628
rect 3564 13572 3568 13628
rect 3504 13568 3568 13572
rect 3584 13628 3648 13632
rect 3584 13572 3588 13628
rect 3588 13572 3644 13628
rect 3644 13572 3648 13628
rect 3584 13568 3648 13572
rect 3664 13628 3728 13632
rect 3664 13572 3668 13628
rect 3668 13572 3724 13628
rect 3724 13572 3728 13628
rect 3664 13568 3728 13572
rect 8369 13628 8433 13632
rect 8369 13572 8373 13628
rect 8373 13572 8429 13628
rect 8429 13572 8433 13628
rect 8369 13568 8433 13572
rect 8449 13628 8513 13632
rect 8449 13572 8453 13628
rect 8453 13572 8509 13628
rect 8509 13572 8513 13628
rect 8449 13568 8513 13572
rect 8529 13628 8593 13632
rect 8529 13572 8533 13628
rect 8533 13572 8589 13628
rect 8589 13572 8593 13628
rect 8529 13568 8593 13572
rect 8609 13628 8673 13632
rect 8609 13572 8613 13628
rect 8613 13572 8669 13628
rect 8669 13572 8673 13628
rect 8609 13568 8673 13572
rect 13314 13628 13378 13632
rect 13314 13572 13318 13628
rect 13318 13572 13374 13628
rect 13374 13572 13378 13628
rect 13314 13568 13378 13572
rect 13394 13628 13458 13632
rect 13394 13572 13398 13628
rect 13398 13572 13454 13628
rect 13454 13572 13458 13628
rect 13394 13568 13458 13572
rect 13474 13628 13538 13632
rect 13474 13572 13478 13628
rect 13478 13572 13534 13628
rect 13534 13572 13538 13628
rect 13474 13568 13538 13572
rect 13554 13628 13618 13632
rect 13554 13572 13558 13628
rect 13558 13572 13614 13628
rect 13614 13572 13618 13628
rect 13554 13568 13618 13572
rect 18259 13628 18323 13632
rect 18259 13572 18263 13628
rect 18263 13572 18319 13628
rect 18319 13572 18323 13628
rect 18259 13568 18323 13572
rect 18339 13628 18403 13632
rect 18339 13572 18343 13628
rect 18343 13572 18399 13628
rect 18399 13572 18403 13628
rect 18339 13568 18403 13572
rect 18419 13628 18483 13632
rect 18419 13572 18423 13628
rect 18423 13572 18479 13628
rect 18479 13572 18483 13628
rect 18419 13568 18483 13572
rect 18499 13628 18563 13632
rect 18499 13572 18503 13628
rect 18503 13572 18559 13628
rect 18559 13572 18563 13628
rect 18499 13568 18563 13572
rect 5896 13084 5960 13088
rect 5896 13028 5900 13084
rect 5900 13028 5956 13084
rect 5956 13028 5960 13084
rect 5896 13024 5960 13028
rect 5976 13084 6040 13088
rect 5976 13028 5980 13084
rect 5980 13028 6036 13084
rect 6036 13028 6040 13084
rect 5976 13024 6040 13028
rect 6056 13084 6120 13088
rect 6056 13028 6060 13084
rect 6060 13028 6116 13084
rect 6116 13028 6120 13084
rect 6056 13024 6120 13028
rect 6136 13084 6200 13088
rect 6136 13028 6140 13084
rect 6140 13028 6196 13084
rect 6196 13028 6200 13084
rect 6136 13024 6200 13028
rect 10841 13084 10905 13088
rect 10841 13028 10845 13084
rect 10845 13028 10901 13084
rect 10901 13028 10905 13084
rect 10841 13024 10905 13028
rect 10921 13084 10985 13088
rect 10921 13028 10925 13084
rect 10925 13028 10981 13084
rect 10981 13028 10985 13084
rect 10921 13024 10985 13028
rect 11001 13084 11065 13088
rect 11001 13028 11005 13084
rect 11005 13028 11061 13084
rect 11061 13028 11065 13084
rect 11001 13024 11065 13028
rect 11081 13084 11145 13088
rect 11081 13028 11085 13084
rect 11085 13028 11141 13084
rect 11141 13028 11145 13084
rect 11081 13024 11145 13028
rect 15786 13084 15850 13088
rect 15786 13028 15790 13084
rect 15790 13028 15846 13084
rect 15846 13028 15850 13084
rect 15786 13024 15850 13028
rect 15866 13084 15930 13088
rect 15866 13028 15870 13084
rect 15870 13028 15926 13084
rect 15926 13028 15930 13084
rect 15866 13024 15930 13028
rect 15946 13084 16010 13088
rect 15946 13028 15950 13084
rect 15950 13028 16006 13084
rect 16006 13028 16010 13084
rect 15946 13024 16010 13028
rect 16026 13084 16090 13088
rect 16026 13028 16030 13084
rect 16030 13028 16086 13084
rect 16086 13028 16090 13084
rect 16026 13024 16090 13028
rect 20731 13084 20795 13088
rect 20731 13028 20735 13084
rect 20735 13028 20791 13084
rect 20791 13028 20795 13084
rect 20731 13024 20795 13028
rect 20811 13084 20875 13088
rect 20811 13028 20815 13084
rect 20815 13028 20871 13084
rect 20871 13028 20875 13084
rect 20811 13024 20875 13028
rect 20891 13084 20955 13088
rect 20891 13028 20895 13084
rect 20895 13028 20951 13084
rect 20951 13028 20955 13084
rect 20891 13024 20955 13028
rect 20971 13084 21035 13088
rect 20971 13028 20975 13084
rect 20975 13028 21031 13084
rect 21031 13028 21035 13084
rect 20971 13024 21035 13028
rect 3424 12540 3488 12544
rect 3424 12484 3428 12540
rect 3428 12484 3484 12540
rect 3484 12484 3488 12540
rect 3424 12480 3488 12484
rect 3504 12540 3568 12544
rect 3504 12484 3508 12540
rect 3508 12484 3564 12540
rect 3564 12484 3568 12540
rect 3504 12480 3568 12484
rect 3584 12540 3648 12544
rect 3584 12484 3588 12540
rect 3588 12484 3644 12540
rect 3644 12484 3648 12540
rect 3584 12480 3648 12484
rect 3664 12540 3728 12544
rect 3664 12484 3668 12540
rect 3668 12484 3724 12540
rect 3724 12484 3728 12540
rect 3664 12480 3728 12484
rect 8369 12540 8433 12544
rect 8369 12484 8373 12540
rect 8373 12484 8429 12540
rect 8429 12484 8433 12540
rect 8369 12480 8433 12484
rect 8449 12540 8513 12544
rect 8449 12484 8453 12540
rect 8453 12484 8509 12540
rect 8509 12484 8513 12540
rect 8449 12480 8513 12484
rect 8529 12540 8593 12544
rect 8529 12484 8533 12540
rect 8533 12484 8589 12540
rect 8589 12484 8593 12540
rect 8529 12480 8593 12484
rect 8609 12540 8673 12544
rect 8609 12484 8613 12540
rect 8613 12484 8669 12540
rect 8669 12484 8673 12540
rect 8609 12480 8673 12484
rect 13314 12540 13378 12544
rect 13314 12484 13318 12540
rect 13318 12484 13374 12540
rect 13374 12484 13378 12540
rect 13314 12480 13378 12484
rect 13394 12540 13458 12544
rect 13394 12484 13398 12540
rect 13398 12484 13454 12540
rect 13454 12484 13458 12540
rect 13394 12480 13458 12484
rect 13474 12540 13538 12544
rect 13474 12484 13478 12540
rect 13478 12484 13534 12540
rect 13534 12484 13538 12540
rect 13474 12480 13538 12484
rect 13554 12540 13618 12544
rect 13554 12484 13558 12540
rect 13558 12484 13614 12540
rect 13614 12484 13618 12540
rect 13554 12480 13618 12484
rect 18259 12540 18323 12544
rect 18259 12484 18263 12540
rect 18263 12484 18319 12540
rect 18319 12484 18323 12540
rect 18259 12480 18323 12484
rect 18339 12540 18403 12544
rect 18339 12484 18343 12540
rect 18343 12484 18399 12540
rect 18399 12484 18403 12540
rect 18339 12480 18403 12484
rect 18419 12540 18483 12544
rect 18419 12484 18423 12540
rect 18423 12484 18479 12540
rect 18479 12484 18483 12540
rect 18419 12480 18483 12484
rect 18499 12540 18563 12544
rect 18499 12484 18503 12540
rect 18503 12484 18559 12540
rect 18559 12484 18563 12540
rect 18499 12480 18563 12484
rect 5896 11996 5960 12000
rect 5896 11940 5900 11996
rect 5900 11940 5956 11996
rect 5956 11940 5960 11996
rect 5896 11936 5960 11940
rect 5976 11996 6040 12000
rect 5976 11940 5980 11996
rect 5980 11940 6036 11996
rect 6036 11940 6040 11996
rect 5976 11936 6040 11940
rect 6056 11996 6120 12000
rect 6056 11940 6060 11996
rect 6060 11940 6116 11996
rect 6116 11940 6120 11996
rect 6056 11936 6120 11940
rect 6136 11996 6200 12000
rect 6136 11940 6140 11996
rect 6140 11940 6196 11996
rect 6196 11940 6200 11996
rect 6136 11936 6200 11940
rect 10841 11996 10905 12000
rect 10841 11940 10845 11996
rect 10845 11940 10901 11996
rect 10901 11940 10905 11996
rect 10841 11936 10905 11940
rect 10921 11996 10985 12000
rect 10921 11940 10925 11996
rect 10925 11940 10981 11996
rect 10981 11940 10985 11996
rect 10921 11936 10985 11940
rect 11001 11996 11065 12000
rect 11001 11940 11005 11996
rect 11005 11940 11061 11996
rect 11061 11940 11065 11996
rect 11001 11936 11065 11940
rect 11081 11996 11145 12000
rect 11081 11940 11085 11996
rect 11085 11940 11141 11996
rect 11141 11940 11145 11996
rect 11081 11936 11145 11940
rect 15786 11996 15850 12000
rect 15786 11940 15790 11996
rect 15790 11940 15846 11996
rect 15846 11940 15850 11996
rect 15786 11936 15850 11940
rect 15866 11996 15930 12000
rect 15866 11940 15870 11996
rect 15870 11940 15926 11996
rect 15926 11940 15930 11996
rect 15866 11936 15930 11940
rect 15946 11996 16010 12000
rect 15946 11940 15950 11996
rect 15950 11940 16006 11996
rect 16006 11940 16010 11996
rect 15946 11936 16010 11940
rect 16026 11996 16090 12000
rect 16026 11940 16030 11996
rect 16030 11940 16086 11996
rect 16086 11940 16090 11996
rect 16026 11936 16090 11940
rect 20731 11996 20795 12000
rect 20731 11940 20735 11996
rect 20735 11940 20791 11996
rect 20791 11940 20795 11996
rect 20731 11936 20795 11940
rect 20811 11996 20875 12000
rect 20811 11940 20815 11996
rect 20815 11940 20871 11996
rect 20871 11940 20875 11996
rect 20811 11936 20875 11940
rect 20891 11996 20955 12000
rect 20891 11940 20895 11996
rect 20895 11940 20951 11996
rect 20951 11940 20955 11996
rect 20891 11936 20955 11940
rect 20971 11996 21035 12000
rect 20971 11940 20975 11996
rect 20975 11940 21031 11996
rect 21031 11940 21035 11996
rect 20971 11936 21035 11940
rect 3424 11452 3488 11456
rect 3424 11396 3428 11452
rect 3428 11396 3484 11452
rect 3484 11396 3488 11452
rect 3424 11392 3488 11396
rect 3504 11452 3568 11456
rect 3504 11396 3508 11452
rect 3508 11396 3564 11452
rect 3564 11396 3568 11452
rect 3504 11392 3568 11396
rect 3584 11452 3648 11456
rect 3584 11396 3588 11452
rect 3588 11396 3644 11452
rect 3644 11396 3648 11452
rect 3584 11392 3648 11396
rect 3664 11452 3728 11456
rect 3664 11396 3668 11452
rect 3668 11396 3724 11452
rect 3724 11396 3728 11452
rect 3664 11392 3728 11396
rect 8369 11452 8433 11456
rect 8369 11396 8373 11452
rect 8373 11396 8429 11452
rect 8429 11396 8433 11452
rect 8369 11392 8433 11396
rect 8449 11452 8513 11456
rect 8449 11396 8453 11452
rect 8453 11396 8509 11452
rect 8509 11396 8513 11452
rect 8449 11392 8513 11396
rect 8529 11452 8593 11456
rect 8529 11396 8533 11452
rect 8533 11396 8589 11452
rect 8589 11396 8593 11452
rect 8529 11392 8593 11396
rect 8609 11452 8673 11456
rect 8609 11396 8613 11452
rect 8613 11396 8669 11452
rect 8669 11396 8673 11452
rect 8609 11392 8673 11396
rect 13314 11452 13378 11456
rect 13314 11396 13318 11452
rect 13318 11396 13374 11452
rect 13374 11396 13378 11452
rect 13314 11392 13378 11396
rect 13394 11452 13458 11456
rect 13394 11396 13398 11452
rect 13398 11396 13454 11452
rect 13454 11396 13458 11452
rect 13394 11392 13458 11396
rect 13474 11452 13538 11456
rect 13474 11396 13478 11452
rect 13478 11396 13534 11452
rect 13534 11396 13538 11452
rect 13474 11392 13538 11396
rect 13554 11452 13618 11456
rect 13554 11396 13558 11452
rect 13558 11396 13614 11452
rect 13614 11396 13618 11452
rect 13554 11392 13618 11396
rect 18259 11452 18323 11456
rect 18259 11396 18263 11452
rect 18263 11396 18319 11452
rect 18319 11396 18323 11452
rect 18259 11392 18323 11396
rect 18339 11452 18403 11456
rect 18339 11396 18343 11452
rect 18343 11396 18399 11452
rect 18399 11396 18403 11452
rect 18339 11392 18403 11396
rect 18419 11452 18483 11456
rect 18419 11396 18423 11452
rect 18423 11396 18479 11452
rect 18479 11396 18483 11452
rect 18419 11392 18483 11396
rect 18499 11452 18563 11456
rect 18499 11396 18503 11452
rect 18503 11396 18559 11452
rect 18559 11396 18563 11452
rect 18499 11392 18563 11396
rect 5896 10908 5960 10912
rect 5896 10852 5900 10908
rect 5900 10852 5956 10908
rect 5956 10852 5960 10908
rect 5896 10848 5960 10852
rect 5976 10908 6040 10912
rect 5976 10852 5980 10908
rect 5980 10852 6036 10908
rect 6036 10852 6040 10908
rect 5976 10848 6040 10852
rect 6056 10908 6120 10912
rect 6056 10852 6060 10908
rect 6060 10852 6116 10908
rect 6116 10852 6120 10908
rect 6056 10848 6120 10852
rect 6136 10908 6200 10912
rect 6136 10852 6140 10908
rect 6140 10852 6196 10908
rect 6196 10852 6200 10908
rect 6136 10848 6200 10852
rect 10841 10908 10905 10912
rect 10841 10852 10845 10908
rect 10845 10852 10901 10908
rect 10901 10852 10905 10908
rect 10841 10848 10905 10852
rect 10921 10908 10985 10912
rect 10921 10852 10925 10908
rect 10925 10852 10981 10908
rect 10981 10852 10985 10908
rect 10921 10848 10985 10852
rect 11001 10908 11065 10912
rect 11001 10852 11005 10908
rect 11005 10852 11061 10908
rect 11061 10852 11065 10908
rect 11001 10848 11065 10852
rect 11081 10908 11145 10912
rect 11081 10852 11085 10908
rect 11085 10852 11141 10908
rect 11141 10852 11145 10908
rect 11081 10848 11145 10852
rect 15786 10908 15850 10912
rect 15786 10852 15790 10908
rect 15790 10852 15846 10908
rect 15846 10852 15850 10908
rect 15786 10848 15850 10852
rect 15866 10908 15930 10912
rect 15866 10852 15870 10908
rect 15870 10852 15926 10908
rect 15926 10852 15930 10908
rect 15866 10848 15930 10852
rect 15946 10908 16010 10912
rect 15946 10852 15950 10908
rect 15950 10852 16006 10908
rect 16006 10852 16010 10908
rect 15946 10848 16010 10852
rect 16026 10908 16090 10912
rect 16026 10852 16030 10908
rect 16030 10852 16086 10908
rect 16086 10852 16090 10908
rect 16026 10848 16090 10852
rect 20731 10908 20795 10912
rect 20731 10852 20735 10908
rect 20735 10852 20791 10908
rect 20791 10852 20795 10908
rect 20731 10848 20795 10852
rect 20811 10908 20875 10912
rect 20811 10852 20815 10908
rect 20815 10852 20871 10908
rect 20871 10852 20875 10908
rect 20811 10848 20875 10852
rect 20891 10908 20955 10912
rect 20891 10852 20895 10908
rect 20895 10852 20951 10908
rect 20951 10852 20955 10908
rect 20891 10848 20955 10852
rect 20971 10908 21035 10912
rect 20971 10852 20975 10908
rect 20975 10852 21031 10908
rect 21031 10852 21035 10908
rect 20971 10848 21035 10852
rect 3424 10364 3488 10368
rect 3424 10308 3428 10364
rect 3428 10308 3484 10364
rect 3484 10308 3488 10364
rect 3424 10304 3488 10308
rect 3504 10364 3568 10368
rect 3504 10308 3508 10364
rect 3508 10308 3564 10364
rect 3564 10308 3568 10364
rect 3504 10304 3568 10308
rect 3584 10364 3648 10368
rect 3584 10308 3588 10364
rect 3588 10308 3644 10364
rect 3644 10308 3648 10364
rect 3584 10304 3648 10308
rect 3664 10364 3728 10368
rect 3664 10308 3668 10364
rect 3668 10308 3724 10364
rect 3724 10308 3728 10364
rect 3664 10304 3728 10308
rect 8369 10364 8433 10368
rect 8369 10308 8373 10364
rect 8373 10308 8429 10364
rect 8429 10308 8433 10364
rect 8369 10304 8433 10308
rect 8449 10364 8513 10368
rect 8449 10308 8453 10364
rect 8453 10308 8509 10364
rect 8509 10308 8513 10364
rect 8449 10304 8513 10308
rect 8529 10364 8593 10368
rect 8529 10308 8533 10364
rect 8533 10308 8589 10364
rect 8589 10308 8593 10364
rect 8529 10304 8593 10308
rect 8609 10364 8673 10368
rect 8609 10308 8613 10364
rect 8613 10308 8669 10364
rect 8669 10308 8673 10364
rect 8609 10304 8673 10308
rect 13314 10364 13378 10368
rect 13314 10308 13318 10364
rect 13318 10308 13374 10364
rect 13374 10308 13378 10364
rect 13314 10304 13378 10308
rect 13394 10364 13458 10368
rect 13394 10308 13398 10364
rect 13398 10308 13454 10364
rect 13454 10308 13458 10364
rect 13394 10304 13458 10308
rect 13474 10364 13538 10368
rect 13474 10308 13478 10364
rect 13478 10308 13534 10364
rect 13534 10308 13538 10364
rect 13474 10304 13538 10308
rect 13554 10364 13618 10368
rect 13554 10308 13558 10364
rect 13558 10308 13614 10364
rect 13614 10308 13618 10364
rect 13554 10304 13618 10308
rect 18259 10364 18323 10368
rect 18259 10308 18263 10364
rect 18263 10308 18319 10364
rect 18319 10308 18323 10364
rect 18259 10304 18323 10308
rect 18339 10364 18403 10368
rect 18339 10308 18343 10364
rect 18343 10308 18399 10364
rect 18399 10308 18403 10364
rect 18339 10304 18403 10308
rect 18419 10364 18483 10368
rect 18419 10308 18423 10364
rect 18423 10308 18479 10364
rect 18479 10308 18483 10364
rect 18419 10304 18483 10308
rect 18499 10364 18563 10368
rect 18499 10308 18503 10364
rect 18503 10308 18559 10364
rect 18559 10308 18563 10364
rect 18499 10304 18563 10308
rect 5896 9820 5960 9824
rect 5896 9764 5900 9820
rect 5900 9764 5956 9820
rect 5956 9764 5960 9820
rect 5896 9760 5960 9764
rect 5976 9820 6040 9824
rect 5976 9764 5980 9820
rect 5980 9764 6036 9820
rect 6036 9764 6040 9820
rect 5976 9760 6040 9764
rect 6056 9820 6120 9824
rect 6056 9764 6060 9820
rect 6060 9764 6116 9820
rect 6116 9764 6120 9820
rect 6056 9760 6120 9764
rect 6136 9820 6200 9824
rect 6136 9764 6140 9820
rect 6140 9764 6196 9820
rect 6196 9764 6200 9820
rect 6136 9760 6200 9764
rect 10841 9820 10905 9824
rect 10841 9764 10845 9820
rect 10845 9764 10901 9820
rect 10901 9764 10905 9820
rect 10841 9760 10905 9764
rect 10921 9820 10985 9824
rect 10921 9764 10925 9820
rect 10925 9764 10981 9820
rect 10981 9764 10985 9820
rect 10921 9760 10985 9764
rect 11001 9820 11065 9824
rect 11001 9764 11005 9820
rect 11005 9764 11061 9820
rect 11061 9764 11065 9820
rect 11001 9760 11065 9764
rect 11081 9820 11145 9824
rect 11081 9764 11085 9820
rect 11085 9764 11141 9820
rect 11141 9764 11145 9820
rect 11081 9760 11145 9764
rect 15786 9820 15850 9824
rect 15786 9764 15790 9820
rect 15790 9764 15846 9820
rect 15846 9764 15850 9820
rect 15786 9760 15850 9764
rect 15866 9820 15930 9824
rect 15866 9764 15870 9820
rect 15870 9764 15926 9820
rect 15926 9764 15930 9820
rect 15866 9760 15930 9764
rect 15946 9820 16010 9824
rect 15946 9764 15950 9820
rect 15950 9764 16006 9820
rect 16006 9764 16010 9820
rect 15946 9760 16010 9764
rect 16026 9820 16090 9824
rect 16026 9764 16030 9820
rect 16030 9764 16086 9820
rect 16086 9764 16090 9820
rect 16026 9760 16090 9764
rect 20731 9820 20795 9824
rect 20731 9764 20735 9820
rect 20735 9764 20791 9820
rect 20791 9764 20795 9820
rect 20731 9760 20795 9764
rect 20811 9820 20875 9824
rect 20811 9764 20815 9820
rect 20815 9764 20871 9820
rect 20871 9764 20875 9820
rect 20811 9760 20875 9764
rect 20891 9820 20955 9824
rect 20891 9764 20895 9820
rect 20895 9764 20951 9820
rect 20951 9764 20955 9820
rect 20891 9760 20955 9764
rect 20971 9820 21035 9824
rect 20971 9764 20975 9820
rect 20975 9764 21031 9820
rect 21031 9764 21035 9820
rect 20971 9760 21035 9764
rect 3424 9276 3488 9280
rect 3424 9220 3428 9276
rect 3428 9220 3484 9276
rect 3484 9220 3488 9276
rect 3424 9216 3488 9220
rect 3504 9276 3568 9280
rect 3504 9220 3508 9276
rect 3508 9220 3564 9276
rect 3564 9220 3568 9276
rect 3504 9216 3568 9220
rect 3584 9276 3648 9280
rect 3584 9220 3588 9276
rect 3588 9220 3644 9276
rect 3644 9220 3648 9276
rect 3584 9216 3648 9220
rect 3664 9276 3728 9280
rect 3664 9220 3668 9276
rect 3668 9220 3724 9276
rect 3724 9220 3728 9276
rect 3664 9216 3728 9220
rect 8369 9276 8433 9280
rect 8369 9220 8373 9276
rect 8373 9220 8429 9276
rect 8429 9220 8433 9276
rect 8369 9216 8433 9220
rect 8449 9276 8513 9280
rect 8449 9220 8453 9276
rect 8453 9220 8509 9276
rect 8509 9220 8513 9276
rect 8449 9216 8513 9220
rect 8529 9276 8593 9280
rect 8529 9220 8533 9276
rect 8533 9220 8589 9276
rect 8589 9220 8593 9276
rect 8529 9216 8593 9220
rect 8609 9276 8673 9280
rect 8609 9220 8613 9276
rect 8613 9220 8669 9276
rect 8669 9220 8673 9276
rect 8609 9216 8673 9220
rect 13314 9276 13378 9280
rect 13314 9220 13318 9276
rect 13318 9220 13374 9276
rect 13374 9220 13378 9276
rect 13314 9216 13378 9220
rect 13394 9276 13458 9280
rect 13394 9220 13398 9276
rect 13398 9220 13454 9276
rect 13454 9220 13458 9276
rect 13394 9216 13458 9220
rect 13474 9276 13538 9280
rect 13474 9220 13478 9276
rect 13478 9220 13534 9276
rect 13534 9220 13538 9276
rect 13474 9216 13538 9220
rect 13554 9276 13618 9280
rect 13554 9220 13558 9276
rect 13558 9220 13614 9276
rect 13614 9220 13618 9276
rect 13554 9216 13618 9220
rect 18259 9276 18323 9280
rect 18259 9220 18263 9276
rect 18263 9220 18319 9276
rect 18319 9220 18323 9276
rect 18259 9216 18323 9220
rect 18339 9276 18403 9280
rect 18339 9220 18343 9276
rect 18343 9220 18399 9276
rect 18399 9220 18403 9276
rect 18339 9216 18403 9220
rect 18419 9276 18483 9280
rect 18419 9220 18423 9276
rect 18423 9220 18479 9276
rect 18479 9220 18483 9276
rect 18419 9216 18483 9220
rect 18499 9276 18563 9280
rect 18499 9220 18503 9276
rect 18503 9220 18559 9276
rect 18559 9220 18563 9276
rect 18499 9216 18563 9220
rect 5896 8732 5960 8736
rect 5896 8676 5900 8732
rect 5900 8676 5956 8732
rect 5956 8676 5960 8732
rect 5896 8672 5960 8676
rect 5976 8732 6040 8736
rect 5976 8676 5980 8732
rect 5980 8676 6036 8732
rect 6036 8676 6040 8732
rect 5976 8672 6040 8676
rect 6056 8732 6120 8736
rect 6056 8676 6060 8732
rect 6060 8676 6116 8732
rect 6116 8676 6120 8732
rect 6056 8672 6120 8676
rect 6136 8732 6200 8736
rect 6136 8676 6140 8732
rect 6140 8676 6196 8732
rect 6196 8676 6200 8732
rect 6136 8672 6200 8676
rect 10841 8732 10905 8736
rect 10841 8676 10845 8732
rect 10845 8676 10901 8732
rect 10901 8676 10905 8732
rect 10841 8672 10905 8676
rect 10921 8732 10985 8736
rect 10921 8676 10925 8732
rect 10925 8676 10981 8732
rect 10981 8676 10985 8732
rect 10921 8672 10985 8676
rect 11001 8732 11065 8736
rect 11001 8676 11005 8732
rect 11005 8676 11061 8732
rect 11061 8676 11065 8732
rect 11001 8672 11065 8676
rect 11081 8732 11145 8736
rect 11081 8676 11085 8732
rect 11085 8676 11141 8732
rect 11141 8676 11145 8732
rect 11081 8672 11145 8676
rect 15786 8732 15850 8736
rect 15786 8676 15790 8732
rect 15790 8676 15846 8732
rect 15846 8676 15850 8732
rect 15786 8672 15850 8676
rect 15866 8732 15930 8736
rect 15866 8676 15870 8732
rect 15870 8676 15926 8732
rect 15926 8676 15930 8732
rect 15866 8672 15930 8676
rect 15946 8732 16010 8736
rect 15946 8676 15950 8732
rect 15950 8676 16006 8732
rect 16006 8676 16010 8732
rect 15946 8672 16010 8676
rect 16026 8732 16090 8736
rect 16026 8676 16030 8732
rect 16030 8676 16086 8732
rect 16086 8676 16090 8732
rect 16026 8672 16090 8676
rect 20731 8732 20795 8736
rect 20731 8676 20735 8732
rect 20735 8676 20791 8732
rect 20791 8676 20795 8732
rect 20731 8672 20795 8676
rect 20811 8732 20875 8736
rect 20811 8676 20815 8732
rect 20815 8676 20871 8732
rect 20871 8676 20875 8732
rect 20811 8672 20875 8676
rect 20891 8732 20955 8736
rect 20891 8676 20895 8732
rect 20895 8676 20951 8732
rect 20951 8676 20955 8732
rect 20891 8672 20955 8676
rect 20971 8732 21035 8736
rect 20971 8676 20975 8732
rect 20975 8676 21031 8732
rect 21031 8676 21035 8732
rect 20971 8672 21035 8676
rect 3424 8188 3488 8192
rect 3424 8132 3428 8188
rect 3428 8132 3484 8188
rect 3484 8132 3488 8188
rect 3424 8128 3488 8132
rect 3504 8188 3568 8192
rect 3504 8132 3508 8188
rect 3508 8132 3564 8188
rect 3564 8132 3568 8188
rect 3504 8128 3568 8132
rect 3584 8188 3648 8192
rect 3584 8132 3588 8188
rect 3588 8132 3644 8188
rect 3644 8132 3648 8188
rect 3584 8128 3648 8132
rect 3664 8188 3728 8192
rect 3664 8132 3668 8188
rect 3668 8132 3724 8188
rect 3724 8132 3728 8188
rect 3664 8128 3728 8132
rect 8369 8188 8433 8192
rect 8369 8132 8373 8188
rect 8373 8132 8429 8188
rect 8429 8132 8433 8188
rect 8369 8128 8433 8132
rect 8449 8188 8513 8192
rect 8449 8132 8453 8188
rect 8453 8132 8509 8188
rect 8509 8132 8513 8188
rect 8449 8128 8513 8132
rect 8529 8188 8593 8192
rect 8529 8132 8533 8188
rect 8533 8132 8589 8188
rect 8589 8132 8593 8188
rect 8529 8128 8593 8132
rect 8609 8188 8673 8192
rect 8609 8132 8613 8188
rect 8613 8132 8669 8188
rect 8669 8132 8673 8188
rect 8609 8128 8673 8132
rect 13314 8188 13378 8192
rect 13314 8132 13318 8188
rect 13318 8132 13374 8188
rect 13374 8132 13378 8188
rect 13314 8128 13378 8132
rect 13394 8188 13458 8192
rect 13394 8132 13398 8188
rect 13398 8132 13454 8188
rect 13454 8132 13458 8188
rect 13394 8128 13458 8132
rect 13474 8188 13538 8192
rect 13474 8132 13478 8188
rect 13478 8132 13534 8188
rect 13534 8132 13538 8188
rect 13474 8128 13538 8132
rect 13554 8188 13618 8192
rect 13554 8132 13558 8188
rect 13558 8132 13614 8188
rect 13614 8132 13618 8188
rect 13554 8128 13618 8132
rect 18259 8188 18323 8192
rect 18259 8132 18263 8188
rect 18263 8132 18319 8188
rect 18319 8132 18323 8188
rect 18259 8128 18323 8132
rect 18339 8188 18403 8192
rect 18339 8132 18343 8188
rect 18343 8132 18399 8188
rect 18399 8132 18403 8188
rect 18339 8128 18403 8132
rect 18419 8188 18483 8192
rect 18419 8132 18423 8188
rect 18423 8132 18479 8188
rect 18479 8132 18483 8188
rect 18419 8128 18483 8132
rect 18499 8188 18563 8192
rect 18499 8132 18503 8188
rect 18503 8132 18559 8188
rect 18559 8132 18563 8188
rect 18499 8128 18563 8132
rect 5896 7644 5960 7648
rect 5896 7588 5900 7644
rect 5900 7588 5956 7644
rect 5956 7588 5960 7644
rect 5896 7584 5960 7588
rect 5976 7644 6040 7648
rect 5976 7588 5980 7644
rect 5980 7588 6036 7644
rect 6036 7588 6040 7644
rect 5976 7584 6040 7588
rect 6056 7644 6120 7648
rect 6056 7588 6060 7644
rect 6060 7588 6116 7644
rect 6116 7588 6120 7644
rect 6056 7584 6120 7588
rect 6136 7644 6200 7648
rect 6136 7588 6140 7644
rect 6140 7588 6196 7644
rect 6196 7588 6200 7644
rect 6136 7584 6200 7588
rect 10841 7644 10905 7648
rect 10841 7588 10845 7644
rect 10845 7588 10901 7644
rect 10901 7588 10905 7644
rect 10841 7584 10905 7588
rect 10921 7644 10985 7648
rect 10921 7588 10925 7644
rect 10925 7588 10981 7644
rect 10981 7588 10985 7644
rect 10921 7584 10985 7588
rect 11001 7644 11065 7648
rect 11001 7588 11005 7644
rect 11005 7588 11061 7644
rect 11061 7588 11065 7644
rect 11001 7584 11065 7588
rect 11081 7644 11145 7648
rect 11081 7588 11085 7644
rect 11085 7588 11141 7644
rect 11141 7588 11145 7644
rect 11081 7584 11145 7588
rect 15786 7644 15850 7648
rect 15786 7588 15790 7644
rect 15790 7588 15846 7644
rect 15846 7588 15850 7644
rect 15786 7584 15850 7588
rect 15866 7644 15930 7648
rect 15866 7588 15870 7644
rect 15870 7588 15926 7644
rect 15926 7588 15930 7644
rect 15866 7584 15930 7588
rect 15946 7644 16010 7648
rect 15946 7588 15950 7644
rect 15950 7588 16006 7644
rect 16006 7588 16010 7644
rect 15946 7584 16010 7588
rect 16026 7644 16090 7648
rect 16026 7588 16030 7644
rect 16030 7588 16086 7644
rect 16086 7588 16090 7644
rect 16026 7584 16090 7588
rect 20731 7644 20795 7648
rect 20731 7588 20735 7644
rect 20735 7588 20791 7644
rect 20791 7588 20795 7644
rect 20731 7584 20795 7588
rect 20811 7644 20875 7648
rect 20811 7588 20815 7644
rect 20815 7588 20871 7644
rect 20871 7588 20875 7644
rect 20811 7584 20875 7588
rect 20891 7644 20955 7648
rect 20891 7588 20895 7644
rect 20895 7588 20951 7644
rect 20951 7588 20955 7644
rect 20891 7584 20955 7588
rect 20971 7644 21035 7648
rect 20971 7588 20975 7644
rect 20975 7588 21031 7644
rect 21031 7588 21035 7644
rect 20971 7584 21035 7588
rect 3424 7100 3488 7104
rect 3424 7044 3428 7100
rect 3428 7044 3484 7100
rect 3484 7044 3488 7100
rect 3424 7040 3488 7044
rect 3504 7100 3568 7104
rect 3504 7044 3508 7100
rect 3508 7044 3564 7100
rect 3564 7044 3568 7100
rect 3504 7040 3568 7044
rect 3584 7100 3648 7104
rect 3584 7044 3588 7100
rect 3588 7044 3644 7100
rect 3644 7044 3648 7100
rect 3584 7040 3648 7044
rect 3664 7100 3728 7104
rect 3664 7044 3668 7100
rect 3668 7044 3724 7100
rect 3724 7044 3728 7100
rect 3664 7040 3728 7044
rect 8369 7100 8433 7104
rect 8369 7044 8373 7100
rect 8373 7044 8429 7100
rect 8429 7044 8433 7100
rect 8369 7040 8433 7044
rect 8449 7100 8513 7104
rect 8449 7044 8453 7100
rect 8453 7044 8509 7100
rect 8509 7044 8513 7100
rect 8449 7040 8513 7044
rect 8529 7100 8593 7104
rect 8529 7044 8533 7100
rect 8533 7044 8589 7100
rect 8589 7044 8593 7100
rect 8529 7040 8593 7044
rect 8609 7100 8673 7104
rect 8609 7044 8613 7100
rect 8613 7044 8669 7100
rect 8669 7044 8673 7100
rect 8609 7040 8673 7044
rect 13314 7100 13378 7104
rect 13314 7044 13318 7100
rect 13318 7044 13374 7100
rect 13374 7044 13378 7100
rect 13314 7040 13378 7044
rect 13394 7100 13458 7104
rect 13394 7044 13398 7100
rect 13398 7044 13454 7100
rect 13454 7044 13458 7100
rect 13394 7040 13458 7044
rect 13474 7100 13538 7104
rect 13474 7044 13478 7100
rect 13478 7044 13534 7100
rect 13534 7044 13538 7100
rect 13474 7040 13538 7044
rect 13554 7100 13618 7104
rect 13554 7044 13558 7100
rect 13558 7044 13614 7100
rect 13614 7044 13618 7100
rect 13554 7040 13618 7044
rect 18259 7100 18323 7104
rect 18259 7044 18263 7100
rect 18263 7044 18319 7100
rect 18319 7044 18323 7100
rect 18259 7040 18323 7044
rect 18339 7100 18403 7104
rect 18339 7044 18343 7100
rect 18343 7044 18399 7100
rect 18399 7044 18403 7100
rect 18339 7040 18403 7044
rect 18419 7100 18483 7104
rect 18419 7044 18423 7100
rect 18423 7044 18479 7100
rect 18479 7044 18483 7100
rect 18419 7040 18483 7044
rect 18499 7100 18563 7104
rect 18499 7044 18503 7100
rect 18503 7044 18559 7100
rect 18559 7044 18563 7100
rect 18499 7040 18563 7044
rect 5896 6556 5960 6560
rect 5896 6500 5900 6556
rect 5900 6500 5956 6556
rect 5956 6500 5960 6556
rect 5896 6496 5960 6500
rect 5976 6556 6040 6560
rect 5976 6500 5980 6556
rect 5980 6500 6036 6556
rect 6036 6500 6040 6556
rect 5976 6496 6040 6500
rect 6056 6556 6120 6560
rect 6056 6500 6060 6556
rect 6060 6500 6116 6556
rect 6116 6500 6120 6556
rect 6056 6496 6120 6500
rect 6136 6556 6200 6560
rect 6136 6500 6140 6556
rect 6140 6500 6196 6556
rect 6196 6500 6200 6556
rect 6136 6496 6200 6500
rect 10841 6556 10905 6560
rect 10841 6500 10845 6556
rect 10845 6500 10901 6556
rect 10901 6500 10905 6556
rect 10841 6496 10905 6500
rect 10921 6556 10985 6560
rect 10921 6500 10925 6556
rect 10925 6500 10981 6556
rect 10981 6500 10985 6556
rect 10921 6496 10985 6500
rect 11001 6556 11065 6560
rect 11001 6500 11005 6556
rect 11005 6500 11061 6556
rect 11061 6500 11065 6556
rect 11001 6496 11065 6500
rect 11081 6556 11145 6560
rect 11081 6500 11085 6556
rect 11085 6500 11141 6556
rect 11141 6500 11145 6556
rect 11081 6496 11145 6500
rect 15786 6556 15850 6560
rect 15786 6500 15790 6556
rect 15790 6500 15846 6556
rect 15846 6500 15850 6556
rect 15786 6496 15850 6500
rect 15866 6556 15930 6560
rect 15866 6500 15870 6556
rect 15870 6500 15926 6556
rect 15926 6500 15930 6556
rect 15866 6496 15930 6500
rect 15946 6556 16010 6560
rect 15946 6500 15950 6556
rect 15950 6500 16006 6556
rect 16006 6500 16010 6556
rect 15946 6496 16010 6500
rect 16026 6556 16090 6560
rect 16026 6500 16030 6556
rect 16030 6500 16086 6556
rect 16086 6500 16090 6556
rect 16026 6496 16090 6500
rect 20731 6556 20795 6560
rect 20731 6500 20735 6556
rect 20735 6500 20791 6556
rect 20791 6500 20795 6556
rect 20731 6496 20795 6500
rect 20811 6556 20875 6560
rect 20811 6500 20815 6556
rect 20815 6500 20871 6556
rect 20871 6500 20875 6556
rect 20811 6496 20875 6500
rect 20891 6556 20955 6560
rect 20891 6500 20895 6556
rect 20895 6500 20951 6556
rect 20951 6500 20955 6556
rect 20891 6496 20955 6500
rect 20971 6556 21035 6560
rect 20971 6500 20975 6556
rect 20975 6500 21031 6556
rect 21031 6500 21035 6556
rect 20971 6496 21035 6500
rect 3424 6012 3488 6016
rect 3424 5956 3428 6012
rect 3428 5956 3484 6012
rect 3484 5956 3488 6012
rect 3424 5952 3488 5956
rect 3504 6012 3568 6016
rect 3504 5956 3508 6012
rect 3508 5956 3564 6012
rect 3564 5956 3568 6012
rect 3504 5952 3568 5956
rect 3584 6012 3648 6016
rect 3584 5956 3588 6012
rect 3588 5956 3644 6012
rect 3644 5956 3648 6012
rect 3584 5952 3648 5956
rect 3664 6012 3728 6016
rect 3664 5956 3668 6012
rect 3668 5956 3724 6012
rect 3724 5956 3728 6012
rect 3664 5952 3728 5956
rect 8369 6012 8433 6016
rect 8369 5956 8373 6012
rect 8373 5956 8429 6012
rect 8429 5956 8433 6012
rect 8369 5952 8433 5956
rect 8449 6012 8513 6016
rect 8449 5956 8453 6012
rect 8453 5956 8509 6012
rect 8509 5956 8513 6012
rect 8449 5952 8513 5956
rect 8529 6012 8593 6016
rect 8529 5956 8533 6012
rect 8533 5956 8589 6012
rect 8589 5956 8593 6012
rect 8529 5952 8593 5956
rect 8609 6012 8673 6016
rect 8609 5956 8613 6012
rect 8613 5956 8669 6012
rect 8669 5956 8673 6012
rect 8609 5952 8673 5956
rect 13314 6012 13378 6016
rect 13314 5956 13318 6012
rect 13318 5956 13374 6012
rect 13374 5956 13378 6012
rect 13314 5952 13378 5956
rect 13394 6012 13458 6016
rect 13394 5956 13398 6012
rect 13398 5956 13454 6012
rect 13454 5956 13458 6012
rect 13394 5952 13458 5956
rect 13474 6012 13538 6016
rect 13474 5956 13478 6012
rect 13478 5956 13534 6012
rect 13534 5956 13538 6012
rect 13474 5952 13538 5956
rect 13554 6012 13618 6016
rect 13554 5956 13558 6012
rect 13558 5956 13614 6012
rect 13614 5956 13618 6012
rect 13554 5952 13618 5956
rect 18259 6012 18323 6016
rect 18259 5956 18263 6012
rect 18263 5956 18319 6012
rect 18319 5956 18323 6012
rect 18259 5952 18323 5956
rect 18339 6012 18403 6016
rect 18339 5956 18343 6012
rect 18343 5956 18399 6012
rect 18399 5956 18403 6012
rect 18339 5952 18403 5956
rect 18419 6012 18483 6016
rect 18419 5956 18423 6012
rect 18423 5956 18479 6012
rect 18479 5956 18483 6012
rect 18419 5952 18483 5956
rect 18499 6012 18563 6016
rect 18499 5956 18503 6012
rect 18503 5956 18559 6012
rect 18559 5956 18563 6012
rect 18499 5952 18563 5956
rect 5896 5468 5960 5472
rect 5896 5412 5900 5468
rect 5900 5412 5956 5468
rect 5956 5412 5960 5468
rect 5896 5408 5960 5412
rect 5976 5468 6040 5472
rect 5976 5412 5980 5468
rect 5980 5412 6036 5468
rect 6036 5412 6040 5468
rect 5976 5408 6040 5412
rect 6056 5468 6120 5472
rect 6056 5412 6060 5468
rect 6060 5412 6116 5468
rect 6116 5412 6120 5468
rect 6056 5408 6120 5412
rect 6136 5468 6200 5472
rect 6136 5412 6140 5468
rect 6140 5412 6196 5468
rect 6196 5412 6200 5468
rect 6136 5408 6200 5412
rect 10841 5468 10905 5472
rect 10841 5412 10845 5468
rect 10845 5412 10901 5468
rect 10901 5412 10905 5468
rect 10841 5408 10905 5412
rect 10921 5468 10985 5472
rect 10921 5412 10925 5468
rect 10925 5412 10981 5468
rect 10981 5412 10985 5468
rect 10921 5408 10985 5412
rect 11001 5468 11065 5472
rect 11001 5412 11005 5468
rect 11005 5412 11061 5468
rect 11061 5412 11065 5468
rect 11001 5408 11065 5412
rect 11081 5468 11145 5472
rect 11081 5412 11085 5468
rect 11085 5412 11141 5468
rect 11141 5412 11145 5468
rect 11081 5408 11145 5412
rect 15786 5468 15850 5472
rect 15786 5412 15790 5468
rect 15790 5412 15846 5468
rect 15846 5412 15850 5468
rect 15786 5408 15850 5412
rect 15866 5468 15930 5472
rect 15866 5412 15870 5468
rect 15870 5412 15926 5468
rect 15926 5412 15930 5468
rect 15866 5408 15930 5412
rect 15946 5468 16010 5472
rect 15946 5412 15950 5468
rect 15950 5412 16006 5468
rect 16006 5412 16010 5468
rect 15946 5408 16010 5412
rect 16026 5468 16090 5472
rect 16026 5412 16030 5468
rect 16030 5412 16086 5468
rect 16086 5412 16090 5468
rect 16026 5408 16090 5412
rect 20731 5468 20795 5472
rect 20731 5412 20735 5468
rect 20735 5412 20791 5468
rect 20791 5412 20795 5468
rect 20731 5408 20795 5412
rect 20811 5468 20875 5472
rect 20811 5412 20815 5468
rect 20815 5412 20871 5468
rect 20871 5412 20875 5468
rect 20811 5408 20875 5412
rect 20891 5468 20955 5472
rect 20891 5412 20895 5468
rect 20895 5412 20951 5468
rect 20951 5412 20955 5468
rect 20891 5408 20955 5412
rect 20971 5468 21035 5472
rect 20971 5412 20975 5468
rect 20975 5412 21031 5468
rect 21031 5412 21035 5468
rect 20971 5408 21035 5412
rect 3424 4924 3488 4928
rect 3424 4868 3428 4924
rect 3428 4868 3484 4924
rect 3484 4868 3488 4924
rect 3424 4864 3488 4868
rect 3504 4924 3568 4928
rect 3504 4868 3508 4924
rect 3508 4868 3564 4924
rect 3564 4868 3568 4924
rect 3504 4864 3568 4868
rect 3584 4924 3648 4928
rect 3584 4868 3588 4924
rect 3588 4868 3644 4924
rect 3644 4868 3648 4924
rect 3584 4864 3648 4868
rect 3664 4924 3728 4928
rect 3664 4868 3668 4924
rect 3668 4868 3724 4924
rect 3724 4868 3728 4924
rect 3664 4864 3728 4868
rect 8369 4924 8433 4928
rect 8369 4868 8373 4924
rect 8373 4868 8429 4924
rect 8429 4868 8433 4924
rect 8369 4864 8433 4868
rect 8449 4924 8513 4928
rect 8449 4868 8453 4924
rect 8453 4868 8509 4924
rect 8509 4868 8513 4924
rect 8449 4864 8513 4868
rect 8529 4924 8593 4928
rect 8529 4868 8533 4924
rect 8533 4868 8589 4924
rect 8589 4868 8593 4924
rect 8529 4864 8593 4868
rect 8609 4924 8673 4928
rect 8609 4868 8613 4924
rect 8613 4868 8669 4924
rect 8669 4868 8673 4924
rect 8609 4864 8673 4868
rect 13314 4924 13378 4928
rect 13314 4868 13318 4924
rect 13318 4868 13374 4924
rect 13374 4868 13378 4924
rect 13314 4864 13378 4868
rect 13394 4924 13458 4928
rect 13394 4868 13398 4924
rect 13398 4868 13454 4924
rect 13454 4868 13458 4924
rect 13394 4864 13458 4868
rect 13474 4924 13538 4928
rect 13474 4868 13478 4924
rect 13478 4868 13534 4924
rect 13534 4868 13538 4924
rect 13474 4864 13538 4868
rect 13554 4924 13618 4928
rect 13554 4868 13558 4924
rect 13558 4868 13614 4924
rect 13614 4868 13618 4924
rect 13554 4864 13618 4868
rect 18259 4924 18323 4928
rect 18259 4868 18263 4924
rect 18263 4868 18319 4924
rect 18319 4868 18323 4924
rect 18259 4864 18323 4868
rect 18339 4924 18403 4928
rect 18339 4868 18343 4924
rect 18343 4868 18399 4924
rect 18399 4868 18403 4924
rect 18339 4864 18403 4868
rect 18419 4924 18483 4928
rect 18419 4868 18423 4924
rect 18423 4868 18479 4924
rect 18479 4868 18483 4924
rect 18419 4864 18483 4868
rect 18499 4924 18563 4928
rect 18499 4868 18503 4924
rect 18503 4868 18559 4924
rect 18559 4868 18563 4924
rect 18499 4864 18563 4868
rect 5896 4380 5960 4384
rect 5896 4324 5900 4380
rect 5900 4324 5956 4380
rect 5956 4324 5960 4380
rect 5896 4320 5960 4324
rect 5976 4380 6040 4384
rect 5976 4324 5980 4380
rect 5980 4324 6036 4380
rect 6036 4324 6040 4380
rect 5976 4320 6040 4324
rect 6056 4380 6120 4384
rect 6056 4324 6060 4380
rect 6060 4324 6116 4380
rect 6116 4324 6120 4380
rect 6056 4320 6120 4324
rect 6136 4380 6200 4384
rect 6136 4324 6140 4380
rect 6140 4324 6196 4380
rect 6196 4324 6200 4380
rect 6136 4320 6200 4324
rect 10841 4380 10905 4384
rect 10841 4324 10845 4380
rect 10845 4324 10901 4380
rect 10901 4324 10905 4380
rect 10841 4320 10905 4324
rect 10921 4380 10985 4384
rect 10921 4324 10925 4380
rect 10925 4324 10981 4380
rect 10981 4324 10985 4380
rect 10921 4320 10985 4324
rect 11001 4380 11065 4384
rect 11001 4324 11005 4380
rect 11005 4324 11061 4380
rect 11061 4324 11065 4380
rect 11001 4320 11065 4324
rect 11081 4380 11145 4384
rect 11081 4324 11085 4380
rect 11085 4324 11141 4380
rect 11141 4324 11145 4380
rect 11081 4320 11145 4324
rect 15786 4380 15850 4384
rect 15786 4324 15790 4380
rect 15790 4324 15846 4380
rect 15846 4324 15850 4380
rect 15786 4320 15850 4324
rect 15866 4380 15930 4384
rect 15866 4324 15870 4380
rect 15870 4324 15926 4380
rect 15926 4324 15930 4380
rect 15866 4320 15930 4324
rect 15946 4380 16010 4384
rect 15946 4324 15950 4380
rect 15950 4324 16006 4380
rect 16006 4324 16010 4380
rect 15946 4320 16010 4324
rect 16026 4380 16090 4384
rect 16026 4324 16030 4380
rect 16030 4324 16086 4380
rect 16086 4324 16090 4380
rect 16026 4320 16090 4324
rect 20731 4380 20795 4384
rect 20731 4324 20735 4380
rect 20735 4324 20791 4380
rect 20791 4324 20795 4380
rect 20731 4320 20795 4324
rect 20811 4380 20875 4384
rect 20811 4324 20815 4380
rect 20815 4324 20871 4380
rect 20871 4324 20875 4380
rect 20811 4320 20875 4324
rect 20891 4380 20955 4384
rect 20891 4324 20895 4380
rect 20895 4324 20951 4380
rect 20951 4324 20955 4380
rect 20891 4320 20955 4324
rect 20971 4380 21035 4384
rect 20971 4324 20975 4380
rect 20975 4324 21031 4380
rect 21031 4324 21035 4380
rect 20971 4320 21035 4324
rect 3424 3836 3488 3840
rect 3424 3780 3428 3836
rect 3428 3780 3484 3836
rect 3484 3780 3488 3836
rect 3424 3776 3488 3780
rect 3504 3836 3568 3840
rect 3504 3780 3508 3836
rect 3508 3780 3564 3836
rect 3564 3780 3568 3836
rect 3504 3776 3568 3780
rect 3584 3836 3648 3840
rect 3584 3780 3588 3836
rect 3588 3780 3644 3836
rect 3644 3780 3648 3836
rect 3584 3776 3648 3780
rect 3664 3836 3728 3840
rect 3664 3780 3668 3836
rect 3668 3780 3724 3836
rect 3724 3780 3728 3836
rect 3664 3776 3728 3780
rect 8369 3836 8433 3840
rect 8369 3780 8373 3836
rect 8373 3780 8429 3836
rect 8429 3780 8433 3836
rect 8369 3776 8433 3780
rect 8449 3836 8513 3840
rect 8449 3780 8453 3836
rect 8453 3780 8509 3836
rect 8509 3780 8513 3836
rect 8449 3776 8513 3780
rect 8529 3836 8593 3840
rect 8529 3780 8533 3836
rect 8533 3780 8589 3836
rect 8589 3780 8593 3836
rect 8529 3776 8593 3780
rect 8609 3836 8673 3840
rect 8609 3780 8613 3836
rect 8613 3780 8669 3836
rect 8669 3780 8673 3836
rect 8609 3776 8673 3780
rect 13314 3836 13378 3840
rect 13314 3780 13318 3836
rect 13318 3780 13374 3836
rect 13374 3780 13378 3836
rect 13314 3776 13378 3780
rect 13394 3836 13458 3840
rect 13394 3780 13398 3836
rect 13398 3780 13454 3836
rect 13454 3780 13458 3836
rect 13394 3776 13458 3780
rect 13474 3836 13538 3840
rect 13474 3780 13478 3836
rect 13478 3780 13534 3836
rect 13534 3780 13538 3836
rect 13474 3776 13538 3780
rect 13554 3836 13618 3840
rect 13554 3780 13558 3836
rect 13558 3780 13614 3836
rect 13614 3780 13618 3836
rect 13554 3776 13618 3780
rect 18259 3836 18323 3840
rect 18259 3780 18263 3836
rect 18263 3780 18319 3836
rect 18319 3780 18323 3836
rect 18259 3776 18323 3780
rect 18339 3836 18403 3840
rect 18339 3780 18343 3836
rect 18343 3780 18399 3836
rect 18399 3780 18403 3836
rect 18339 3776 18403 3780
rect 18419 3836 18483 3840
rect 18419 3780 18423 3836
rect 18423 3780 18479 3836
rect 18479 3780 18483 3836
rect 18419 3776 18483 3780
rect 18499 3836 18563 3840
rect 18499 3780 18503 3836
rect 18503 3780 18559 3836
rect 18559 3780 18563 3836
rect 18499 3776 18563 3780
rect 5896 3292 5960 3296
rect 5896 3236 5900 3292
rect 5900 3236 5956 3292
rect 5956 3236 5960 3292
rect 5896 3232 5960 3236
rect 5976 3292 6040 3296
rect 5976 3236 5980 3292
rect 5980 3236 6036 3292
rect 6036 3236 6040 3292
rect 5976 3232 6040 3236
rect 6056 3292 6120 3296
rect 6056 3236 6060 3292
rect 6060 3236 6116 3292
rect 6116 3236 6120 3292
rect 6056 3232 6120 3236
rect 6136 3292 6200 3296
rect 6136 3236 6140 3292
rect 6140 3236 6196 3292
rect 6196 3236 6200 3292
rect 6136 3232 6200 3236
rect 10841 3292 10905 3296
rect 10841 3236 10845 3292
rect 10845 3236 10901 3292
rect 10901 3236 10905 3292
rect 10841 3232 10905 3236
rect 10921 3292 10985 3296
rect 10921 3236 10925 3292
rect 10925 3236 10981 3292
rect 10981 3236 10985 3292
rect 10921 3232 10985 3236
rect 11001 3292 11065 3296
rect 11001 3236 11005 3292
rect 11005 3236 11061 3292
rect 11061 3236 11065 3292
rect 11001 3232 11065 3236
rect 11081 3292 11145 3296
rect 11081 3236 11085 3292
rect 11085 3236 11141 3292
rect 11141 3236 11145 3292
rect 11081 3232 11145 3236
rect 15786 3292 15850 3296
rect 15786 3236 15790 3292
rect 15790 3236 15846 3292
rect 15846 3236 15850 3292
rect 15786 3232 15850 3236
rect 15866 3292 15930 3296
rect 15866 3236 15870 3292
rect 15870 3236 15926 3292
rect 15926 3236 15930 3292
rect 15866 3232 15930 3236
rect 15946 3292 16010 3296
rect 15946 3236 15950 3292
rect 15950 3236 16006 3292
rect 16006 3236 16010 3292
rect 15946 3232 16010 3236
rect 16026 3292 16090 3296
rect 16026 3236 16030 3292
rect 16030 3236 16086 3292
rect 16086 3236 16090 3292
rect 16026 3232 16090 3236
rect 20731 3292 20795 3296
rect 20731 3236 20735 3292
rect 20735 3236 20791 3292
rect 20791 3236 20795 3292
rect 20731 3232 20795 3236
rect 20811 3292 20875 3296
rect 20811 3236 20815 3292
rect 20815 3236 20871 3292
rect 20871 3236 20875 3292
rect 20811 3232 20875 3236
rect 20891 3292 20955 3296
rect 20891 3236 20895 3292
rect 20895 3236 20951 3292
rect 20951 3236 20955 3292
rect 20891 3232 20955 3236
rect 20971 3292 21035 3296
rect 20971 3236 20975 3292
rect 20975 3236 21031 3292
rect 21031 3236 21035 3292
rect 20971 3232 21035 3236
rect 3424 2748 3488 2752
rect 3424 2692 3428 2748
rect 3428 2692 3484 2748
rect 3484 2692 3488 2748
rect 3424 2688 3488 2692
rect 3504 2748 3568 2752
rect 3504 2692 3508 2748
rect 3508 2692 3564 2748
rect 3564 2692 3568 2748
rect 3504 2688 3568 2692
rect 3584 2748 3648 2752
rect 3584 2692 3588 2748
rect 3588 2692 3644 2748
rect 3644 2692 3648 2748
rect 3584 2688 3648 2692
rect 3664 2748 3728 2752
rect 3664 2692 3668 2748
rect 3668 2692 3724 2748
rect 3724 2692 3728 2748
rect 3664 2688 3728 2692
rect 8369 2748 8433 2752
rect 8369 2692 8373 2748
rect 8373 2692 8429 2748
rect 8429 2692 8433 2748
rect 8369 2688 8433 2692
rect 8449 2748 8513 2752
rect 8449 2692 8453 2748
rect 8453 2692 8509 2748
rect 8509 2692 8513 2748
rect 8449 2688 8513 2692
rect 8529 2748 8593 2752
rect 8529 2692 8533 2748
rect 8533 2692 8589 2748
rect 8589 2692 8593 2748
rect 8529 2688 8593 2692
rect 8609 2748 8673 2752
rect 8609 2692 8613 2748
rect 8613 2692 8669 2748
rect 8669 2692 8673 2748
rect 8609 2688 8673 2692
rect 13314 2748 13378 2752
rect 13314 2692 13318 2748
rect 13318 2692 13374 2748
rect 13374 2692 13378 2748
rect 13314 2688 13378 2692
rect 13394 2748 13458 2752
rect 13394 2692 13398 2748
rect 13398 2692 13454 2748
rect 13454 2692 13458 2748
rect 13394 2688 13458 2692
rect 13474 2748 13538 2752
rect 13474 2692 13478 2748
rect 13478 2692 13534 2748
rect 13534 2692 13538 2748
rect 13474 2688 13538 2692
rect 13554 2748 13618 2752
rect 13554 2692 13558 2748
rect 13558 2692 13614 2748
rect 13614 2692 13618 2748
rect 13554 2688 13618 2692
rect 18259 2748 18323 2752
rect 18259 2692 18263 2748
rect 18263 2692 18319 2748
rect 18319 2692 18323 2748
rect 18259 2688 18323 2692
rect 18339 2748 18403 2752
rect 18339 2692 18343 2748
rect 18343 2692 18399 2748
rect 18399 2692 18403 2748
rect 18339 2688 18403 2692
rect 18419 2748 18483 2752
rect 18419 2692 18423 2748
rect 18423 2692 18479 2748
rect 18479 2692 18483 2748
rect 18419 2688 18483 2692
rect 18499 2748 18563 2752
rect 18499 2692 18503 2748
rect 18503 2692 18559 2748
rect 18559 2692 18563 2748
rect 18499 2688 18563 2692
rect 5896 2204 5960 2208
rect 5896 2148 5900 2204
rect 5900 2148 5956 2204
rect 5956 2148 5960 2204
rect 5896 2144 5960 2148
rect 5976 2204 6040 2208
rect 5976 2148 5980 2204
rect 5980 2148 6036 2204
rect 6036 2148 6040 2204
rect 5976 2144 6040 2148
rect 6056 2204 6120 2208
rect 6056 2148 6060 2204
rect 6060 2148 6116 2204
rect 6116 2148 6120 2204
rect 6056 2144 6120 2148
rect 6136 2204 6200 2208
rect 6136 2148 6140 2204
rect 6140 2148 6196 2204
rect 6196 2148 6200 2204
rect 6136 2144 6200 2148
rect 10841 2204 10905 2208
rect 10841 2148 10845 2204
rect 10845 2148 10901 2204
rect 10901 2148 10905 2204
rect 10841 2144 10905 2148
rect 10921 2204 10985 2208
rect 10921 2148 10925 2204
rect 10925 2148 10981 2204
rect 10981 2148 10985 2204
rect 10921 2144 10985 2148
rect 11001 2204 11065 2208
rect 11001 2148 11005 2204
rect 11005 2148 11061 2204
rect 11061 2148 11065 2204
rect 11001 2144 11065 2148
rect 11081 2204 11145 2208
rect 11081 2148 11085 2204
rect 11085 2148 11141 2204
rect 11141 2148 11145 2204
rect 11081 2144 11145 2148
rect 15786 2204 15850 2208
rect 15786 2148 15790 2204
rect 15790 2148 15846 2204
rect 15846 2148 15850 2204
rect 15786 2144 15850 2148
rect 15866 2204 15930 2208
rect 15866 2148 15870 2204
rect 15870 2148 15926 2204
rect 15926 2148 15930 2204
rect 15866 2144 15930 2148
rect 15946 2204 16010 2208
rect 15946 2148 15950 2204
rect 15950 2148 16006 2204
rect 16006 2148 16010 2204
rect 15946 2144 16010 2148
rect 16026 2204 16090 2208
rect 16026 2148 16030 2204
rect 16030 2148 16086 2204
rect 16086 2148 16090 2204
rect 16026 2144 16090 2148
rect 20731 2204 20795 2208
rect 20731 2148 20735 2204
rect 20735 2148 20791 2204
rect 20791 2148 20795 2204
rect 20731 2144 20795 2148
rect 20811 2204 20875 2208
rect 20811 2148 20815 2204
rect 20815 2148 20871 2204
rect 20871 2148 20875 2204
rect 20811 2144 20875 2148
rect 20891 2204 20955 2208
rect 20891 2148 20895 2204
rect 20895 2148 20951 2204
rect 20951 2148 20955 2204
rect 20891 2144 20955 2148
rect 20971 2204 21035 2208
rect 20971 2148 20975 2204
rect 20975 2148 21031 2204
rect 21031 2148 21035 2204
rect 20971 2144 21035 2148
<< metal4 >>
rect 3416 19072 3736 19632
rect 3416 19008 3424 19072
rect 3488 19008 3504 19072
rect 3568 19008 3584 19072
rect 3648 19008 3664 19072
rect 3728 19008 3736 19072
rect 3416 17984 3736 19008
rect 3416 17920 3424 17984
rect 3488 17920 3504 17984
rect 3568 17920 3584 17984
rect 3648 17920 3664 17984
rect 3728 17920 3736 17984
rect 3416 16896 3736 17920
rect 3416 16832 3424 16896
rect 3488 16832 3504 16896
rect 3568 16832 3584 16896
rect 3648 16832 3664 16896
rect 3728 16832 3736 16896
rect 3416 15808 3736 16832
rect 3416 15744 3424 15808
rect 3488 15744 3504 15808
rect 3568 15744 3584 15808
rect 3648 15744 3664 15808
rect 3728 15744 3736 15808
rect 3416 14720 3736 15744
rect 3416 14656 3424 14720
rect 3488 14656 3504 14720
rect 3568 14656 3584 14720
rect 3648 14656 3664 14720
rect 3728 14656 3736 14720
rect 3416 13632 3736 14656
rect 3416 13568 3424 13632
rect 3488 13568 3504 13632
rect 3568 13568 3584 13632
rect 3648 13568 3664 13632
rect 3728 13568 3736 13632
rect 3416 12544 3736 13568
rect 3416 12480 3424 12544
rect 3488 12480 3504 12544
rect 3568 12480 3584 12544
rect 3648 12480 3664 12544
rect 3728 12480 3736 12544
rect 3416 11456 3736 12480
rect 3416 11392 3424 11456
rect 3488 11392 3504 11456
rect 3568 11392 3584 11456
rect 3648 11392 3664 11456
rect 3728 11392 3736 11456
rect 3416 10368 3736 11392
rect 3416 10304 3424 10368
rect 3488 10304 3504 10368
rect 3568 10304 3584 10368
rect 3648 10304 3664 10368
rect 3728 10304 3736 10368
rect 3416 9280 3736 10304
rect 3416 9216 3424 9280
rect 3488 9216 3504 9280
rect 3568 9216 3584 9280
rect 3648 9216 3664 9280
rect 3728 9216 3736 9280
rect 3416 8192 3736 9216
rect 3416 8128 3424 8192
rect 3488 8128 3504 8192
rect 3568 8128 3584 8192
rect 3648 8128 3664 8192
rect 3728 8128 3736 8192
rect 3416 7104 3736 8128
rect 3416 7040 3424 7104
rect 3488 7040 3504 7104
rect 3568 7040 3584 7104
rect 3648 7040 3664 7104
rect 3728 7040 3736 7104
rect 3416 6016 3736 7040
rect 3416 5952 3424 6016
rect 3488 5952 3504 6016
rect 3568 5952 3584 6016
rect 3648 5952 3664 6016
rect 3728 5952 3736 6016
rect 3416 4928 3736 5952
rect 3416 4864 3424 4928
rect 3488 4864 3504 4928
rect 3568 4864 3584 4928
rect 3648 4864 3664 4928
rect 3728 4864 3736 4928
rect 3416 3840 3736 4864
rect 3416 3776 3424 3840
rect 3488 3776 3504 3840
rect 3568 3776 3584 3840
rect 3648 3776 3664 3840
rect 3728 3776 3736 3840
rect 3416 2752 3736 3776
rect 3416 2688 3424 2752
rect 3488 2688 3504 2752
rect 3568 2688 3584 2752
rect 3648 2688 3664 2752
rect 3728 2688 3736 2752
rect 3416 2128 3736 2688
rect 5888 19616 6208 19632
rect 5888 19552 5896 19616
rect 5960 19552 5976 19616
rect 6040 19552 6056 19616
rect 6120 19552 6136 19616
rect 6200 19552 6208 19616
rect 5888 18528 6208 19552
rect 5888 18464 5896 18528
rect 5960 18464 5976 18528
rect 6040 18464 6056 18528
rect 6120 18464 6136 18528
rect 6200 18464 6208 18528
rect 5888 17440 6208 18464
rect 5888 17376 5896 17440
rect 5960 17376 5976 17440
rect 6040 17376 6056 17440
rect 6120 17376 6136 17440
rect 6200 17376 6208 17440
rect 5888 16352 6208 17376
rect 5888 16288 5896 16352
rect 5960 16288 5976 16352
rect 6040 16288 6056 16352
rect 6120 16288 6136 16352
rect 6200 16288 6208 16352
rect 5888 15264 6208 16288
rect 5888 15200 5896 15264
rect 5960 15200 5976 15264
rect 6040 15200 6056 15264
rect 6120 15200 6136 15264
rect 6200 15200 6208 15264
rect 5888 14176 6208 15200
rect 5888 14112 5896 14176
rect 5960 14112 5976 14176
rect 6040 14112 6056 14176
rect 6120 14112 6136 14176
rect 6200 14112 6208 14176
rect 5888 13088 6208 14112
rect 5888 13024 5896 13088
rect 5960 13024 5976 13088
rect 6040 13024 6056 13088
rect 6120 13024 6136 13088
rect 6200 13024 6208 13088
rect 5888 12000 6208 13024
rect 5888 11936 5896 12000
rect 5960 11936 5976 12000
rect 6040 11936 6056 12000
rect 6120 11936 6136 12000
rect 6200 11936 6208 12000
rect 5888 10912 6208 11936
rect 5888 10848 5896 10912
rect 5960 10848 5976 10912
rect 6040 10848 6056 10912
rect 6120 10848 6136 10912
rect 6200 10848 6208 10912
rect 5888 9824 6208 10848
rect 5888 9760 5896 9824
rect 5960 9760 5976 9824
rect 6040 9760 6056 9824
rect 6120 9760 6136 9824
rect 6200 9760 6208 9824
rect 5888 8736 6208 9760
rect 5888 8672 5896 8736
rect 5960 8672 5976 8736
rect 6040 8672 6056 8736
rect 6120 8672 6136 8736
rect 6200 8672 6208 8736
rect 5888 7648 6208 8672
rect 5888 7584 5896 7648
rect 5960 7584 5976 7648
rect 6040 7584 6056 7648
rect 6120 7584 6136 7648
rect 6200 7584 6208 7648
rect 5888 6560 6208 7584
rect 5888 6496 5896 6560
rect 5960 6496 5976 6560
rect 6040 6496 6056 6560
rect 6120 6496 6136 6560
rect 6200 6496 6208 6560
rect 5888 5472 6208 6496
rect 5888 5408 5896 5472
rect 5960 5408 5976 5472
rect 6040 5408 6056 5472
rect 6120 5408 6136 5472
rect 6200 5408 6208 5472
rect 5888 4384 6208 5408
rect 5888 4320 5896 4384
rect 5960 4320 5976 4384
rect 6040 4320 6056 4384
rect 6120 4320 6136 4384
rect 6200 4320 6208 4384
rect 5888 3296 6208 4320
rect 5888 3232 5896 3296
rect 5960 3232 5976 3296
rect 6040 3232 6056 3296
rect 6120 3232 6136 3296
rect 6200 3232 6208 3296
rect 5888 2208 6208 3232
rect 5888 2144 5896 2208
rect 5960 2144 5976 2208
rect 6040 2144 6056 2208
rect 6120 2144 6136 2208
rect 6200 2144 6208 2208
rect 5888 2128 6208 2144
rect 8361 19072 8681 19632
rect 8361 19008 8369 19072
rect 8433 19008 8449 19072
rect 8513 19008 8529 19072
rect 8593 19008 8609 19072
rect 8673 19008 8681 19072
rect 8361 17984 8681 19008
rect 8361 17920 8369 17984
rect 8433 17920 8449 17984
rect 8513 17920 8529 17984
rect 8593 17920 8609 17984
rect 8673 17920 8681 17984
rect 8361 16896 8681 17920
rect 8361 16832 8369 16896
rect 8433 16832 8449 16896
rect 8513 16832 8529 16896
rect 8593 16832 8609 16896
rect 8673 16832 8681 16896
rect 8361 15808 8681 16832
rect 8361 15744 8369 15808
rect 8433 15744 8449 15808
rect 8513 15744 8529 15808
rect 8593 15744 8609 15808
rect 8673 15744 8681 15808
rect 8361 14720 8681 15744
rect 8361 14656 8369 14720
rect 8433 14656 8449 14720
rect 8513 14656 8529 14720
rect 8593 14656 8609 14720
rect 8673 14656 8681 14720
rect 8361 13632 8681 14656
rect 8361 13568 8369 13632
rect 8433 13568 8449 13632
rect 8513 13568 8529 13632
rect 8593 13568 8609 13632
rect 8673 13568 8681 13632
rect 8361 12544 8681 13568
rect 8361 12480 8369 12544
rect 8433 12480 8449 12544
rect 8513 12480 8529 12544
rect 8593 12480 8609 12544
rect 8673 12480 8681 12544
rect 8361 11456 8681 12480
rect 8361 11392 8369 11456
rect 8433 11392 8449 11456
rect 8513 11392 8529 11456
rect 8593 11392 8609 11456
rect 8673 11392 8681 11456
rect 8361 10368 8681 11392
rect 8361 10304 8369 10368
rect 8433 10304 8449 10368
rect 8513 10304 8529 10368
rect 8593 10304 8609 10368
rect 8673 10304 8681 10368
rect 8361 9280 8681 10304
rect 8361 9216 8369 9280
rect 8433 9216 8449 9280
rect 8513 9216 8529 9280
rect 8593 9216 8609 9280
rect 8673 9216 8681 9280
rect 8361 8192 8681 9216
rect 8361 8128 8369 8192
rect 8433 8128 8449 8192
rect 8513 8128 8529 8192
rect 8593 8128 8609 8192
rect 8673 8128 8681 8192
rect 8361 7104 8681 8128
rect 8361 7040 8369 7104
rect 8433 7040 8449 7104
rect 8513 7040 8529 7104
rect 8593 7040 8609 7104
rect 8673 7040 8681 7104
rect 8361 6016 8681 7040
rect 8361 5952 8369 6016
rect 8433 5952 8449 6016
rect 8513 5952 8529 6016
rect 8593 5952 8609 6016
rect 8673 5952 8681 6016
rect 8361 4928 8681 5952
rect 8361 4864 8369 4928
rect 8433 4864 8449 4928
rect 8513 4864 8529 4928
rect 8593 4864 8609 4928
rect 8673 4864 8681 4928
rect 8361 3840 8681 4864
rect 8361 3776 8369 3840
rect 8433 3776 8449 3840
rect 8513 3776 8529 3840
rect 8593 3776 8609 3840
rect 8673 3776 8681 3840
rect 8361 2752 8681 3776
rect 8361 2688 8369 2752
rect 8433 2688 8449 2752
rect 8513 2688 8529 2752
rect 8593 2688 8609 2752
rect 8673 2688 8681 2752
rect 8361 2128 8681 2688
rect 10833 19616 11153 19632
rect 10833 19552 10841 19616
rect 10905 19552 10921 19616
rect 10985 19552 11001 19616
rect 11065 19552 11081 19616
rect 11145 19552 11153 19616
rect 10833 18528 11153 19552
rect 10833 18464 10841 18528
rect 10905 18464 10921 18528
rect 10985 18464 11001 18528
rect 11065 18464 11081 18528
rect 11145 18464 11153 18528
rect 10833 17440 11153 18464
rect 10833 17376 10841 17440
rect 10905 17376 10921 17440
rect 10985 17376 11001 17440
rect 11065 17376 11081 17440
rect 11145 17376 11153 17440
rect 10833 16352 11153 17376
rect 10833 16288 10841 16352
rect 10905 16288 10921 16352
rect 10985 16288 11001 16352
rect 11065 16288 11081 16352
rect 11145 16288 11153 16352
rect 10833 15264 11153 16288
rect 10833 15200 10841 15264
rect 10905 15200 10921 15264
rect 10985 15200 11001 15264
rect 11065 15200 11081 15264
rect 11145 15200 11153 15264
rect 10833 14176 11153 15200
rect 10833 14112 10841 14176
rect 10905 14112 10921 14176
rect 10985 14112 11001 14176
rect 11065 14112 11081 14176
rect 11145 14112 11153 14176
rect 10833 13088 11153 14112
rect 10833 13024 10841 13088
rect 10905 13024 10921 13088
rect 10985 13024 11001 13088
rect 11065 13024 11081 13088
rect 11145 13024 11153 13088
rect 10833 12000 11153 13024
rect 10833 11936 10841 12000
rect 10905 11936 10921 12000
rect 10985 11936 11001 12000
rect 11065 11936 11081 12000
rect 11145 11936 11153 12000
rect 10833 10912 11153 11936
rect 10833 10848 10841 10912
rect 10905 10848 10921 10912
rect 10985 10848 11001 10912
rect 11065 10848 11081 10912
rect 11145 10848 11153 10912
rect 10833 9824 11153 10848
rect 10833 9760 10841 9824
rect 10905 9760 10921 9824
rect 10985 9760 11001 9824
rect 11065 9760 11081 9824
rect 11145 9760 11153 9824
rect 10833 8736 11153 9760
rect 10833 8672 10841 8736
rect 10905 8672 10921 8736
rect 10985 8672 11001 8736
rect 11065 8672 11081 8736
rect 11145 8672 11153 8736
rect 10833 7648 11153 8672
rect 10833 7584 10841 7648
rect 10905 7584 10921 7648
rect 10985 7584 11001 7648
rect 11065 7584 11081 7648
rect 11145 7584 11153 7648
rect 10833 6560 11153 7584
rect 10833 6496 10841 6560
rect 10905 6496 10921 6560
rect 10985 6496 11001 6560
rect 11065 6496 11081 6560
rect 11145 6496 11153 6560
rect 10833 5472 11153 6496
rect 10833 5408 10841 5472
rect 10905 5408 10921 5472
rect 10985 5408 11001 5472
rect 11065 5408 11081 5472
rect 11145 5408 11153 5472
rect 10833 4384 11153 5408
rect 10833 4320 10841 4384
rect 10905 4320 10921 4384
rect 10985 4320 11001 4384
rect 11065 4320 11081 4384
rect 11145 4320 11153 4384
rect 10833 3296 11153 4320
rect 10833 3232 10841 3296
rect 10905 3232 10921 3296
rect 10985 3232 11001 3296
rect 11065 3232 11081 3296
rect 11145 3232 11153 3296
rect 10833 2208 11153 3232
rect 10833 2144 10841 2208
rect 10905 2144 10921 2208
rect 10985 2144 11001 2208
rect 11065 2144 11081 2208
rect 11145 2144 11153 2208
rect 10833 2128 11153 2144
rect 13306 19072 13626 19632
rect 13306 19008 13314 19072
rect 13378 19008 13394 19072
rect 13458 19008 13474 19072
rect 13538 19008 13554 19072
rect 13618 19008 13626 19072
rect 13306 17984 13626 19008
rect 13306 17920 13314 17984
rect 13378 17920 13394 17984
rect 13458 17920 13474 17984
rect 13538 17920 13554 17984
rect 13618 17920 13626 17984
rect 13306 16896 13626 17920
rect 13306 16832 13314 16896
rect 13378 16832 13394 16896
rect 13458 16832 13474 16896
rect 13538 16832 13554 16896
rect 13618 16832 13626 16896
rect 13306 15808 13626 16832
rect 13306 15744 13314 15808
rect 13378 15744 13394 15808
rect 13458 15744 13474 15808
rect 13538 15744 13554 15808
rect 13618 15744 13626 15808
rect 13306 14720 13626 15744
rect 13306 14656 13314 14720
rect 13378 14656 13394 14720
rect 13458 14656 13474 14720
rect 13538 14656 13554 14720
rect 13618 14656 13626 14720
rect 13306 13632 13626 14656
rect 13306 13568 13314 13632
rect 13378 13568 13394 13632
rect 13458 13568 13474 13632
rect 13538 13568 13554 13632
rect 13618 13568 13626 13632
rect 13306 12544 13626 13568
rect 13306 12480 13314 12544
rect 13378 12480 13394 12544
rect 13458 12480 13474 12544
rect 13538 12480 13554 12544
rect 13618 12480 13626 12544
rect 13306 11456 13626 12480
rect 13306 11392 13314 11456
rect 13378 11392 13394 11456
rect 13458 11392 13474 11456
rect 13538 11392 13554 11456
rect 13618 11392 13626 11456
rect 13306 10368 13626 11392
rect 13306 10304 13314 10368
rect 13378 10304 13394 10368
rect 13458 10304 13474 10368
rect 13538 10304 13554 10368
rect 13618 10304 13626 10368
rect 13306 9280 13626 10304
rect 13306 9216 13314 9280
rect 13378 9216 13394 9280
rect 13458 9216 13474 9280
rect 13538 9216 13554 9280
rect 13618 9216 13626 9280
rect 13306 8192 13626 9216
rect 13306 8128 13314 8192
rect 13378 8128 13394 8192
rect 13458 8128 13474 8192
rect 13538 8128 13554 8192
rect 13618 8128 13626 8192
rect 13306 7104 13626 8128
rect 13306 7040 13314 7104
rect 13378 7040 13394 7104
rect 13458 7040 13474 7104
rect 13538 7040 13554 7104
rect 13618 7040 13626 7104
rect 13306 6016 13626 7040
rect 13306 5952 13314 6016
rect 13378 5952 13394 6016
rect 13458 5952 13474 6016
rect 13538 5952 13554 6016
rect 13618 5952 13626 6016
rect 13306 4928 13626 5952
rect 13306 4864 13314 4928
rect 13378 4864 13394 4928
rect 13458 4864 13474 4928
rect 13538 4864 13554 4928
rect 13618 4864 13626 4928
rect 13306 3840 13626 4864
rect 13306 3776 13314 3840
rect 13378 3776 13394 3840
rect 13458 3776 13474 3840
rect 13538 3776 13554 3840
rect 13618 3776 13626 3840
rect 13306 2752 13626 3776
rect 13306 2688 13314 2752
rect 13378 2688 13394 2752
rect 13458 2688 13474 2752
rect 13538 2688 13554 2752
rect 13618 2688 13626 2752
rect 13306 2128 13626 2688
rect 15778 19616 16098 19632
rect 15778 19552 15786 19616
rect 15850 19552 15866 19616
rect 15930 19552 15946 19616
rect 16010 19552 16026 19616
rect 16090 19552 16098 19616
rect 15778 18528 16098 19552
rect 15778 18464 15786 18528
rect 15850 18464 15866 18528
rect 15930 18464 15946 18528
rect 16010 18464 16026 18528
rect 16090 18464 16098 18528
rect 15778 17440 16098 18464
rect 15778 17376 15786 17440
rect 15850 17376 15866 17440
rect 15930 17376 15946 17440
rect 16010 17376 16026 17440
rect 16090 17376 16098 17440
rect 15778 16352 16098 17376
rect 15778 16288 15786 16352
rect 15850 16288 15866 16352
rect 15930 16288 15946 16352
rect 16010 16288 16026 16352
rect 16090 16288 16098 16352
rect 15778 15264 16098 16288
rect 15778 15200 15786 15264
rect 15850 15200 15866 15264
rect 15930 15200 15946 15264
rect 16010 15200 16026 15264
rect 16090 15200 16098 15264
rect 15778 14176 16098 15200
rect 15778 14112 15786 14176
rect 15850 14112 15866 14176
rect 15930 14112 15946 14176
rect 16010 14112 16026 14176
rect 16090 14112 16098 14176
rect 15778 13088 16098 14112
rect 15778 13024 15786 13088
rect 15850 13024 15866 13088
rect 15930 13024 15946 13088
rect 16010 13024 16026 13088
rect 16090 13024 16098 13088
rect 15778 12000 16098 13024
rect 15778 11936 15786 12000
rect 15850 11936 15866 12000
rect 15930 11936 15946 12000
rect 16010 11936 16026 12000
rect 16090 11936 16098 12000
rect 15778 10912 16098 11936
rect 15778 10848 15786 10912
rect 15850 10848 15866 10912
rect 15930 10848 15946 10912
rect 16010 10848 16026 10912
rect 16090 10848 16098 10912
rect 15778 9824 16098 10848
rect 15778 9760 15786 9824
rect 15850 9760 15866 9824
rect 15930 9760 15946 9824
rect 16010 9760 16026 9824
rect 16090 9760 16098 9824
rect 15778 8736 16098 9760
rect 15778 8672 15786 8736
rect 15850 8672 15866 8736
rect 15930 8672 15946 8736
rect 16010 8672 16026 8736
rect 16090 8672 16098 8736
rect 15778 7648 16098 8672
rect 15778 7584 15786 7648
rect 15850 7584 15866 7648
rect 15930 7584 15946 7648
rect 16010 7584 16026 7648
rect 16090 7584 16098 7648
rect 15778 6560 16098 7584
rect 15778 6496 15786 6560
rect 15850 6496 15866 6560
rect 15930 6496 15946 6560
rect 16010 6496 16026 6560
rect 16090 6496 16098 6560
rect 15778 5472 16098 6496
rect 15778 5408 15786 5472
rect 15850 5408 15866 5472
rect 15930 5408 15946 5472
rect 16010 5408 16026 5472
rect 16090 5408 16098 5472
rect 15778 4384 16098 5408
rect 15778 4320 15786 4384
rect 15850 4320 15866 4384
rect 15930 4320 15946 4384
rect 16010 4320 16026 4384
rect 16090 4320 16098 4384
rect 15778 3296 16098 4320
rect 15778 3232 15786 3296
rect 15850 3232 15866 3296
rect 15930 3232 15946 3296
rect 16010 3232 16026 3296
rect 16090 3232 16098 3296
rect 15778 2208 16098 3232
rect 15778 2144 15786 2208
rect 15850 2144 15866 2208
rect 15930 2144 15946 2208
rect 16010 2144 16026 2208
rect 16090 2144 16098 2208
rect 15778 2128 16098 2144
rect 18251 19072 18571 19632
rect 18251 19008 18259 19072
rect 18323 19008 18339 19072
rect 18403 19008 18419 19072
rect 18483 19008 18499 19072
rect 18563 19008 18571 19072
rect 18251 17984 18571 19008
rect 18251 17920 18259 17984
rect 18323 17920 18339 17984
rect 18403 17920 18419 17984
rect 18483 17920 18499 17984
rect 18563 17920 18571 17984
rect 18251 16896 18571 17920
rect 18251 16832 18259 16896
rect 18323 16832 18339 16896
rect 18403 16832 18419 16896
rect 18483 16832 18499 16896
rect 18563 16832 18571 16896
rect 18251 15808 18571 16832
rect 18251 15744 18259 15808
rect 18323 15744 18339 15808
rect 18403 15744 18419 15808
rect 18483 15744 18499 15808
rect 18563 15744 18571 15808
rect 18251 14720 18571 15744
rect 18251 14656 18259 14720
rect 18323 14656 18339 14720
rect 18403 14656 18419 14720
rect 18483 14656 18499 14720
rect 18563 14656 18571 14720
rect 18251 13632 18571 14656
rect 18251 13568 18259 13632
rect 18323 13568 18339 13632
rect 18403 13568 18419 13632
rect 18483 13568 18499 13632
rect 18563 13568 18571 13632
rect 18251 12544 18571 13568
rect 18251 12480 18259 12544
rect 18323 12480 18339 12544
rect 18403 12480 18419 12544
rect 18483 12480 18499 12544
rect 18563 12480 18571 12544
rect 18251 11456 18571 12480
rect 18251 11392 18259 11456
rect 18323 11392 18339 11456
rect 18403 11392 18419 11456
rect 18483 11392 18499 11456
rect 18563 11392 18571 11456
rect 18251 10368 18571 11392
rect 18251 10304 18259 10368
rect 18323 10304 18339 10368
rect 18403 10304 18419 10368
rect 18483 10304 18499 10368
rect 18563 10304 18571 10368
rect 18251 9280 18571 10304
rect 18251 9216 18259 9280
rect 18323 9216 18339 9280
rect 18403 9216 18419 9280
rect 18483 9216 18499 9280
rect 18563 9216 18571 9280
rect 18251 8192 18571 9216
rect 18251 8128 18259 8192
rect 18323 8128 18339 8192
rect 18403 8128 18419 8192
rect 18483 8128 18499 8192
rect 18563 8128 18571 8192
rect 18251 7104 18571 8128
rect 18251 7040 18259 7104
rect 18323 7040 18339 7104
rect 18403 7040 18419 7104
rect 18483 7040 18499 7104
rect 18563 7040 18571 7104
rect 18251 6016 18571 7040
rect 18251 5952 18259 6016
rect 18323 5952 18339 6016
rect 18403 5952 18419 6016
rect 18483 5952 18499 6016
rect 18563 5952 18571 6016
rect 18251 4928 18571 5952
rect 18251 4864 18259 4928
rect 18323 4864 18339 4928
rect 18403 4864 18419 4928
rect 18483 4864 18499 4928
rect 18563 4864 18571 4928
rect 18251 3840 18571 4864
rect 18251 3776 18259 3840
rect 18323 3776 18339 3840
rect 18403 3776 18419 3840
rect 18483 3776 18499 3840
rect 18563 3776 18571 3840
rect 18251 2752 18571 3776
rect 18251 2688 18259 2752
rect 18323 2688 18339 2752
rect 18403 2688 18419 2752
rect 18483 2688 18499 2752
rect 18563 2688 18571 2752
rect 18251 2128 18571 2688
rect 20723 19616 21043 19632
rect 20723 19552 20731 19616
rect 20795 19552 20811 19616
rect 20875 19552 20891 19616
rect 20955 19552 20971 19616
rect 21035 19552 21043 19616
rect 20723 18528 21043 19552
rect 20723 18464 20731 18528
rect 20795 18464 20811 18528
rect 20875 18464 20891 18528
rect 20955 18464 20971 18528
rect 21035 18464 21043 18528
rect 20723 17440 21043 18464
rect 20723 17376 20731 17440
rect 20795 17376 20811 17440
rect 20875 17376 20891 17440
rect 20955 17376 20971 17440
rect 21035 17376 21043 17440
rect 20723 16352 21043 17376
rect 20723 16288 20731 16352
rect 20795 16288 20811 16352
rect 20875 16288 20891 16352
rect 20955 16288 20971 16352
rect 21035 16288 21043 16352
rect 20723 15264 21043 16288
rect 20723 15200 20731 15264
rect 20795 15200 20811 15264
rect 20875 15200 20891 15264
rect 20955 15200 20971 15264
rect 21035 15200 21043 15264
rect 20723 14176 21043 15200
rect 20723 14112 20731 14176
rect 20795 14112 20811 14176
rect 20875 14112 20891 14176
rect 20955 14112 20971 14176
rect 21035 14112 21043 14176
rect 20723 13088 21043 14112
rect 20723 13024 20731 13088
rect 20795 13024 20811 13088
rect 20875 13024 20891 13088
rect 20955 13024 20971 13088
rect 21035 13024 21043 13088
rect 20723 12000 21043 13024
rect 20723 11936 20731 12000
rect 20795 11936 20811 12000
rect 20875 11936 20891 12000
rect 20955 11936 20971 12000
rect 21035 11936 21043 12000
rect 20723 10912 21043 11936
rect 20723 10848 20731 10912
rect 20795 10848 20811 10912
rect 20875 10848 20891 10912
rect 20955 10848 20971 10912
rect 21035 10848 21043 10912
rect 20723 9824 21043 10848
rect 20723 9760 20731 9824
rect 20795 9760 20811 9824
rect 20875 9760 20891 9824
rect 20955 9760 20971 9824
rect 21035 9760 21043 9824
rect 20723 8736 21043 9760
rect 20723 8672 20731 8736
rect 20795 8672 20811 8736
rect 20875 8672 20891 8736
rect 20955 8672 20971 8736
rect 21035 8672 21043 8736
rect 20723 7648 21043 8672
rect 20723 7584 20731 7648
rect 20795 7584 20811 7648
rect 20875 7584 20891 7648
rect 20955 7584 20971 7648
rect 21035 7584 21043 7648
rect 20723 6560 21043 7584
rect 20723 6496 20731 6560
rect 20795 6496 20811 6560
rect 20875 6496 20891 6560
rect 20955 6496 20971 6560
rect 21035 6496 21043 6560
rect 20723 5472 21043 6496
rect 20723 5408 20731 5472
rect 20795 5408 20811 5472
rect 20875 5408 20891 5472
rect 20955 5408 20971 5472
rect 21035 5408 21043 5472
rect 20723 4384 21043 5408
rect 20723 4320 20731 4384
rect 20795 4320 20811 4384
rect 20875 4320 20891 4384
rect 20955 4320 20971 4384
rect 21035 4320 21043 4384
rect 20723 3296 21043 4320
rect 20723 3232 20731 3296
rect 20795 3232 20811 3296
rect 20875 3232 20891 3296
rect 20955 3232 20971 3296
rect 21035 3232 21043 3296
rect 20723 2208 21043 3232
rect 20723 2144 20731 2208
rect 20795 2144 20811 2208
rect 20875 2144 20891 2208
rect 20955 2144 20971 2208
rect 21035 2144 21043 2208
rect 20723 2128 21043 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2576 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1676037725
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74
timestamp 1676037725
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91
timestamp 1676037725
transform 1 0 9476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1676037725
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121
timestamp 1676037725
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133
timestamp 1676037725
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1676037725
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155
timestamp 1676037725
transform 1 0 15364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_10
timestamp 1676037725
transform 1 0 2024 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_36
timestamp 1676037725
transform 1 0 4416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_44
timestamp 1676037725
transform 1 0 5152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_68
timestamp 1676037725
transform 1 0 7360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_72
timestamp 1676037725
transform 1 0 7728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_103
timestamp 1676037725
transform 1 0 10580 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1676037725
transform 1 0 12236 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_128
timestamp 1676037725
transform 1 0 12880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_144
timestamp 1676037725
transform 1 0 14352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1676037725
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1676037725
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_178
timestamp 1676037725
transform 1 0 17480 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_190
timestamp 1676037725
transform 1 0 18584 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_202
timestamp 1676037725
transform 1 0 19688 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_210
timestamp 1676037725
transform 1 0 20424 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_9
timestamp 1676037725
transform 1 0 1932 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_61
timestamp 1676037725
transform 1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1676037725
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_115
timestamp 1676037725
transform 1 0 11684 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_120
timestamp 1676037725
transform 1 0 12144 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_128
timestamp 1676037725
transform 1 0 12880 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1676037725
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_151
timestamp 1676037725
transform 1 0 14996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_163
timestamp 1676037725
transform 1 0 16100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_169
timestamp 1676037725
transform 1 0 16652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_188
timestamp 1676037725
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_22
timestamp 1676037725
transform 1 0 3128 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_34
timestamp 1676037725
transform 1 0 4232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1676037725
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_89
timestamp 1676037725
transform 1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1676037725
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_141
timestamp 1676037725
transform 1 0 14076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_152
timestamp 1676037725
transform 1 0 15088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1676037725
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_179
timestamp 1676037725
transform 1 0 17572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_191
timestamp 1676037725
transform 1 0 18676 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_203
timestamp 1676037725
transform 1 0 19780 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_211
timestamp 1676037725
transform 1 0 20516 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_9
timestamp 1676037725
transform 1 0 1932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1676037725
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_61
timestamp 1676037725
transform 1 0 6716 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1676037725
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1676037725
transform 1 0 9660 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_110
timestamp 1676037725
transform 1 0 11224 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_122
timestamp 1676037725
transform 1 0 12328 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_134
timestamp 1676037725
transform 1 0 13432 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1676037725
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_160
timestamp 1676037725
transform 1 0 15824 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_180
timestamp 1676037725
transform 1 0 17664 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_187
timestamp 1676037725
transform 1 0 18308 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_11
timestamp 1676037725
transform 1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_16
timestamp 1676037725
transform 1 0 2576 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_34
timestamp 1676037725
transform 1 0 4232 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1676037725
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1676037725
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_121
timestamp 1676037725
transform 1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_133
timestamp 1676037725
transform 1 0 13340 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_146
timestamp 1676037725
transform 1 0 14536 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_158
timestamp 1676037725
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_175
timestamp 1676037725
transform 1 0 17204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_187
timestamp 1676037725
transform 1 0 18308 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_199
timestamp 1676037725
transform 1 0 19412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_211
timestamp 1676037725
transform 1 0 20516 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1676037725
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_45
timestamp 1676037725
transform 1 0 5244 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_62
timestamp 1676037725
transform 1 0 6808 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_74
timestamp 1676037725
transform 1 0 7912 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1676037725
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_93
timestamp 1676037725
transform 1 0 9660 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_110
timestamp 1676037725
transform 1 0 11224 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_122
timestamp 1676037725
transform 1 0 12328 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_134
timestamp 1676037725
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_148
timestamp 1676037725
transform 1 0 14720 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_160
timestamp 1676037725
transform 1 0 15824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_172
timestamp 1676037725
transform 1 0 16928 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_179
timestamp 1676037725
transform 1 0 17572 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_191
timestamp 1676037725
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_204
timestamp 1676037725
transform 1 0 19872 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_35
timestamp 1676037725
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1676037725
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_101
timestamp 1676037725
transform 1 0 10396 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1676037725
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_121
timestamp 1676037725
transform 1 0 12236 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_133
timestamp 1676037725
transform 1 0 13340 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_150
timestamp 1676037725
transform 1 0 14904 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_158
timestamp 1676037725
transform 1 0 15640 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1676037725
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_195
timestamp 1676037725
transform 1 0 19044 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_207
timestamp 1676037725
transform 1 0 20148 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_211
timestamp 1676037725
transform 1 0 20516 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_21
timestamp 1676037725
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_73
timestamp 1676037725
transform 1 0 7820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1676037725
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_93
timestamp 1676037725
transform 1 0 9660 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_110
timestamp 1676037725
transform 1 0 11224 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_122
timestamp 1676037725
transform 1 0 12328 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_130
timestamp 1676037725
transform 1 0 13064 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_151
timestamp 1676037725
transform 1 0 14996 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_155
timestamp 1676037725
transform 1 0 15364 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_163
timestamp 1676037725
transform 1 0 16100 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_171
timestamp 1676037725
transform 1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_181
timestamp 1676037725
transform 1 0 17756 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_185
timestamp 1676037725
transform 1 0 18124 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1676037725
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_36
timestamp 1676037725
transform 1 0 4416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_48
timestamp 1676037725
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_134
timestamp 1676037725
transform 1 0 13432 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_146
timestamp 1676037725
transform 1 0 14536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_158
timestamp 1676037725
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1676037725
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_177
timestamp 1676037725
transform 1 0 17388 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_183
timestamp 1676037725
transform 1 0 17940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_195
timestamp 1676037725
transform 1 0 19044 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_207
timestamp 1676037725
transform 1 0 20148 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_211
timestamp 1676037725
transform 1 0 20516 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_37
timestamp 1676037725
transform 1 0 4508 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_56
timestamp 1676037725
transform 1 0 6256 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp 1676037725
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_93
timestamp 1676037725
transform 1 0 9660 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_112
timestamp 1676037725
transform 1 0 11408 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_124
timestamp 1676037725
transform 1 0 12512 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 1676037725
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_160
timestamp 1676037725
transform 1 0 15824 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_168
timestamp 1676037725
transform 1 0 16560 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_174
timestamp 1676037725
transform 1 0 17112 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_181
timestamp 1676037725
transform 1 0 17756 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_202
timestamp 1676037725
transform 1 0 19688 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_210
timestamp 1676037725
transform 1 0 20424 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_19
timestamp 1676037725
transform 1 0 2852 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_36
timestamp 1676037725
transform 1 0 4416 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_48
timestamp 1676037725
transform 1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_134
timestamp 1676037725
transform 1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_146
timestamp 1676037725
transform 1 0 14536 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_158
timestamp 1676037725
transform 1 0 15640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_176
timestamp 1676037725
transform 1 0 17296 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1676037725
transform 1 0 18032 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_194
timestamp 1676037725
transform 1 0 18952 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_206
timestamp 1676037725
transform 1 0 20056 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1676037725
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_37
timestamp 1676037725
transform 1 0 4508 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_54
timestamp 1676037725
transform 1 0 6072 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_62
timestamp 1676037725
transform 1 0 6808 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1676037725
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_117
timestamp 1676037725
transform 1 0 11868 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_129
timestamp 1676037725
transform 1 0 12972 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1676037725
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_149
timestamp 1676037725
transform 1 0 14812 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_161
timestamp 1676037725
transform 1 0 15916 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_167
timestamp 1676037725
transform 1 0 16468 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_184
timestamp 1676037725
transform 1 0 18032 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_205
timestamp 1676037725
transform 1 0 19964 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_211
timestamp 1676037725
transform 1 0 20516 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_35
timestamp 1676037725
transform 1 0 4324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1676037725
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_91
timestamp 1676037725
transform 1 0 9476 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_103
timestamp 1676037725
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_132
timestamp 1676037725
transform 1 0 13248 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_140
timestamp 1676037725
transform 1 0 13984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_146
timestamp 1676037725
transform 1 0 14536 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_157
timestamp 1676037725
transform 1 0 15548 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_175
timestamp 1676037725
transform 1 0 17204 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_187
timestamp 1676037725
transform 1 0 18308 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_210
timestamp 1676037725
transform 1 0 20424 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1676037725
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_60
timestamp 1676037725
transform 1 0 6624 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1676037725
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_116
timestamp 1676037725
transform 1 0 11776 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_124
timestamp 1676037725
transform 1 0 12512 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_150
timestamp 1676037725
transform 1 0 14904 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_154
timestamp 1676037725
transform 1 0 15272 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_163
timestamp 1676037725
transform 1 0 16100 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_172
timestamp 1676037725
transform 1 0 16928 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_176
timestamp 1676037725
transform 1 0 17296 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1676037725
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_204
timestamp 1676037725
transform 1 0 19872 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_9
timestamp 1676037725
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_21
timestamp 1676037725
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_33
timestamp 1676037725
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1676037725
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1676037725
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_89
timestamp 1676037725
transform 1 0 9292 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1676037725
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_143
timestamp 1676037725
transform 1 0 14260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_155
timestamp 1676037725
transform 1 0 15364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_174
timestamp 1676037725
transform 1 0 17112 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_186
timestamp 1676037725
transform 1 0 18216 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_195
timestamp 1676037725
transform 1 0 19044 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_206
timestamp 1676037725
transform 1 0 20056 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1676037725
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_12
timestamp 1676037725
transform 1 0 2208 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1676037725
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_37
timestamp 1676037725
transform 1 0 4508 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_49
timestamp 1676037725
transform 1 0 5612 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_70
timestamp 1676037725
transform 1 0 7544 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1676037725
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_125
timestamp 1676037725
transform 1 0 12604 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_150
timestamp 1676037725
transform 1 0 14904 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_158
timestamp 1676037725
transform 1 0 15640 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_182
timestamp 1676037725
transform 1 0 17848 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_208
timestamp 1676037725
transform 1 0 20240 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1676037725
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_33
timestamp 1676037725
transform 1 0 4140 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_41
timestamp 1676037725
transform 1 0 4876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_74
timestamp 1676037725
transform 1 0 7912 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_82
timestamp 1676037725
transform 1 0 8648 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_91
timestamp 1676037725
transform 1 0 9476 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_99
timestamp 1676037725
transform 1 0 10212 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1676037725
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_124
timestamp 1676037725
transform 1 0 12512 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_132
timestamp 1676037725
transform 1 0 13248 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_144
timestamp 1676037725
transform 1 0 14352 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_150
timestamp 1676037725
transform 1 0 14904 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_154
timestamp 1676037725
transform 1 0 15272 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_175
timestamp 1676037725
transform 1 0 17204 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_182
timestamp 1676037725
transform 1 0 17848 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_199
timestamp 1676037725
transform 1 0 19412 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_210
timestamp 1676037725
transform 1 0 20424 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1676037725
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_17
timestamp 1676037725
transform 1 0 2668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1676037725
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_37
timestamp 1676037725
transform 1 0 4508 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_49
timestamp 1676037725
transform 1 0 5612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_74
timestamp 1676037725
transform 1 0 7912 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1676037725
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_95
timestamp 1676037725
transform 1 0 9844 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1676037725
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_123
timestamp 1676037725
transform 1 0 12420 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_129
timestamp 1676037725
transform 1 0 12972 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1676037725
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_151
timestamp 1676037725
transform 1 0 14996 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_158
timestamp 1676037725
transform 1 0 15640 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_162
timestamp 1676037725
transform 1 0 16008 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_170
timestamp 1676037725
transform 1 0 16744 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_178
timestamp 1676037725
transform 1 0 17480 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_187
timestamp 1676037725
transform 1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_201
timestamp 1676037725
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_208
timestamp 1676037725
transform 1 0 20240 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_11
timestamp 1676037725
transform 1 0 2116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_23
timestamp 1676037725
transform 1 0 3220 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_37
timestamp 1676037725
transform 1 0 4508 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1676037725
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_68
timestamp 1676037725
transform 1 0 7360 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_80
timestamp 1676037725
transform 1 0 8464 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_90
timestamp 1676037725
transform 1 0 9384 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_102
timestamp 1676037725
transform 1 0 10488 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_119
timestamp 1676037725
transform 1 0 12052 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_131
timestamp 1676037725
transform 1 0 13156 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_139
timestamp 1676037725
transform 1 0 13892 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_151
timestamp 1676037725
transform 1 0 14996 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1676037725
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_178
timestamp 1676037725
transform 1 0 17480 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_186
timestamp 1676037725
transform 1 0 18216 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_192
timestamp 1676037725
transform 1 0 18768 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_200
timestamp 1676037725
transform 1 0 19504 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_208
timestamp 1676037725
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_18
timestamp 1676037725
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1676037725
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_33
timestamp 1676037725
transform 1 0 4140 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_43
timestamp 1676037725
transform 1 0 5060 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_55
timestamp 1676037725
transform 1 0 6164 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_67
timestamp 1676037725
transform 1 0 7268 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_72
timestamp 1676037725
transform 1 0 7728 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_90
timestamp 1676037725
transform 1 0 9384 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_102
timestamp 1676037725
transform 1 0 10488 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_115
timestamp 1676037725
transform 1 0 11684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_127
timestamp 1676037725
transform 1 0 12788 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1676037725
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_146
timestamp 1676037725
transform 1 0 14536 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_158
timestamp 1676037725
transform 1 0 15640 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_170
timestamp 1676037725
transform 1 0 16744 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_186
timestamp 1676037725
transform 1 0 18216 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_203
timestamp 1676037725
transform 1 0 19780 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_207
timestamp 1676037725
transform 1 0 20148 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_211
timestamp 1676037725
transform 1 0 20516 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_14
timestamp 1676037725
transform 1 0 2392 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_18
timestamp 1676037725
transform 1 0 2760 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_23
timestamp 1676037725
transform 1 0 3220 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_35
timestamp 1676037725
transform 1 0 4324 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_41
timestamp 1676037725
transform 1 0 4876 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1676037725
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_68
timestamp 1676037725
transform 1 0 7360 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_77
timestamp 1676037725
transform 1 0 8188 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_90
timestamp 1676037725
transform 1 0 9384 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_94
timestamp 1676037725
transform 1 0 9752 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_102
timestamp 1676037725
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_124
timestamp 1676037725
transform 1 0 12512 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_132
timestamp 1676037725
transform 1 0 13248 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1676037725
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_177
timestamp 1676037725
transform 1 0 17388 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_192
timestamp 1676037725
transform 1 0 18768 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_198
timestamp 1676037725
transform 1 0 19320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_207
timestamp 1676037725
transform 1 0 20148 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_211
timestamp 1676037725
transform 1 0 20516 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_14
timestamp 1676037725
transform 1 0 2392 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1676037725
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_38
timestamp 1676037725
transform 1 0 4600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_49
timestamp 1676037725
transform 1 0 5612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1676037725
transform 1 0 6256 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_62
timestamp 1676037725
transform 1 0 6808 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_71
timestamp 1676037725
transform 1 0 7636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1676037725
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_95
timestamp 1676037725
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_107
timestamp 1676037725
transform 1 0 10948 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_124
timestamp 1676037725
transform 1 0 12512 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_130
timestamp 1676037725
transform 1 0 13064 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1676037725
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1676037725
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_170
timestamp 1676037725
transform 1 0 16744 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_182
timestamp 1676037725
transform 1 0 17848 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_190
timestamp 1676037725
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_11
timestamp 1676037725
transform 1 0 2116 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_16
timestamp 1676037725
transform 1 0 2576 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_28
timestamp 1676037725
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_40
timestamp 1676037725
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1676037725
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_70
timestamp 1676037725
transform 1 0 7544 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_78
timestamp 1676037725
transform 1 0 8280 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_90
timestamp 1676037725
transform 1 0 9384 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_102
timestamp 1676037725
transform 1 0 10488 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_122
timestamp 1676037725
transform 1 0 12328 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_126
timestamp 1676037725
transform 1 0 12696 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_136
timestamp 1676037725
transform 1 0 13616 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_144
timestamp 1676037725
transform 1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_157
timestamp 1676037725
transform 1 0 15548 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1676037725
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_177
timestamp 1676037725
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_187
timestamp 1676037725
transform 1 0 18308 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_195
timestamp 1676037725
transform 1 0 19044 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_207
timestamp 1676037725
transform 1 0 20148 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_211
timestamp 1676037725
transform 1 0 20516 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_18
timestamp 1676037725
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1676037725
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_74
timestamp 1676037725
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1676037725
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_92
timestamp 1676037725
transform 1 0 9568 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_100
timestamp 1676037725
transform 1 0 10304 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_108
timestamp 1676037725
transform 1 0 11040 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_115
timestamp 1676037725
transform 1 0 11684 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_123
timestamp 1676037725
transform 1 0 12420 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_128
timestamp 1676037725
transform 1 0 12880 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1676037725
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_148
timestamp 1676037725
transform 1 0 14720 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_160
timestamp 1676037725
transform 1 0 15824 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_169
timestamp 1676037725
transform 1 0 16652 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_181
timestamp 1676037725
transform 1 0 17756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1676037725
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_32
timestamp 1676037725
transform 1 0 4048 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_43
timestamp 1676037725
transform 1 0 5060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_50
timestamp 1676037725
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_63
timestamp 1676037725
transform 1 0 6900 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_75
timestamp 1676037725
transform 1 0 8004 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_95
timestamp 1676037725
transform 1 0 9844 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_106
timestamp 1676037725
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_124
timestamp 1676037725
transform 1 0 12512 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp 1676037725
transform 1 0 13524 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_143
timestamp 1676037725
transform 1 0 14260 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_154
timestamp 1676037725
transform 1 0 15272 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1676037725
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_205
timestamp 1676037725
transform 1 0 19964 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_211
timestamp 1676037725
transform 1 0 20516 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1676037725
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_37
timestamp 1676037725
transform 1 0 4508 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_43
timestamp 1676037725
transform 1 0 5060 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_51
timestamp 1676037725
transform 1 0 5796 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_59
timestamp 1676037725
transform 1 0 6532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_73
timestamp 1676037725
transform 1 0 7820 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_105
timestamp 1676037725
transform 1 0 10764 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_113
timestamp 1676037725
transform 1 0 11500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_125
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1676037725
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_147
timestamp 1676037725
transform 1 0 14628 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_151
timestamp 1676037725
transform 1 0 14996 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_163
timestamp 1676037725
transform 1 0 16100 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_175
timestamp 1676037725
transform 1 0 17204 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_187
timestamp 1676037725
transform 1 0 18308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_62
timestamp 1676037725
transform 1 0 6808 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_70
timestamp 1676037725
transform 1 0 7544 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_75
timestamp 1676037725
transform 1 0 8004 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_87
timestamp 1676037725
transform 1 0 9108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_99
timestamp 1676037725
transform 1 0 10212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1676037725
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_205
timestamp 1676037725
transform 1 0 19964 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_211
timestamp 1676037725
transform 1 0 20516 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1676037725
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_209
timestamp 1676037725
transform 1 0 20332 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1676037725
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_205
timestamp 1676037725
transform 1 0 19964 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_211
timestamp 1676037725
transform 1 0 20516 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_11
timestamp 1676037725
transform 1 0 2116 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 1676037725
transform 1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_209
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_29
timestamp 1676037725
transform 1 0 3772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_41
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1676037725
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_85
timestamp 1676037725
transform 1 0 8924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_97
timestamp 1676037725
transform 1 0 10028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 1676037725
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_141
timestamp 1676037725
transform 1 0 14076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_153
timestamp 1676037725
transform 1 0 15180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1676037725
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_197
timestamp 1676037725
transform 1 0 19228 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_209
timestamp 1676037725
transform 1 0 20332 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 20884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 20884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 20884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 20884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 20884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 20884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 20884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 20884 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 20884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 20884 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 20884 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 20884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 20884 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 20884 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 20884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 20884 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 20884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 20884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 20884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 20884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 20884 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 20884 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 20884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 20884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 3680 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 8832 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 13984 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 19136 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16928 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp 1676037725
transform 1 0 19872 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 1676037725
transform 1 0 12328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp 1676037725
transform 1 0 16100 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1676037725
transform 1 0 15548 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1676037725
transform 1 0 13524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _206_
timestamp 1676037725
transform 1 0 7452 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5428 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and4_4  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12328 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13248 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _211_
timestamp 1676037725
transform 1 0 15824 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_2  _213_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14168 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_2  _214_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14444 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _216_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14444 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1676037725
transform 1 0 17480 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_2  _221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1676037725
transform 1 0 17664 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18308 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_4  _225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16560 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__xnor2_4  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18400 0 -1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_4  _227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19780 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1676037725
transform 1 0 17572 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _229_
timestamp 1676037725
transform 1 0 15364 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19688 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18216 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_4  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__and2_2  _234_
timestamp 1676037725
transform 1 0 13064 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _235_
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _236_
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11776 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8740 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _239_
timestamp 1676037725
transform 1 0 9844 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1676037725
transform 1 0 11408 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _241_
timestamp 1676037725
transform 1 0 17296 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _242_
timestamp 1676037725
transform 1 0 15088 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _244_
timestamp 1676037725
transform 1 0 18400 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _245_
timestamp 1676037725
transform 1 0 11776 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _246_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11224 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1676037725
transform 1 0 13432 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _249_
timestamp 1676037725
transform 1 0 13248 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _250_
timestamp 1676037725
transform 1 0 16468 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8280 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _252_
timestamp 1676037725
transform 1 0 8740 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _253_
timestamp 1676037725
transform 1 0 8832 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  _254_
timestamp 1676037725
transform 1 0 10212 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1676037725
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15916 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _258_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15364 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _260_
timestamp 1676037725
transform 1 0 19688 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18584 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _262_
timestamp 1676037725
transform 1 0 16100 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _263_
timestamp 1676037725
transform 1 0 14076 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13156 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _266_
timestamp 1676037725
transform 1 0 13340 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13800 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _268_
timestamp 1676037725
transform 1 0 12972 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12788 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _270_
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10580 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12788 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _274_
timestamp 1676037725
transform 1 0 15732 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _275_
timestamp 1676037725
transform 1 0 14720 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _276_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10304 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _280_
timestamp 1676037725
transform 1 0 14536 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _283_
timestamp 1676037725
transform 1 0 18400 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _284_
timestamp 1676037725
transform 1 0 18676 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17480 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17020 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _287_
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _288_
timestamp 1676037725
transform 1 0 15824 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _289_
timestamp 1676037725
transform 1 0 16008 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _290_
timestamp 1676037725
transform 1 0 14444 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _291_
timestamp 1676037725
transform 1 0 14536 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _292_
timestamp 1676037725
transform 1 0 15640 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _293_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _294_
timestamp 1676037725
transform 1 0 18216 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _295_
timestamp 1676037725
transform 1 0 18124 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _296_
timestamp 1676037725
transform 1 0 17572 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _297_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17480 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15456 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _300_
timestamp 1676037725
transform 1 0 16468 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13984 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15180 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _304_
timestamp 1676037725
transform 1 0 12880 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _305_
timestamp 1676037725
transform 1 0 9200 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _306_
timestamp 1676037725
transform 1 0 11684 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _307_
timestamp 1676037725
transform 1 0 12512 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10396 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _309_
timestamp 1676037725
transform 1 0 9108 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _310_
timestamp 1676037725
transform 1 0 9108 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _311_
timestamp 1676037725
transform 1 0 9108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _312_
timestamp 1676037725
transform 1 0 10212 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _313_
timestamp 1676037725
transform 1 0 9108 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _314_
timestamp 1676037725
transform 1 0 2024 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16928 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _316_
timestamp 1676037725
transform 1 0 13156 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _317_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13248 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _318_
timestamp 1676037725
transform 1 0 12512 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _319_
timestamp 1676037725
transform 1 0 14260 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _320_
timestamp 1676037725
transform 1 0 14352 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _321_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13800 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _322_
timestamp 1676037725
transform 1 0 12604 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _323_
timestamp 1676037725
transform 1 0 15824 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _324_
timestamp 1676037725
transform 1 0 15456 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _325_
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _326_
timestamp 1676037725
transform 1 0 14352 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _327_
timestamp 1676037725
transform 1 0 14260 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _328_
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _329_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18308 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _330_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18216 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _331_
timestamp 1676037725
transform 1 0 1932 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_2  _332_
timestamp 1676037725
transform 1 0 6624 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_4  _333_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ai_1  _334_
timestamp 1676037725
transform 1 0 3036 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _335_
timestamp 1676037725
transform 1 0 1840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _336_
timestamp 1676037725
transform 1 0 7452 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _337_
timestamp 1676037725
transform 1 0 4324 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _338_
timestamp 1676037725
transform 1 0 7728 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _340_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3128 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1676037725
transform 1 0 1932 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _342_
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _343_
timestamp 1676037725
transform 1 0 6532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _344_
timestamp 1676037725
transform 1 0 4600 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _345_
timestamp 1676037725
transform 1 0 6532 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _346_
timestamp 1676037725
transform 1 0 7084 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _347_
timestamp 1676037725
transform 1 0 6624 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _348_
timestamp 1676037725
transform 1 0 1840 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _349_
timestamp 1676037725
transform 1 0 7728 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _350_
timestamp 1676037725
transform 1 0 7912 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1676037725
transform 1 0 7084 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1676037725
transform 1 0 6716 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _354_
timestamp 1676037725
transform 1 0 4968 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _355_
timestamp 1676037725
transform 1 0 5428 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _356_
timestamp 1676037725
transform 1 0 4968 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1676037725
transform 1 0 4876 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1676037725
transform 1 0 4784 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _359_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6900 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _360_
timestamp 1676037725
transform 1 0 4416 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _361_
timestamp 1676037725
transform 1 0 3680 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1676037725
transform 1 0 4232 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1676037725
transform 1 0 3680 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _364_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6900 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _365_
timestamp 1676037725
transform 1 0 5888 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _366_
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _367_
timestamp 1676037725
transform 1 0 5244 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _368_
timestamp 1676037725
transform 1 0 4232 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _369_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4048 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _370_
timestamp 1676037725
transform 1 0 2300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _371_
timestamp 1676037725
transform 1 0 2852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _372_
timestamp 1676037725
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _373_
timestamp 1676037725
transform 1 0 2852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1676037725
transform 1 0 12512 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _375_
timestamp 1676037725
transform 1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _376_
timestamp 1676037725
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _377_
timestamp 1676037725
transform 1 0 2944 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _378_
timestamp 1676037725
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _379_
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _380_
timestamp 1676037725
transform 1 0 7636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _381_
timestamp 1676037725
transform 1 0 5520 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _382_
timestamp 1676037725
transform 1 0 8280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _383_
timestamp 1676037725
transform 1 0 10028 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _384_
timestamp 1676037725
transform 1 0 11776 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _385_
timestamp 1676037725
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _386_
timestamp 1676037725
transform 1 0 14076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _387_
timestamp 1676037725
transform 1 0 12972 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _388_
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _389_
timestamp 1676037725
transform 1 0 14720 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _390_
timestamp 1676037725
transform 1 0 14904 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _391_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17112 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp 1676037725
transform 1 0 18032 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _393_
timestamp 1676037725
transform 1 0 16744 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _394_
timestamp 1676037725
transform 1 0 17296 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _395_
timestamp 1676037725
transform 1 0 16100 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _396_
timestamp 1676037725
transform 1 0 16928 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _397_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _398_
timestamp 1676037725
transform 1 0 17756 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _399_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9936 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1676037725
transform 1 0 9752 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _401_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6992 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _402_
timestamp 1676037725
transform 1 0 5060 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _403_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7728 0 -1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _404_
timestamp 1676037725
transform 1 0 4784 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _405_
timestamp 1676037725
transform 1 0 7084 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _406_
timestamp 1676037725
transform 1 0 5336 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _407_
timestamp 1676037725
transform 1 0 9752 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _408_
timestamp 1676037725
transform 1 0 9752 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _409_
timestamp 1676037725
transform 1 0 9752 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _410_
timestamp 1676037725
transform 1 0 10120 0 1 8704
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _411_
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _412_
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _413_
timestamp 1676037725
transform 1 0 7728 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _414_
timestamp 1676037725
transform 1 0 8924 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _415_
timestamp 1676037725
transform -1 0 4232 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _416_
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _417_
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _418_
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _419_
timestamp 1676037725
transform 1 0 6992 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _420_
timestamp 1676037725
transform 1 0 4600 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _421_
timestamp 1676037725
transform 1 0 2760 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _422_
timestamp 1676037725
transform 1 0 2760 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _423_
timestamp 1676037725
transform 1 0 2944 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _424_
timestamp 1676037725
transform 1 0 9660 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _425_
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _426_
timestamp 1676037725
transform 1 0 2024 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _427_
timestamp 1676037725
transform 1 0 2024 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _428_
timestamp 1676037725
transform 1 0 4600 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _429_
timestamp 1676037725
transform 1 0 6992 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _430_
timestamp 1676037725
transform 1 0 9568 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _431_
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _432_
timestamp 1676037725
transform 1 0 4508 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _433_
timestamp 1676037725
transform 1 0 5244 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _434_
timestamp 1676037725
transform 1 0 7084 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _435_
timestamp 1676037725
transform 1 0 9752 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _436_
timestamp 1676037725
transform 1 0 9752 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _437_
timestamp 1676037725
transform 1 0 9568 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _438_
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1676037725
transform 1 0 2576 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1676037725
transform 1 0 2576 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1676037725
transform 1 0 7820 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1676037725
transform 1 0 7820 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout4
timestamp 1676037725
transform 1 0 13340 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12880 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8004 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2392 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout8
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout9
timestamp 1676037725
transform 1 0 3956 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output2
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 590 592
<< labels >>
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 OP
port 0 nsew signal tristate
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 clk
port 1 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 rst
port 2 nsew signal input
flabel metal4 s 3416 2128 3736 19632 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 8361 2128 8681 19632 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 13306 2128 13626 19632 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 18251 2128 18571 19632 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 5888 2128 6208 19632 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
flabel metal4 s 10833 2128 11153 19632 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
flabel metal4 s 15778 2128 16098 19632 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
flabel metal4 s 20723 2128 21043 19632 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 22000 22000
<< end >>
